magic
tech sky130A
magscale 1 2
timestamp 1656996701
<< viali >>
rect 4721 20553 4755 20587
rect 5181 20553 5215 20587
rect 5825 20553 5859 20587
rect 6193 20553 6227 20587
rect 6929 20553 6963 20587
rect 10701 20553 10735 20587
rect 11713 20553 11747 20587
rect 14933 20553 14967 20587
rect 16865 20553 16899 20587
rect 18705 20553 18739 20587
rect 20085 20553 20119 20587
rect 18889 20485 18923 20519
rect 21005 20485 21039 20519
rect 4997 20417 5031 20451
rect 5733 20417 5767 20451
rect 7021 20417 7055 20451
rect 7665 20417 7699 20451
rect 10425 20417 10459 20451
rect 10517 20417 10551 20451
rect 10885 20417 10919 20451
rect 11529 20417 11563 20451
rect 14197 20417 14231 20451
rect 14749 20417 14783 20451
rect 16681 20417 16715 20451
rect 17325 20417 17359 20451
rect 18521 20417 18555 20451
rect 19441 20417 19475 20451
rect 19717 20417 19751 20451
rect 19901 20417 19935 20451
rect 20177 20417 20211 20451
rect 20729 20417 20763 20451
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 10241 20349 10275 20383
rect 20453 20349 20487 20383
rect 11069 20281 11103 20315
rect 17785 20281 17819 20315
rect 19073 20281 19107 20315
rect 21465 20281 21499 20315
rect 5273 20213 5307 20247
rect 6377 20213 6411 20247
rect 7389 20213 7423 20247
rect 7481 20213 7515 20247
rect 11253 20213 11287 20247
rect 12909 20213 12943 20247
rect 14381 20213 14415 20247
rect 15117 20213 15151 20247
rect 15485 20213 15519 20247
rect 17141 20213 17175 20247
rect 21281 20213 21315 20247
rect 4077 20009 4111 20043
rect 5641 20009 5675 20043
rect 7113 20009 7147 20043
rect 11989 20009 12023 20043
rect 13185 20009 13219 20043
rect 14197 20009 14231 20043
rect 14565 20009 14599 20043
rect 14933 20009 14967 20043
rect 15393 20009 15427 20043
rect 15761 20009 15795 20043
rect 16129 20009 16163 20043
rect 18797 20009 18831 20043
rect 19073 20009 19107 20043
rect 21465 20009 21499 20043
rect 9597 19941 9631 19975
rect 13461 19941 13495 19975
rect 7297 19873 7331 19907
rect 7481 19873 7515 19907
rect 8217 19873 8251 19907
rect 11253 19873 11287 19907
rect 17325 19873 17359 19907
rect 17877 19873 17911 19907
rect 18429 19873 18463 19907
rect 19625 19873 19659 19907
rect 20545 19873 20579 19907
rect 21097 19873 21131 19907
rect 4261 19805 4295 19839
rect 5733 19805 5767 19839
rect 5989 19805 6023 19839
rect 9045 19805 9079 19839
rect 10977 19805 11011 19839
rect 11079 19805 11113 19839
rect 11805 19805 11839 19839
rect 12909 19805 12943 19839
rect 13001 19805 13035 19839
rect 13645 19805 13679 19839
rect 14381 19805 14415 19839
rect 14749 19805 14783 19839
rect 15117 19805 15151 19839
rect 15209 19805 15243 19839
rect 15577 19805 15611 19839
rect 15945 19805 15979 19839
rect 16773 19805 16807 19839
rect 17049 19805 17083 19839
rect 17601 19805 17635 19839
rect 18153 19805 18187 19839
rect 18705 19805 18739 19839
rect 20085 19805 20119 19839
rect 20361 19805 20395 19839
rect 20913 19805 20947 19839
rect 4506 19737 4540 19771
rect 9321 19737 9355 19771
rect 10732 19737 10766 19771
rect 12633 19737 12667 19771
rect 13737 19737 13771 19771
rect 2237 19669 2271 19703
rect 2605 19669 2639 19703
rect 2881 19669 2915 19703
rect 3801 19669 3835 19703
rect 7573 19669 7607 19703
rect 7941 19669 7975 19703
rect 8309 19669 8343 19703
rect 8401 19669 8435 19703
rect 8769 19669 8803 19703
rect 11713 19669 11747 19703
rect 1961 19465 1995 19499
rect 2329 19465 2363 19499
rect 3341 19465 3375 19499
rect 3893 19465 3927 19499
rect 5365 19465 5399 19499
rect 5825 19465 5859 19499
rect 6837 19465 6871 19499
rect 7205 19465 7239 19499
rect 8677 19465 8711 19499
rect 10241 19465 10275 19499
rect 11253 19465 11287 19499
rect 13369 19465 13403 19499
rect 15301 19465 15335 19499
rect 15945 19465 15979 19499
rect 16773 19465 16807 19499
rect 17233 19465 17267 19499
rect 17877 19465 17911 19499
rect 18337 19465 18371 19499
rect 18521 19465 18555 19499
rect 2697 19397 2731 19431
rect 7564 19397 7598 19431
rect 10701 19397 10735 19431
rect 11774 19397 11808 19431
rect 14473 19397 14507 19431
rect 15025 19397 15059 19431
rect 19073 19397 19107 19431
rect 19717 19397 19751 19431
rect 20269 19397 20303 19431
rect 20821 19397 20855 19431
rect 21373 19397 21407 19431
rect 2145 19329 2179 19363
rect 2513 19329 2547 19363
rect 3249 19329 3283 19363
rect 5017 19329 5051 19363
rect 5284 19329 5318 19363
rect 5733 19329 5767 19363
rect 9025 19329 9059 19363
rect 10609 19329 10643 19363
rect 11069 19329 11103 19363
rect 11529 19329 11563 19363
rect 13185 19329 13219 19363
rect 14197 19329 14231 19363
rect 14749 19329 14783 19363
rect 15761 19329 15795 19363
rect 16957 19329 16991 19363
rect 17049 19329 17083 19363
rect 17417 19329 17451 19363
rect 18061 19329 18095 19363
rect 19349 19329 19383 19363
rect 19441 19329 19475 19363
rect 19993 19329 20027 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 3433 19261 3467 19295
rect 3801 19261 3835 19295
rect 5917 19261 5951 19295
rect 6653 19261 6687 19295
rect 6745 19261 6779 19295
rect 7297 19261 7331 19295
rect 8769 19261 8803 19295
rect 10793 19261 10827 19295
rect 13001 19261 13035 19295
rect 16497 19261 16531 19295
rect 10149 19193 10183 19227
rect 12909 19193 12943 19227
rect 2881 19125 2915 19159
rect 13921 19125 13955 19159
rect 15669 19125 15703 19159
rect 17601 19125 17635 19159
rect 18797 19125 18831 19159
rect 1593 18921 1627 18955
rect 4261 18921 4295 18955
rect 5181 18921 5215 18955
rect 8309 18921 8343 18955
rect 8493 18921 8527 18955
rect 8769 18921 8803 18955
rect 9689 18921 9723 18955
rect 10701 18921 10735 18955
rect 13001 18921 13035 18955
rect 18981 18921 19015 18955
rect 19349 18921 19383 18955
rect 21373 18921 21407 18955
rect 4169 18853 4203 18887
rect 2053 18785 2087 18819
rect 2789 18785 2823 18819
rect 3893 18785 3927 18819
rect 4629 18785 4663 18819
rect 4721 18785 4755 18819
rect 5733 18785 5767 18819
rect 5825 18785 5859 18819
rect 6193 18785 6227 18819
rect 6377 18785 6411 18819
rect 6929 18785 6963 18819
rect 9045 18785 9079 18819
rect 10057 18785 10091 18819
rect 12081 18785 12115 18819
rect 12817 18785 12851 18819
rect 13553 18785 13587 18819
rect 14197 18785 14231 18819
rect 14381 18785 14415 18819
rect 18889 18785 18923 18819
rect 1777 18717 1811 18751
rect 3065 18717 3099 18751
rect 7196 18717 7230 18751
rect 9781 18717 9815 18751
rect 13829 18717 13863 18751
rect 14473 18717 14507 18751
rect 19533 18717 19567 18751
rect 20085 18717 20119 18751
rect 20361 18717 20395 18751
rect 20637 18717 20671 18751
rect 21189 18717 21223 18751
rect 4813 18649 4847 18683
rect 6469 18649 6503 18683
rect 11814 18649 11848 18683
rect 13461 18649 13495 18683
rect 19809 18649 19843 18683
rect 20913 18649 20947 18683
rect 2145 18581 2179 18615
rect 2237 18581 2271 18615
rect 2605 18581 2639 18615
rect 2973 18581 3007 18615
rect 3433 18581 3467 18615
rect 3617 18581 3651 18615
rect 5273 18581 5307 18615
rect 5641 18581 5675 18615
rect 6837 18581 6871 18615
rect 9229 18581 9263 18615
rect 9321 18581 9355 18615
rect 10333 18581 10367 18615
rect 12173 18581 12207 18615
rect 12541 18581 12575 18615
rect 12633 18581 12667 18615
rect 13369 18581 13403 18615
rect 14841 18581 14875 18615
rect 1685 18377 1719 18411
rect 1961 18377 1995 18411
rect 4353 18377 4387 18411
rect 7389 18377 7423 18411
rect 7757 18377 7791 18411
rect 8217 18377 8251 18411
rect 8677 18377 8711 18411
rect 9137 18377 9171 18411
rect 10057 18377 10091 18411
rect 10885 18377 10919 18411
rect 10977 18377 11011 18411
rect 11897 18377 11931 18411
rect 12265 18377 12299 18411
rect 14565 18377 14599 18411
rect 15577 18377 15611 18411
rect 19809 18377 19843 18411
rect 20545 18377 20579 18411
rect 21465 18377 21499 18411
rect 1501 18309 1535 18343
rect 5558 18309 5592 18343
rect 6193 18309 6227 18343
rect 9505 18309 9539 18343
rect 13093 18309 13127 18343
rect 13452 18309 13486 18343
rect 21005 18309 21039 18343
rect 2145 18241 2179 18275
rect 3157 18241 3191 18275
rect 3985 18241 4019 18275
rect 6561 18241 6595 18275
rect 6929 18241 6963 18275
rect 7021 18241 7055 18275
rect 7849 18241 7883 18275
rect 10149 18241 10183 18275
rect 14657 18241 14691 18275
rect 19625 18241 19659 18275
rect 19993 18241 20027 18275
rect 20729 18241 20763 18275
rect 21281 18241 21315 18275
rect 2881 18173 2915 18207
rect 3065 18173 3099 18207
rect 3801 18173 3835 18207
rect 3893 18173 3927 18207
rect 5825 18173 5859 18207
rect 6837 18173 6871 18207
rect 7573 18173 7607 18207
rect 8401 18173 8435 18207
rect 8585 18173 8619 18207
rect 9597 18173 9631 18207
rect 9689 18173 9723 18207
rect 10793 18173 10827 18207
rect 11621 18173 11655 18207
rect 12357 18173 12391 18207
rect 12541 18173 12575 18207
rect 12725 18173 12759 18207
rect 13185 18173 13219 18207
rect 20177 18173 20211 18207
rect 3525 18105 3559 18139
rect 9045 18105 9079 18139
rect 11345 18105 11379 18139
rect 19349 18105 19383 18139
rect 2237 18037 2271 18071
rect 4445 18037 4479 18071
rect 6009 18037 6043 18071
rect 11713 18037 11747 18071
rect 19533 18037 19567 18071
rect 1777 17833 1811 17867
rect 4537 17833 4571 17867
rect 5365 17833 5399 17867
rect 6193 17833 6227 17867
rect 6561 17833 6595 17867
rect 7849 17833 7883 17867
rect 8769 17833 8803 17867
rect 12265 17833 12299 17867
rect 20085 17833 20119 17867
rect 21557 17833 21591 17867
rect 6469 17765 6503 17799
rect 7665 17765 7699 17799
rect 8953 17765 8987 17799
rect 9873 17765 9907 17799
rect 11345 17765 11379 17799
rect 20177 17765 20211 17799
rect 4997 17697 5031 17731
rect 5181 17697 5215 17731
rect 5917 17697 5951 17731
rect 6745 17697 6779 17731
rect 7113 17697 7147 17731
rect 7205 17697 7239 17731
rect 8217 17697 8251 17731
rect 9505 17697 9539 17731
rect 10149 17697 10183 17731
rect 10793 17697 10827 17731
rect 11989 17697 12023 17731
rect 12817 17697 12851 17731
rect 16221 17697 16255 17731
rect 1593 17629 1627 17663
rect 1961 17629 1995 17663
rect 3166 17629 3200 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 3893 17629 3927 17663
rect 7297 17629 7331 17663
rect 11805 17629 11839 17663
rect 14197 17629 14231 17663
rect 14464 17629 14498 17663
rect 16129 17629 16163 17663
rect 20361 17629 20395 17663
rect 20913 17629 20947 17663
rect 4905 17561 4939 17595
rect 9413 17561 9447 17595
rect 10977 17561 11011 17595
rect 12633 17561 12667 17595
rect 16037 17561 16071 17595
rect 20637 17561 20671 17595
rect 21189 17561 21223 17595
rect 2053 17493 2087 17527
rect 5733 17493 5767 17527
rect 5825 17493 5859 17527
rect 8309 17493 8343 17527
rect 8401 17493 8435 17527
rect 9321 17493 9355 17527
rect 10241 17493 10275 17527
rect 10885 17493 10919 17527
rect 11437 17493 11471 17527
rect 11897 17493 11931 17527
rect 12725 17493 12759 17527
rect 13093 17493 13127 17527
rect 15577 17493 15611 17527
rect 15669 17493 15703 17527
rect 16589 17493 16623 17527
rect 1777 17289 1811 17323
rect 3433 17289 3467 17323
rect 5457 17289 5491 17323
rect 7021 17289 7055 17323
rect 8217 17289 8251 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 9505 17289 9539 17323
rect 11253 17289 11287 17323
rect 11805 17289 11839 17323
rect 12449 17289 12483 17323
rect 13829 17289 13863 17323
rect 14197 17289 14231 17323
rect 14657 17289 14691 17323
rect 15025 17289 15059 17323
rect 15761 17289 15795 17323
rect 16405 17289 16439 17323
rect 20177 17289 20211 17323
rect 21005 17289 21039 17323
rect 21373 17289 21407 17323
rect 2298 17221 2332 17255
rect 3770 17221 3804 17255
rect 12909 17221 12943 17255
rect 14289 17221 14323 17255
rect 1593 17153 1627 17187
rect 1961 17153 1995 17187
rect 5273 17153 5307 17187
rect 5825 17153 5859 17187
rect 6929 17153 6963 17187
rect 7389 17153 7423 17187
rect 8585 17153 8619 17187
rect 10129 17153 10163 17187
rect 11897 17153 11931 17187
rect 12725 17153 12759 17187
rect 15117 17153 15151 17187
rect 15853 17153 15887 17187
rect 19993 17153 20027 17187
rect 20821 17153 20855 17187
rect 21189 17153 21223 17187
rect 2053 17085 2087 17119
rect 3525 17085 3559 17119
rect 5917 17085 5951 17119
rect 6009 17085 6043 17119
rect 6469 17085 6503 17119
rect 7113 17085 7147 17119
rect 7757 17085 7791 17119
rect 8125 17085 8159 17119
rect 8677 17085 8711 17119
rect 8769 17085 8803 17119
rect 9597 17085 9631 17119
rect 9873 17085 9907 17119
rect 11713 17085 11747 17119
rect 14381 17085 14415 17119
rect 15209 17085 15243 17119
rect 15577 17085 15611 17119
rect 4905 17017 4939 17051
rect 12265 17017 12299 17051
rect 12633 17017 12667 17051
rect 5089 16949 5123 16983
rect 6561 16949 6595 16983
rect 7665 16949 7699 16983
rect 16221 16949 16255 16983
rect 16773 16949 16807 16983
rect 20453 16949 20487 16983
rect 20729 16949 20763 16983
rect 1869 16745 1903 16779
rect 2789 16745 2823 16779
rect 6561 16745 6595 16779
rect 8769 16745 8803 16779
rect 9045 16745 9079 16779
rect 10885 16745 10919 16779
rect 14105 16745 14139 16779
rect 15577 16745 15611 16779
rect 17233 16745 17267 16779
rect 21005 16745 21039 16779
rect 6101 16677 6135 16711
rect 7389 16677 7423 16711
rect 17417 16677 17451 16711
rect 3525 16609 3559 16643
rect 4353 16609 4387 16643
rect 4721 16609 4755 16643
rect 7021 16609 7055 16643
rect 7205 16609 7239 16643
rect 7941 16609 7975 16643
rect 8217 16609 8251 16643
rect 8309 16609 8343 16643
rect 9965 16609 9999 16643
rect 10057 16609 10091 16643
rect 10793 16609 10827 16643
rect 11621 16609 11655 16643
rect 13277 16609 13311 16643
rect 13553 16609 13587 16643
rect 16037 16609 16071 16643
rect 16129 16609 16163 16643
rect 16957 16609 16991 16643
rect 19533 16609 19567 16643
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 2605 16541 2639 16575
rect 3341 16541 3375 16575
rect 4977 16541 5011 16575
rect 7573 16541 7607 16575
rect 8401 16541 8435 16575
rect 11529 16541 11563 16575
rect 13021 16541 13055 16575
rect 15485 16541 15519 16575
rect 19257 16541 19291 16575
rect 20821 16541 20855 16575
rect 4261 16473 4295 16507
rect 6193 16473 6227 16507
rect 13461 16473 13495 16507
rect 15218 16473 15252 16507
rect 15945 16473 15979 16507
rect 16773 16473 16807 16507
rect 20729 16473 20763 16507
rect 2881 16405 2915 16439
rect 3249 16405 3283 16439
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 6929 16405 6963 16439
rect 9505 16405 9539 16439
rect 9873 16405 9907 16439
rect 11069 16405 11103 16439
rect 11437 16405 11471 16439
rect 11897 16405 11931 16439
rect 16405 16405 16439 16439
rect 16865 16405 16899 16439
rect 21189 16405 21223 16439
rect 1961 16201 1995 16235
rect 3709 16201 3743 16235
rect 4169 16201 4203 16235
rect 4629 16201 4663 16235
rect 5457 16201 5491 16235
rect 5825 16201 5859 16235
rect 7205 16201 7239 16235
rect 7849 16201 7883 16235
rect 8401 16201 8435 16235
rect 8861 16201 8895 16235
rect 10885 16201 10919 16235
rect 11069 16201 11103 16235
rect 12909 16201 12943 16235
rect 13093 16201 13127 16235
rect 15301 16201 15335 16235
rect 15669 16201 15703 16235
rect 16129 16201 16163 16235
rect 16221 16201 16255 16235
rect 17049 16201 17083 16235
rect 17509 16201 17543 16235
rect 17969 16201 18003 16235
rect 20637 16201 20671 16235
rect 21005 16201 21039 16235
rect 21373 16201 21407 16235
rect 6561 16133 6595 16167
rect 8033 16133 8067 16167
rect 9680 16133 9714 16167
rect 12449 16133 12483 16167
rect 14228 16133 14262 16167
rect 18337 16133 18371 16167
rect 20361 16133 20395 16167
rect 2145 16065 2179 16099
rect 3341 16065 3375 16099
rect 4997 16065 5031 16099
rect 8953 16065 8987 16099
rect 9402 16065 9436 16099
rect 12541 16065 12575 16099
rect 14473 16065 14507 16099
rect 14933 16065 14967 16099
rect 15761 16065 15795 16099
rect 17877 16065 17911 16099
rect 20453 16065 20487 16099
rect 20821 16065 20855 16099
rect 21189 16065 21223 16099
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 4261 15997 4295 16031
rect 4353 15997 4387 16031
rect 5089 15997 5123 16031
rect 5181 15997 5215 16031
rect 5917 15997 5951 16031
rect 6009 15997 6043 16031
rect 7297 15997 7331 16031
rect 7481 15997 7515 16031
rect 8769 15997 8803 16031
rect 12357 15997 12391 16031
rect 14657 15997 14691 16031
rect 14841 15997 14875 16031
rect 15485 15997 15519 16031
rect 16773 15997 16807 16031
rect 16957 15997 16991 16031
rect 18153 15997 18187 16031
rect 3801 15929 3835 15963
rect 9321 15929 9355 15963
rect 2237 15861 2271 15895
rect 2513 15861 2547 15895
rect 2881 15861 2915 15895
rect 6377 15861 6411 15895
rect 6837 15861 6871 15895
rect 7665 15861 7699 15895
rect 10793 15861 10827 15895
rect 17417 15861 17451 15895
rect 1961 15657 1995 15691
rect 2329 15657 2363 15691
rect 2789 15657 2823 15691
rect 4169 15657 4203 15691
rect 6009 15657 6043 15691
rect 11897 15657 11931 15691
rect 13461 15657 13495 15691
rect 14565 15657 14599 15691
rect 15853 15657 15887 15691
rect 17877 15657 17911 15691
rect 21373 15657 21407 15691
rect 8953 15589 8987 15623
rect 13369 15589 13403 15623
rect 3433 15521 3467 15555
rect 6469 15521 6503 15555
rect 6561 15521 6595 15555
rect 7297 15521 7331 15555
rect 12541 15521 12575 15555
rect 12633 15521 12667 15555
rect 14381 15521 14415 15555
rect 15301 15521 15335 15555
rect 16405 15521 16439 15555
rect 18429 15521 18463 15555
rect 2145 15453 2179 15487
rect 2513 15453 2547 15487
rect 2605 15453 2639 15487
rect 7553 15453 7587 15487
rect 10333 15453 10367 15487
rect 10517 15453 10551 15487
rect 10784 15453 10818 15487
rect 14933 15453 14967 15487
rect 16672 15453 16706 15487
rect 18245 15453 18279 15487
rect 18337 15453 18371 15487
rect 18705 15453 18739 15487
rect 19625 15453 19659 15487
rect 19901 15453 19935 15487
rect 20821 15453 20855 15487
rect 21189 15453 21223 15487
rect 2973 15385 3007 15419
rect 5457 15385 5491 15419
rect 6377 15385 6411 15419
rect 10066 15385 10100 15419
rect 12725 15385 12759 15419
rect 14289 15385 14323 15419
rect 15393 15385 15427 15419
rect 15945 15385 15979 15419
rect 20729 15385 20763 15419
rect 4353 15317 4387 15351
rect 5273 15317 5307 15351
rect 5641 15317 5675 15351
rect 8677 15317 8711 15351
rect 12081 15317 12115 15351
rect 13093 15317 13127 15351
rect 15485 15317 15519 15351
rect 16221 15317 16255 15351
rect 17785 15317 17819 15351
rect 18889 15317 18923 15351
rect 21005 15317 21039 15351
rect 1777 15113 1811 15147
rect 4077 15113 4111 15147
rect 7941 15113 7975 15147
rect 9045 15113 9079 15147
rect 9505 15113 9539 15147
rect 9597 15113 9631 15147
rect 9965 15113 9999 15147
rect 11529 15113 11563 15147
rect 11989 15113 12023 15147
rect 13001 15113 13035 15147
rect 13461 15113 13495 15147
rect 13921 15113 13955 15147
rect 16497 15113 16531 15147
rect 17141 15113 17175 15147
rect 8677 15045 8711 15079
rect 10425 15045 10459 15079
rect 11345 15045 11379 15079
rect 16681 15045 16715 15079
rect 17500 15045 17534 15079
rect 19993 15045 20027 15079
rect 1961 14977 1995 15011
rect 2237 14977 2271 15011
rect 2513 14977 2547 15011
rect 2605 14977 2639 15011
rect 2872 14977 2906 15011
rect 4445 14977 4479 15011
rect 4537 14977 4571 15011
rect 5365 14977 5399 15011
rect 6745 14977 6779 15011
rect 7389 14977 7423 15011
rect 10333 14977 10367 15011
rect 10793 14977 10827 15011
rect 11897 14977 11931 15011
rect 13829 14977 13863 15011
rect 14933 14977 14967 15011
rect 15384 14977 15418 15011
rect 17233 14977 17267 15011
rect 18705 14977 18739 15011
rect 19717 14977 19751 15011
rect 4629 14909 4663 14943
rect 5457 14909 5491 14943
rect 5549 14909 5583 14943
rect 6929 14909 6963 14943
rect 7481 14909 7515 14943
rect 7665 14909 7699 14943
rect 8401 14909 8435 14943
rect 8585 14909 8619 14943
rect 9689 14909 9723 14943
rect 10609 14909 10643 14943
rect 11069 14909 11103 14943
rect 12081 14909 12115 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 14105 14909 14139 14943
rect 15117 14909 15151 14943
rect 3985 14841 4019 14875
rect 6561 14841 6595 14875
rect 14749 14841 14783 14875
rect 4997 14773 5031 14807
rect 7021 14773 7055 14807
rect 8217 14773 8251 14807
rect 9137 14773 9171 14807
rect 12449 14773 12483 14807
rect 13369 14773 13403 14807
rect 18613 14773 18647 14807
rect 21097 14773 21131 14807
rect 2881 14569 2915 14603
rect 4169 14569 4203 14603
rect 9873 14569 9907 14603
rect 10701 14569 10735 14603
rect 12173 14569 12207 14603
rect 19349 14569 19383 14603
rect 21373 14569 21407 14603
rect 1593 14501 1627 14535
rect 3617 14501 3651 14535
rect 15485 14501 15519 14535
rect 21005 14501 21039 14535
rect 2145 14433 2179 14467
rect 4629 14433 4663 14467
rect 4813 14433 4847 14467
rect 6377 14433 6411 14467
rect 8585 14433 8619 14467
rect 9229 14433 9263 14467
rect 9413 14433 9447 14467
rect 10057 14433 10091 14467
rect 10241 14433 10275 14467
rect 13921 14433 13955 14467
rect 15669 14433 15703 14467
rect 15853 14433 15887 14467
rect 16589 14433 16623 14467
rect 17693 14433 17727 14467
rect 1777 14365 1811 14399
rect 2329 14365 2363 14399
rect 2697 14365 2731 14399
rect 3065 14365 3099 14399
rect 3157 14365 3191 14399
rect 4537 14365 4571 14399
rect 6110 14365 6144 14399
rect 7941 14365 7975 14399
rect 8401 14365 8435 14399
rect 8493 14365 8527 14399
rect 10793 14365 10827 14399
rect 12265 14365 12299 14399
rect 12532 14365 12566 14399
rect 14105 14365 14139 14399
rect 20729 14365 20763 14399
rect 20821 14365 20855 14399
rect 21189 14365 21223 14399
rect 3433 14297 3467 14331
rect 7696 14297 7730 14331
rect 11060 14297 11094 14331
rect 14350 14297 14384 14331
rect 16681 14297 16715 14331
rect 17960 14297 17994 14331
rect 19441 14297 19475 14331
rect 2513 14229 2547 14263
rect 3985 14229 4019 14263
rect 4997 14229 5031 14263
rect 6561 14229 6595 14263
rect 8033 14229 8067 14263
rect 8953 14229 8987 14263
rect 9505 14229 9539 14263
rect 10333 14229 10367 14263
rect 13645 14229 13679 14263
rect 15945 14229 15979 14263
rect 16313 14229 16347 14263
rect 16773 14229 16807 14263
rect 17141 14229 17175 14263
rect 19073 14229 19107 14263
rect 3617 14025 3651 14059
rect 5917 14025 5951 14059
rect 6745 14025 6779 14059
rect 6837 14025 6871 14059
rect 9413 14025 9447 14059
rect 9873 14025 9907 14059
rect 10977 14025 11011 14059
rect 13369 14025 13403 14059
rect 13461 14025 13495 14059
rect 16681 14025 16715 14059
rect 17785 14025 17819 14059
rect 17877 14025 17911 14059
rect 18245 14025 18279 14059
rect 19349 14025 19383 14059
rect 19809 14025 19843 14059
rect 21005 14025 21039 14059
rect 2820 13957 2854 13991
rect 3249 13957 3283 13991
rect 3525 13957 3559 13991
rect 7450 13957 7484 13991
rect 8953 13957 8987 13991
rect 9505 13957 9539 13991
rect 10241 13957 10275 13991
rect 12357 13957 12391 13991
rect 13829 13957 13863 13991
rect 17141 13957 17175 13991
rect 3985 13889 4019 13923
rect 4537 13889 4571 13923
rect 4804 13889 4838 13923
rect 7205 13889 7239 13923
rect 11529 13889 11563 13923
rect 13001 13889 13035 13923
rect 13921 13889 13955 13923
rect 14749 13889 14783 13923
rect 15954 13889 15988 13923
rect 17049 13889 17083 13923
rect 18981 13889 19015 13923
rect 19901 13889 19935 13923
rect 20821 13889 20855 13923
rect 3065 13821 3099 13855
rect 4077 13821 4111 13855
rect 4169 13821 4203 13855
rect 6009 13821 6043 13855
rect 6929 13821 6963 13855
rect 9689 13821 9723 13855
rect 10333 13821 10367 13855
rect 10517 13821 10551 13855
rect 10885 13821 10919 13855
rect 12449 13821 12483 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 14105 13821 14139 13855
rect 14565 13821 14599 13855
rect 16221 13821 16255 13855
rect 17233 13821 17267 13855
rect 17693 13821 17727 13855
rect 18337 13821 18371 13855
rect 18705 13821 18739 13855
rect 18889 13821 18923 13855
rect 19993 13821 20027 13855
rect 20729 13821 20763 13855
rect 8585 13753 8619 13787
rect 14381 13753 14415 13787
rect 14841 13753 14875 13787
rect 19441 13753 19475 13787
rect 1685 13685 1719 13719
rect 6377 13685 6411 13719
rect 8677 13685 8711 13719
rect 9045 13685 9079 13719
rect 11161 13685 11195 13719
rect 16313 13685 16347 13719
rect 2145 13481 2179 13515
rect 4353 13481 4387 13515
rect 5181 13481 5215 13515
rect 6009 13481 6043 13515
rect 6929 13481 6963 13515
rect 13461 13481 13495 13515
rect 16773 13481 16807 13515
rect 19257 13481 19291 13515
rect 21465 13481 21499 13515
rect 8033 13413 8067 13447
rect 8953 13413 8987 13447
rect 15945 13413 15979 13447
rect 16865 13413 16899 13447
rect 20085 13413 20119 13447
rect 1593 13345 1627 13379
rect 3617 13345 3651 13379
rect 4905 13345 4939 13379
rect 5641 13345 5675 13379
rect 5825 13345 5859 13379
rect 6469 13345 6503 13379
rect 6561 13345 6595 13379
rect 7573 13345 7607 13379
rect 8585 13345 8619 13379
rect 10977 13345 11011 13379
rect 12817 13345 12851 13379
rect 13001 13345 13035 13379
rect 13645 13345 13679 13379
rect 16221 13345 16255 13379
rect 16313 13345 16347 13379
rect 17417 13345 17451 13379
rect 17693 13345 17727 13379
rect 19809 13345 19843 13379
rect 20637 13345 20671 13379
rect 1685 13277 1719 13311
rect 7481 13277 7515 13311
rect 7941 13277 7975 13311
rect 8401 13277 8435 13311
rect 10066 13277 10100 13311
rect 10333 13277 10367 13311
rect 13093 13277 13127 13311
rect 14565 13277 14599 13311
rect 17325 13277 17359 13311
rect 17960 13277 17994 13311
rect 20545 13277 20579 13311
rect 20913 13277 20947 13311
rect 21281 13277 21315 13311
rect 1777 13209 1811 13243
rect 3372 13209 3406 13243
rect 6377 13209 6411 13243
rect 7389 13209 7423 13243
rect 8493 13209 8527 13243
rect 10793 13209 10827 13243
rect 14832 13209 14866 13243
rect 16405 13209 16439 13243
rect 17233 13209 17267 13243
rect 19625 13209 19659 13243
rect 2237 13141 2271 13175
rect 3801 13141 3835 13175
rect 4261 13141 4295 13175
rect 4721 13141 4755 13175
rect 4813 13141 4847 13175
rect 5549 13141 5583 13175
rect 7021 13141 7055 13175
rect 10425 13141 10459 13175
rect 10885 13141 10919 13175
rect 11345 13141 11379 13175
rect 19073 13141 19107 13175
rect 19717 13141 19751 13175
rect 20453 13141 20487 13175
rect 21097 13141 21131 13175
rect 1593 12937 1627 12971
rect 5641 12937 5675 12971
rect 6101 12937 6135 12971
rect 7849 12937 7883 12971
rect 8309 12937 8343 12971
rect 8677 12937 8711 12971
rect 9137 12937 9171 12971
rect 9505 12937 9539 12971
rect 9965 12937 9999 12971
rect 10701 12937 10735 12971
rect 13369 12937 13403 12971
rect 15853 12937 15887 12971
rect 16773 12937 16807 12971
rect 18245 12937 18279 12971
rect 19717 12937 19751 12971
rect 19993 12937 20027 12971
rect 2850 12869 2884 12903
rect 5181 12869 5215 12903
rect 5273 12869 5307 12903
rect 17141 12869 17175 12903
rect 18582 12869 18616 12903
rect 20177 12869 20211 12903
rect 20729 12869 20763 12903
rect 1777 12801 1811 12835
rect 2053 12801 2087 12835
rect 2329 12801 2363 12835
rect 4445 12801 4479 12835
rect 4537 12801 4571 12835
rect 5917 12801 5951 12835
rect 6377 12801 6411 12835
rect 6633 12801 6667 12835
rect 8217 12801 8251 12835
rect 9045 12801 9079 12835
rect 9873 12801 9907 12835
rect 11529 12801 11563 12835
rect 11796 12801 11830 12835
rect 13921 12801 13955 12835
rect 15126 12801 15160 12835
rect 15393 12801 15427 12835
rect 17877 12801 17911 12835
rect 20453 12801 20487 12835
rect 2605 12733 2639 12767
rect 4629 12733 4663 12767
rect 5089 12733 5123 12767
rect 8401 12733 8435 12767
rect 9229 12733 9263 12767
rect 10057 12733 10091 12767
rect 10333 12733 10367 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 17693 12733 17727 12767
rect 17785 12733 17819 12767
rect 18337 12733 18371 12767
rect 7757 12665 7791 12699
rect 12909 12665 12943 12699
rect 15485 12665 15519 12699
rect 16129 12665 16163 12699
rect 16405 12665 16439 12699
rect 2513 12597 2547 12631
rect 3985 12597 4019 12631
rect 4077 12597 4111 12631
rect 10609 12597 10643 12631
rect 10977 12597 11011 12631
rect 13737 12597 13771 12631
rect 14013 12597 14047 12631
rect 15669 12597 15703 12631
rect 16865 12597 16899 12631
rect 17325 12597 17359 12631
rect 20269 12597 20303 12631
rect 21097 12597 21131 12631
rect 1593 12393 1627 12427
rect 1961 12393 1995 12427
rect 2421 12393 2455 12427
rect 3801 12393 3835 12427
rect 6285 12393 6319 12427
rect 7297 12393 7331 12427
rect 8217 12393 8251 12427
rect 12449 12393 12483 12427
rect 14565 12393 14599 12427
rect 15485 12393 15519 12427
rect 16405 12393 16439 12427
rect 18061 12393 18095 12427
rect 19349 12393 19383 12427
rect 21005 12393 21039 12427
rect 6193 12325 6227 12359
rect 7849 12325 7883 12359
rect 3065 12257 3099 12291
rect 4261 12257 4295 12291
rect 4353 12257 4387 12291
rect 4813 12257 4847 12291
rect 6837 12257 6871 12291
rect 7757 12257 7791 12291
rect 8677 12257 8711 12291
rect 13185 12257 13219 12291
rect 13829 12257 13863 12291
rect 14197 12257 14231 12291
rect 14933 12257 14967 12291
rect 16221 12257 16255 12291
rect 16957 12257 16991 12291
rect 17417 12257 17451 12291
rect 18705 12257 18739 12291
rect 1777 12189 1811 12223
rect 2145 12189 2179 12223
rect 2237 12189 2271 12223
rect 3249 12189 3283 12223
rect 11069 12189 11103 12223
rect 13001 12189 13035 12223
rect 14381 12189 14415 12223
rect 17601 12189 17635 12223
rect 18889 12189 18923 12223
rect 20177 12189 20211 12223
rect 20453 12189 20487 12223
rect 20821 12189 20855 12223
rect 4169 12121 4203 12155
rect 5080 12121 5114 12155
rect 7205 12121 7239 12155
rect 11314 12121 11348 12155
rect 13461 12121 13495 12155
rect 15117 12121 15151 12155
rect 16773 12121 16807 12155
rect 17509 12121 17543 12155
rect 18521 12121 18555 12155
rect 2789 12053 2823 12087
rect 3157 12053 3191 12087
rect 3617 12053 3651 12087
rect 4629 12053 4663 12087
rect 6653 12053 6687 12087
rect 6745 12053 6779 12087
rect 9597 12053 9631 12087
rect 12633 12053 12667 12087
rect 13093 12053 13127 12087
rect 15025 12053 15059 12087
rect 15577 12053 15611 12087
rect 15945 12053 15979 12087
rect 16037 12053 16071 12087
rect 16865 12053 16899 12087
rect 17969 12053 18003 12087
rect 18429 12053 18463 12087
rect 19441 12053 19475 12087
rect 21465 12053 21499 12087
rect 4721 11849 4755 11883
rect 5089 11849 5123 11883
rect 5733 11849 5767 11883
rect 6469 11849 6503 11883
rect 6929 11849 6963 11883
rect 7297 11849 7331 11883
rect 7665 11849 7699 11883
rect 8125 11849 8159 11883
rect 8493 11849 8527 11883
rect 11805 11849 11839 11883
rect 12265 11849 12299 11883
rect 13553 11849 13587 11883
rect 15577 11849 15611 11883
rect 16681 11849 16715 11883
rect 18705 11849 18739 11883
rect 1961 11781 1995 11815
rect 3985 11781 4019 11815
rect 4169 11781 4203 11815
rect 4905 11781 4939 11815
rect 6837 11781 6871 11815
rect 11897 11781 11931 11815
rect 12817 11781 12851 11815
rect 13645 11781 13679 11815
rect 16129 11781 16163 11815
rect 17877 11781 17911 11815
rect 18613 11781 18647 11815
rect 2237 11713 2271 11747
rect 2697 11713 2731 11747
rect 5825 11713 5859 11747
rect 8585 11713 8619 11747
rect 9505 11713 9539 11747
rect 10232 11713 10266 11747
rect 12725 11713 12759 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 14464 11713 14498 11747
rect 16037 11713 16071 11747
rect 17049 11713 17083 11747
rect 19073 11713 19107 11747
rect 19340 11713 19374 11747
rect 21005 11713 21039 11747
rect 2789 11645 2823 11679
rect 2973 11645 3007 11679
rect 5549 11645 5583 11679
rect 7021 11645 7055 11679
rect 7757 11645 7791 11679
rect 7941 11645 7975 11679
rect 8677 11645 8711 11679
rect 9229 11645 9263 11679
rect 9413 11645 9447 11679
rect 9965 11645 9999 11679
rect 11621 11645 11655 11679
rect 13001 11645 13035 11679
rect 13737 11645 13771 11679
rect 16313 11645 16347 11679
rect 17141 11645 17175 11679
rect 17233 11645 17267 11679
rect 17601 11645 17635 11679
rect 17785 11645 17819 11679
rect 18429 11645 18463 11679
rect 20821 11645 20855 11679
rect 20913 11645 20947 11679
rect 2329 11577 2363 11611
rect 6193 11577 6227 11611
rect 11345 11577 11379 11611
rect 18889 11577 18923 11611
rect 21465 11577 21499 11611
rect 5181 11509 5215 11543
rect 9045 11509 9079 11543
rect 9873 11509 9907 11543
rect 12357 11509 12391 11543
rect 13185 11509 13219 11543
rect 15669 11509 15703 11543
rect 18245 11509 18279 11543
rect 20453 11509 20487 11543
rect 21373 11509 21407 11543
rect 3065 11305 3099 11339
rect 3249 11305 3283 11339
rect 3433 11305 3467 11339
rect 4353 11305 4387 11339
rect 6745 11305 6779 11339
rect 8769 11305 8803 11339
rect 10977 11305 11011 11339
rect 14381 11305 14415 11339
rect 15301 11305 15335 11339
rect 17785 11305 17819 11339
rect 18613 11305 18647 11339
rect 19349 11305 19383 11339
rect 21097 11305 21131 11339
rect 6009 11237 6043 11271
rect 12817 11237 12851 11271
rect 15393 11237 15427 11271
rect 19441 11237 19475 11271
rect 7297 11169 7331 11203
rect 8217 11169 8251 11203
rect 9137 11169 9171 11203
rect 11345 11169 11379 11203
rect 12173 11169 12207 11203
rect 12357 11169 12391 11203
rect 13369 11169 13403 11203
rect 13461 11169 13495 11203
rect 13829 11169 13863 11203
rect 14749 11169 14783 11203
rect 14841 11169 14875 11203
rect 15853 11169 15887 11203
rect 16037 11169 16071 11203
rect 16865 11169 16899 11203
rect 17233 11169 17267 11203
rect 18061 11169 18095 11203
rect 20821 11169 20855 11203
rect 1685 11101 1719 11135
rect 4629 11101 4663 11135
rect 8953 11101 8987 11135
rect 9393 11101 9427 11135
rect 11529 11101 11563 11135
rect 12449 11101 12483 11135
rect 16681 11101 16715 11135
rect 18245 11101 18279 11135
rect 20913 11101 20947 11135
rect 1952 11033 1986 11067
rect 4874 11033 4908 11067
rect 7849 11033 7883 11067
rect 8401 11033 8435 11067
rect 11161 11033 11195 11067
rect 15761 11033 15795 11067
rect 17325 11033 17359 11067
rect 18889 11033 18923 11067
rect 20554 11033 20588 11067
rect 21281 11033 21315 11067
rect 21557 11033 21591 11067
rect 6101 10965 6135 10999
rect 6653 10965 6687 10999
rect 7113 10965 7147 10999
rect 7205 10965 7239 10999
rect 7665 10965 7699 10999
rect 8309 10965 8343 10999
rect 10517 10965 10551 10999
rect 10609 10965 10643 10999
rect 11621 10965 11655 10999
rect 11989 10965 12023 10999
rect 12909 10965 12943 10999
rect 13277 10965 13311 10999
rect 14933 10965 14967 10999
rect 16221 10965 16255 10999
rect 16589 10965 16623 10999
rect 17417 10965 17451 10999
rect 18153 10965 18187 10999
rect 18705 10965 18739 10999
rect 4261 10761 4295 10795
rect 5825 10761 5859 10795
rect 7481 10761 7515 10795
rect 8401 10761 8435 10795
rect 9873 10761 9907 10795
rect 10241 10761 10275 10795
rect 10793 10761 10827 10795
rect 12081 10761 12115 10795
rect 13829 10761 13863 10795
rect 14657 10761 14691 10795
rect 16497 10761 16531 10795
rect 17141 10761 17175 10795
rect 19349 10761 19383 10795
rect 20269 10761 20303 10795
rect 21281 10761 21315 10795
rect 3126 10693 3160 10727
rect 6377 10693 6411 10727
rect 7113 10693 7147 10727
rect 10333 10693 10367 10727
rect 10885 10693 10919 10727
rect 12532 10693 12566 10727
rect 15884 10693 15918 10727
rect 17601 10693 17635 10727
rect 1409 10625 1443 10659
rect 1676 10625 1710 10659
rect 2881 10625 2915 10659
rect 4712 10625 4746 10659
rect 7941 10625 7975 10659
rect 9514 10625 9548 10659
rect 12265 10625 12299 10659
rect 14289 10625 14323 10659
rect 17049 10625 17083 10659
rect 18236 10625 18270 10659
rect 19901 10625 19935 10659
rect 20729 10625 20763 10659
rect 4445 10557 4479 10591
rect 5917 10557 5951 10591
rect 6561 10557 6595 10591
rect 6929 10557 6963 10591
rect 7021 10557 7055 10591
rect 7757 10557 7791 10591
rect 7849 10557 7883 10591
rect 9781 10557 9815 10591
rect 10517 10557 10551 10591
rect 14105 10557 14139 10591
rect 14197 10557 14231 10591
rect 16129 10557 16163 10591
rect 17233 10557 17267 10591
rect 17969 10557 18003 10591
rect 19717 10557 19751 10591
rect 19809 10557 19843 10591
rect 20821 10557 20855 10591
rect 20913 10557 20947 10591
rect 8309 10489 8343 10523
rect 14749 10489 14783 10523
rect 16681 10489 16715 10523
rect 20361 10489 20395 10523
rect 2789 10421 2823 10455
rect 11161 10421 11195 10455
rect 13645 10421 13679 10455
rect 17693 10421 17727 10455
rect 2513 10217 2547 10251
rect 2881 10217 2915 10251
rect 5917 10217 5951 10251
rect 8033 10217 8067 10251
rect 12541 10217 12575 10251
rect 13737 10217 13771 10251
rect 15025 10217 15059 10251
rect 16129 10217 16163 10251
rect 17049 10217 17083 10251
rect 18613 10217 18647 10251
rect 18797 10217 18831 10251
rect 18981 10217 19015 10251
rect 20085 10217 20119 10251
rect 20913 10217 20947 10251
rect 7757 10149 7791 10183
rect 10793 10149 10827 10183
rect 14841 10149 14875 10183
rect 1961 10081 1995 10115
rect 3433 10081 3467 10115
rect 4537 10081 4571 10115
rect 5365 10081 5399 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 8585 10081 8619 10115
rect 9505 10081 9539 10115
rect 9597 10081 9631 10115
rect 10241 10081 10275 10115
rect 10517 10081 10551 10115
rect 11253 10081 11287 10115
rect 11437 10081 11471 10115
rect 11897 10081 11931 10115
rect 12081 10081 12115 10115
rect 12725 10081 12759 10115
rect 12909 10081 12943 10115
rect 14197 10081 14231 10115
rect 15669 10081 15703 10115
rect 15945 10081 15979 10115
rect 16405 10081 16439 10115
rect 19533 10081 19567 10115
rect 20269 10081 20303 10115
rect 3341 10013 3375 10047
rect 4721 10013 4755 10047
rect 6377 10013 6411 10047
rect 9689 10013 9723 10047
rect 10609 10013 10643 10047
rect 11161 10013 11195 10047
rect 13001 10013 13035 10047
rect 13645 10013 13679 10047
rect 14473 10013 14507 10047
rect 15485 10013 15519 10047
rect 16497 10013 16531 10047
rect 17233 10013 17267 10047
rect 20453 10013 20487 10047
rect 3249 9945 3283 9979
rect 5549 9945 5583 9979
rect 6469 9945 6503 9979
rect 7205 9945 7239 9979
rect 7941 9945 7975 9979
rect 15393 9945 15427 9979
rect 16589 9945 16623 9979
rect 17478 9945 17512 9979
rect 19625 9945 19659 9979
rect 2053 9877 2087 9911
rect 2145 9877 2179 9911
rect 4261 9877 4295 9911
rect 4629 9877 4663 9911
rect 5089 9877 5123 9911
rect 5457 9877 5491 9911
rect 6009 9877 6043 9911
rect 6837 9877 6871 9911
rect 7297 9877 7331 9911
rect 8401 9877 8435 9911
rect 8493 9877 8527 9911
rect 10057 9877 10091 9911
rect 11713 9877 11747 9911
rect 12173 9877 12207 9911
rect 13369 9877 13403 9911
rect 14381 9877 14415 9911
rect 16957 9877 16991 9911
rect 19717 9877 19751 9911
rect 20545 9877 20579 9911
rect 21005 9877 21039 9911
rect 21281 9877 21315 9911
rect 21557 9877 21591 9911
rect 1777 9673 1811 9707
rect 4169 9673 4203 9707
rect 4629 9673 4663 9707
rect 5089 9673 5123 9707
rect 7941 9673 7975 9707
rect 8309 9673 8343 9707
rect 9781 9673 9815 9707
rect 11069 9673 11103 9707
rect 19901 9673 19935 9707
rect 20729 9673 20763 9707
rect 2850 9605 2884 9639
rect 5825 9605 5859 9639
rect 6837 9605 6871 9639
rect 8668 9605 8702 9639
rect 10425 9605 10459 9639
rect 11989 9605 12023 9639
rect 13706 9605 13740 9639
rect 14933 9605 14967 9639
rect 19542 9605 19576 9639
rect 20361 9605 20395 9639
rect 2145 9537 2179 9571
rect 4997 9537 5031 9571
rect 6745 9537 6779 9571
rect 10977 9537 11011 9571
rect 11897 9537 11931 9571
rect 12817 9537 12851 9571
rect 15485 9537 15519 9571
rect 17325 9537 17359 9571
rect 20269 9537 20303 9571
rect 21097 9537 21131 9571
rect 2237 9469 2271 9503
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 5181 9469 5215 9503
rect 5917 9469 5951 9503
rect 6009 9469 6043 9503
rect 6929 9469 6963 9503
rect 7481 9469 7515 9503
rect 7757 9469 7791 9503
rect 7849 9469 7883 9503
rect 8401 9469 8435 9503
rect 11161 9469 11195 9503
rect 12173 9469 12207 9503
rect 12633 9469 12667 9503
rect 12725 9469 12759 9503
rect 13461 9469 13495 9503
rect 15209 9469 15243 9503
rect 15393 9469 15427 9503
rect 17049 9469 17083 9503
rect 17233 9469 17267 9503
rect 17969 9469 18003 9503
rect 19809 9469 19843 9503
rect 20453 9469 20487 9503
rect 21189 9469 21223 9503
rect 21281 9469 21315 9503
rect 5457 9401 5491 9435
rect 11529 9401 11563 9435
rect 17693 9401 17727 9435
rect 18245 9401 18279 9435
rect 3985 9333 4019 9367
rect 4353 9333 4387 9367
rect 4537 9333 4571 9367
rect 6377 9333 6411 9367
rect 7297 9333 7331 9367
rect 9873 9333 9907 9367
rect 10609 9333 10643 9367
rect 13185 9333 13219 9367
rect 14841 9333 14875 9367
rect 15853 9333 15887 9367
rect 16405 9333 16439 9367
rect 16681 9333 16715 9367
rect 18061 9333 18095 9367
rect 18429 9333 18463 9367
rect 2329 9129 2363 9163
rect 4445 9129 4479 9163
rect 6101 9129 6135 9163
rect 6377 9129 6411 9163
rect 7297 9129 7331 9163
rect 9045 9129 9079 9163
rect 10241 9129 10275 9163
rect 10517 9129 10551 9163
rect 12265 9129 12299 9163
rect 12541 9129 12575 9163
rect 13461 9129 13495 9163
rect 20729 9129 20763 9163
rect 8769 9061 8803 9095
rect 10057 9061 10091 9095
rect 20637 9061 20671 9095
rect 1685 8993 1719 9027
rect 2881 8993 2915 9027
rect 3341 8993 3375 9027
rect 3893 8993 3927 9027
rect 4997 8993 5031 9027
rect 5733 8993 5767 9027
rect 5825 8993 5859 9027
rect 6653 8993 6687 9027
rect 9597 8993 9631 9027
rect 11989 8993 12023 9027
rect 12817 8993 12851 9027
rect 13001 8993 13035 9027
rect 14749 8993 14783 9027
rect 15117 8993 15151 9027
rect 18429 8993 18463 9027
rect 18613 8993 18647 9027
rect 21281 8993 21315 9027
rect 3157 8925 3191 8959
rect 4905 8925 4939 8959
rect 7389 8925 7423 8959
rect 9413 8925 9447 8959
rect 11897 8925 11931 8959
rect 15301 8925 15335 8959
rect 15568 8925 15602 8959
rect 16773 8925 16807 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 1869 8857 1903 8891
rect 2697 8857 2731 8891
rect 4353 8857 4387 8891
rect 7656 8857 7690 8891
rect 11652 8857 11686 8891
rect 17018 8857 17052 8891
rect 19502 8857 19536 8891
rect 21189 8857 21223 8891
rect 1777 8789 1811 8823
rect 2237 8789 2271 8823
rect 2789 8789 2823 8823
rect 4813 8789 4847 8823
rect 5273 8789 5307 8823
rect 5641 8789 5675 8823
rect 6837 8789 6871 8823
rect 6929 8789 6963 8823
rect 9505 8789 9539 8823
rect 9965 8789 9999 8823
rect 13093 8789 13127 8823
rect 13645 8789 13679 8823
rect 14933 8789 14967 8823
rect 16681 8789 16715 8823
rect 18153 8789 18187 8823
rect 18705 8789 18739 8823
rect 19073 8789 19107 8823
rect 2053 8585 2087 8619
rect 2421 8585 2455 8619
rect 2513 8585 2547 8619
rect 4537 8585 4571 8619
rect 5089 8585 5123 8619
rect 5549 8585 5583 8619
rect 5917 8585 5951 8619
rect 6377 8585 6411 8619
rect 8953 8585 8987 8619
rect 9321 8585 9355 8619
rect 9781 8585 9815 8619
rect 12817 8585 12851 8619
rect 13553 8585 13587 8619
rect 14749 8585 14783 8619
rect 16037 8585 16071 8619
rect 16497 8585 16531 8619
rect 16957 8585 16991 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 18429 8585 18463 8619
rect 20269 8585 20303 8619
rect 20637 8585 20671 8619
rect 1593 8517 1627 8551
rect 7941 8517 7975 8551
rect 8401 8517 8435 8551
rect 10905 8517 10939 8551
rect 11805 8517 11839 8551
rect 1961 8449 1995 8483
rect 3240 8449 3274 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 7490 8449 7524 8483
rect 8677 8449 8711 8483
rect 9413 8449 9447 8483
rect 12265 8449 12299 8483
rect 12357 8449 12391 8483
rect 13185 8449 13219 8483
rect 14841 8449 14875 8483
rect 16129 8449 16163 8483
rect 17049 8449 17083 8483
rect 19542 8449 19576 8483
rect 19809 8449 19843 8483
rect 20729 8449 20763 8483
rect 1777 8381 1811 8415
rect 2605 8381 2639 8415
rect 2973 8381 3007 8415
rect 4997 8381 5031 8415
rect 5641 8381 5675 8415
rect 6101 8381 6135 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 9597 8381 9631 8415
rect 11161 8381 11195 8415
rect 12449 8381 12483 8415
rect 14657 8381 14691 8415
rect 15301 8381 15335 8415
rect 15945 8381 15979 8415
rect 16865 8381 16899 8415
rect 17969 8381 18003 8415
rect 18153 8381 18187 8415
rect 20821 8381 20855 8415
rect 21557 8381 21591 8415
rect 4353 8313 4387 8347
rect 13369 8313 13403 8347
rect 14197 8313 14231 8347
rect 15209 8313 15243 8347
rect 17509 8313 17543 8347
rect 19901 8313 19935 8347
rect 20177 8313 20211 8347
rect 8309 8245 8343 8279
rect 8861 8245 8895 8279
rect 11253 8245 11287 8279
rect 11897 8245 11931 8279
rect 13001 8245 13035 8279
rect 14289 8245 14323 8279
rect 15577 8245 15611 8279
rect 21097 8245 21131 8279
rect 21281 8245 21315 8279
rect 2881 8041 2915 8075
rect 6561 8041 6595 8075
rect 6745 8041 6779 8075
rect 7573 8041 7607 8075
rect 8953 8041 8987 8075
rect 11437 8041 11471 8075
rect 12909 8041 12943 8075
rect 13829 8041 13863 8075
rect 19073 8041 19107 8075
rect 19993 8041 20027 8075
rect 7389 7973 7423 8007
rect 17325 7973 17359 8007
rect 20821 7973 20855 8007
rect 2237 7905 2271 7939
rect 3525 7905 3559 7939
rect 4905 7905 4939 7939
rect 6837 7905 6871 7939
rect 8585 7905 8619 7939
rect 9413 7905 9447 7939
rect 9597 7905 9631 7939
rect 9873 7905 9907 7939
rect 11161 7905 11195 7939
rect 13461 7905 13495 7939
rect 16037 7905 16071 7939
rect 16129 7905 16163 7939
rect 20453 7905 20487 7939
rect 20637 7905 20671 7939
rect 21373 7905 21407 7939
rect 3801 7837 3835 7871
rect 4261 7837 4295 7871
rect 4813 7837 4847 7871
rect 5181 7837 5215 7871
rect 8401 7837 8435 7871
rect 9321 7837 9355 7871
rect 10149 7837 10183 7871
rect 11069 7837 11103 7871
rect 12561 7837 12595 7871
rect 12817 7837 12851 7871
rect 13277 7837 13311 7871
rect 14105 7837 14139 7871
rect 16681 7837 16715 7871
rect 17693 7837 17727 7871
rect 19441 7837 19475 7871
rect 20361 7837 20395 7871
rect 2329 7769 2363 7803
rect 3341 7769 3375 7803
rect 5426 7769 5460 7803
rect 10057 7769 10091 7803
rect 14372 7769 14406 7803
rect 17960 7769 17994 7803
rect 19717 7769 19751 7803
rect 1685 7701 1719 7735
rect 1961 7701 1995 7735
rect 2421 7701 2455 7735
rect 2789 7701 2823 7735
rect 3249 7701 3283 7735
rect 4353 7701 4387 7735
rect 4721 7701 4755 7735
rect 7021 7701 7055 7735
rect 7205 7701 7239 7735
rect 7757 7701 7791 7735
rect 8033 7701 8067 7735
rect 8493 7701 8527 7735
rect 10517 7701 10551 7735
rect 10609 7701 10643 7735
rect 10977 7701 11011 7735
rect 13369 7701 13403 7735
rect 15485 7701 15519 7735
rect 15577 7701 15611 7735
rect 15945 7701 15979 7735
rect 16497 7701 16531 7735
rect 16773 7701 16807 7735
rect 19349 7701 19383 7735
rect 21189 7701 21223 7735
rect 21281 7701 21315 7735
rect 2053 7497 2087 7531
rect 3157 7497 3191 7531
rect 3617 7497 3651 7531
rect 5365 7497 5399 7531
rect 7941 7497 7975 7531
rect 9413 7497 9447 7531
rect 10517 7497 10551 7531
rect 10701 7497 10735 7531
rect 11529 7497 11563 7531
rect 12357 7497 12391 7531
rect 14749 7497 14783 7531
rect 15485 7497 15519 7531
rect 16129 7497 16163 7531
rect 17693 7497 17727 7531
rect 18245 7497 18279 7531
rect 19441 7497 19475 7531
rect 21189 7497 21223 7531
rect 1961 7429 1995 7463
rect 2513 7429 2547 7463
rect 5181 7429 5215 7463
rect 5825 7429 5859 7463
rect 8300 7429 8334 7463
rect 9873 7429 9907 7463
rect 9965 7429 9999 7463
rect 10333 7429 10367 7463
rect 12725 7429 12759 7463
rect 20729 7429 20763 7463
rect 21281 7429 21315 7463
rect 1593 7361 1627 7395
rect 2421 7361 2455 7395
rect 3249 7361 3283 7395
rect 4822 7361 4856 7395
rect 5089 7361 5123 7395
rect 5733 7361 5767 7395
rect 6561 7361 6595 7395
rect 6828 7361 6862 7395
rect 8033 7361 8067 7395
rect 11897 7361 11931 7395
rect 13277 7361 13311 7395
rect 13829 7361 13863 7395
rect 14289 7361 14323 7395
rect 15577 7361 15611 7395
rect 17049 7361 17083 7395
rect 19073 7361 19107 7395
rect 19901 7361 19935 7395
rect 20821 7361 20855 7395
rect 2605 7293 2639 7327
rect 3065 7293 3099 7327
rect 5917 7293 5951 7327
rect 10057 7293 10091 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 12817 7293 12851 7327
rect 12909 7293 12943 7327
rect 14105 7293 14139 7327
rect 14841 7293 14875 7327
rect 15025 7293 15059 7327
rect 15393 7293 15427 7327
rect 16773 7293 16807 7327
rect 16957 7293 16991 7327
rect 17969 7293 18003 7327
rect 18153 7293 18187 7327
rect 18889 7293 18923 7327
rect 18981 7293 19015 7327
rect 19993 7293 20027 7327
rect 20085 7293 20119 7327
rect 20637 7293 20671 7327
rect 13461 7225 13495 7259
rect 17417 7225 17451 7259
rect 19533 7225 19567 7259
rect 21465 7225 21499 7259
rect 1777 7157 1811 7191
rect 3709 7157 3743 7191
rect 6469 7157 6503 7191
rect 9505 7157 9539 7191
rect 10977 7157 11011 7191
rect 11069 7157 11103 7191
rect 11345 7157 11379 7191
rect 13737 7157 13771 7191
rect 14381 7157 14415 7191
rect 15945 7157 15979 7191
rect 17509 7157 17543 7191
rect 18613 7157 18647 7191
rect 3065 6953 3099 6987
rect 12081 6953 12115 6987
rect 13921 6953 13955 6987
rect 15669 6953 15703 6987
rect 18889 6953 18923 6987
rect 19257 6953 19291 6987
rect 9597 6885 9631 6919
rect 1501 6817 1535 6851
rect 3617 6817 3651 6851
rect 3801 6817 3835 6851
rect 5733 6817 5767 6851
rect 5825 6817 5859 6851
rect 6929 6817 6963 6851
rect 7389 6817 7423 6851
rect 8125 6817 8159 6851
rect 8309 6817 8343 6851
rect 8953 6817 8987 6851
rect 10977 6817 11011 6851
rect 11713 6817 11747 6851
rect 12633 6817 12667 6851
rect 13001 6817 13035 6851
rect 14289 6817 14323 6851
rect 15025 6817 15059 6851
rect 19717 6817 19751 6851
rect 19809 6817 19843 6851
rect 20637 6817 20671 6851
rect 3249 6749 3283 6783
rect 7481 6749 7515 6783
rect 7573 6749 7607 6783
rect 12541 6749 12575 6783
rect 14473 6749 14507 6783
rect 17150 6749 17184 6783
rect 17417 6749 17451 6783
rect 17509 6749 17543 6783
rect 17776 6749 17810 6783
rect 20545 6749 20579 6783
rect 20913 6749 20947 6783
rect 1768 6681 1802 6715
rect 4057 6681 4091 6715
rect 5641 6681 5675 6715
rect 6837 6681 6871 6715
rect 10710 6681 10744 6715
rect 15301 6681 15335 6715
rect 15761 6681 15795 6715
rect 19625 6681 19659 6715
rect 20453 6681 20487 6715
rect 21281 6681 21315 6715
rect 2881 6613 2915 6647
rect 3341 6613 3375 6647
rect 5181 6613 5215 6647
rect 5273 6613 5307 6647
rect 6285 6613 6319 6647
rect 6377 6613 6411 6647
rect 6745 6613 6779 6647
rect 7941 6613 7975 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 9137 6613 9171 6647
rect 11069 6613 11103 6647
rect 11437 6613 11471 6647
rect 11529 6613 11563 6647
rect 11989 6613 12023 6647
rect 12449 6613 12483 6647
rect 14381 6613 14415 6647
rect 14841 6613 14875 6647
rect 15209 6613 15243 6647
rect 16037 6613 16071 6647
rect 18981 6613 19015 6647
rect 20085 6613 20119 6647
rect 21097 6613 21131 6647
rect 1593 6409 1627 6443
rect 1961 6409 1995 6443
rect 2789 6409 2823 6443
rect 3157 6409 3191 6443
rect 6009 6409 6043 6443
rect 7573 6409 7607 6443
rect 8309 6409 8343 6443
rect 8953 6409 8987 6443
rect 9137 6409 9171 6443
rect 9873 6409 9907 6443
rect 10333 6409 10367 6443
rect 10701 6409 10735 6443
rect 11529 6409 11563 6443
rect 11989 6409 12023 6443
rect 13553 6409 13587 6443
rect 15669 6409 15703 6443
rect 17417 6409 17451 6443
rect 17509 6409 17543 6443
rect 18337 6409 18371 6443
rect 19809 6409 19843 6443
rect 20177 6409 20211 6443
rect 20637 6409 20671 6443
rect 3893 6341 3927 6375
rect 3985 6341 4019 6375
rect 4598 6341 4632 6375
rect 6837 6341 6871 6375
rect 7481 6341 7515 6375
rect 8401 6341 8435 6375
rect 11897 6341 11931 6375
rect 13093 6341 13127 6375
rect 14188 6341 14222 6375
rect 15761 6341 15795 6375
rect 21465 6341 21499 6375
rect 4353 6273 4387 6307
rect 6745 6273 6779 6307
rect 11345 6273 11379 6307
rect 12541 6273 12575 6307
rect 13185 6273 13219 6307
rect 16405 6273 16439 6307
rect 17049 6273 17083 6307
rect 17877 6273 17911 6307
rect 19450 6273 19484 6307
rect 21005 6273 21039 6307
rect 21097 6273 21131 6307
rect 2053 6205 2087 6239
rect 2237 6205 2271 6239
rect 2605 6205 2639 6239
rect 2697 6205 2731 6239
rect 3249 6205 3283 6239
rect 4077 6205 4111 6239
rect 6929 6205 6963 6239
rect 7389 6205 7423 6239
rect 8125 6205 8159 6239
rect 9597 6205 9631 6239
rect 9781 6205 9815 6239
rect 10793 6205 10827 6239
rect 10885 6205 10919 6239
rect 12081 6205 12115 6239
rect 13001 6205 13035 6239
rect 13921 6205 13955 6239
rect 15485 6205 15519 6239
rect 16773 6205 16807 6239
rect 16957 6205 16991 6239
rect 17969 6205 18003 6239
rect 18061 6205 18095 6239
rect 19717 6205 19751 6239
rect 20269 6205 20303 6239
rect 20361 6205 20395 6239
rect 21189 6205 21223 6239
rect 6193 6137 6227 6171
rect 12633 6137 12667 6171
rect 15301 6137 15335 6171
rect 16221 6137 16255 6171
rect 1501 6069 1535 6103
rect 3525 6069 3559 6103
rect 5733 6069 5767 6103
rect 6377 6069 6411 6103
rect 7941 6069 7975 6103
rect 8769 6069 8803 6103
rect 10241 6069 10275 6103
rect 16129 6069 16163 6103
rect 1869 5865 1903 5899
rect 2881 5865 2915 5899
rect 4721 5865 4755 5899
rect 12173 5865 12207 5899
rect 13553 5865 13587 5899
rect 20729 5865 20763 5899
rect 5549 5797 5583 5831
rect 16497 5797 16531 5831
rect 20637 5797 20671 5831
rect 2605 5729 2639 5763
rect 3341 5729 3375 5763
rect 3525 5729 3559 5763
rect 4445 5729 4479 5763
rect 5273 5729 5307 5763
rect 6009 5729 6043 5763
rect 6101 5729 6135 5763
rect 6929 5729 6963 5763
rect 7665 5729 7699 5763
rect 7849 5729 7883 5763
rect 8217 5729 8251 5763
rect 8953 5729 8987 5763
rect 10701 5729 10735 5763
rect 11989 5729 12023 5763
rect 13185 5729 13219 5763
rect 13369 5729 13403 5763
rect 15945 5729 15979 5763
rect 16773 5729 16807 5763
rect 17877 5729 17911 5763
rect 21281 5729 21315 5763
rect 1685 5661 1719 5695
rect 5089 5661 5123 5695
rect 6745 5661 6779 5695
rect 7573 5661 7607 5695
rect 8401 5661 8435 5695
rect 9209 5661 9243 5695
rect 10885 5661 10919 5695
rect 11713 5661 11747 5695
rect 11805 5661 11839 5695
rect 12357 5661 12391 5695
rect 15402 5661 15436 5695
rect 15669 5661 15703 5695
rect 16129 5661 16163 5695
rect 16957 5661 16991 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 19257 5661 19291 5695
rect 2421 5593 2455 5627
rect 2513 5593 2547 5627
rect 5181 5593 5215 5627
rect 12633 5593 12667 5627
rect 13093 5593 13127 5627
rect 16865 5593 16899 5627
rect 18337 5593 18371 5627
rect 19524 5593 19558 5627
rect 1501 5525 1535 5559
rect 2053 5525 2087 5559
rect 3249 5525 3283 5559
rect 3801 5525 3835 5559
rect 4169 5525 4203 5559
rect 4261 5525 4295 5559
rect 5917 5525 5951 5559
rect 6377 5525 6411 5559
rect 6837 5525 6871 5559
rect 7205 5525 7239 5559
rect 8309 5525 8343 5559
rect 8769 5525 8803 5559
rect 10333 5525 10367 5559
rect 10793 5525 10827 5559
rect 11253 5525 11287 5559
rect 11345 5525 11379 5559
rect 12725 5525 12759 5559
rect 14289 5525 14323 5559
rect 16037 5525 16071 5559
rect 17325 5525 17359 5559
rect 18981 5525 19015 5559
rect 21097 5525 21131 5559
rect 21189 5525 21223 5559
rect 2329 5321 2363 5355
rect 2789 5321 2823 5355
rect 4445 5321 4479 5355
rect 5273 5321 5307 5355
rect 5457 5321 5491 5355
rect 5917 5321 5951 5355
rect 7205 5321 7239 5355
rect 7389 5321 7423 5355
rect 8309 5321 8343 5355
rect 10241 5321 10275 5355
rect 10609 5321 10643 5355
rect 10977 5321 11011 5355
rect 12449 5321 12483 5355
rect 15577 5321 15611 5355
rect 16405 5321 16439 5355
rect 17049 5321 17083 5355
rect 19533 5321 19567 5355
rect 21005 5321 21039 5355
rect 1685 5253 1719 5287
rect 3126 5253 3160 5287
rect 5089 5253 5123 5287
rect 5825 5253 5859 5287
rect 7665 5253 7699 5287
rect 9106 5253 9140 5287
rect 10517 5253 10551 5287
rect 14136 5253 14170 5287
rect 20729 5253 20763 5287
rect 1961 5185 1995 5219
rect 2421 5185 2455 5219
rect 2881 5185 2915 5219
rect 4997 5185 5031 5219
rect 6745 5185 6779 5219
rect 8401 5185 8435 5219
rect 11069 5185 11103 5219
rect 12541 5185 12575 5219
rect 14841 5185 14875 5219
rect 15485 5185 15519 5219
rect 18153 5185 18187 5219
rect 18409 5185 18443 5219
rect 19993 5185 20027 5219
rect 20453 5185 20487 5219
rect 21281 5185 21315 5219
rect 2237 5117 2271 5151
rect 4813 5117 4847 5151
rect 6009 5117 6043 5151
rect 6837 5117 6871 5151
rect 7021 5117 7055 5151
rect 8217 5117 8251 5151
rect 8861 5117 8895 5151
rect 11207 5117 11241 5151
rect 11529 5117 11563 5151
rect 12357 5117 12391 5151
rect 14381 5117 14415 5151
rect 15761 5117 15795 5151
rect 16129 5117 16163 5151
rect 16773 5117 16807 5151
rect 16957 5117 16991 5151
rect 18061 5117 18095 5151
rect 19717 5117 19751 5151
rect 19901 5117 19935 5151
rect 4261 5049 4295 5083
rect 12909 5049 12943 5083
rect 16037 5049 16071 5083
rect 17693 5049 17727 5083
rect 20361 5049 20395 5083
rect 4537 4981 4571 5015
rect 6377 4981 6411 5015
rect 7849 4981 7883 5015
rect 8769 4981 8803 5015
rect 11713 4981 11747 5015
rect 11897 4981 11931 5015
rect 13001 4981 13035 5015
rect 14473 4981 14507 5015
rect 14657 4981 14691 5015
rect 17417 4981 17451 5015
rect 21557 4981 21591 5015
rect 1777 4777 1811 4811
rect 3893 4777 3927 4811
rect 6377 4777 6411 4811
rect 8217 4777 8251 4811
rect 8953 4777 8987 4811
rect 9873 4777 9907 4811
rect 10793 4777 10827 4811
rect 11805 4777 11839 4811
rect 12265 4777 12299 4811
rect 16773 4777 16807 4811
rect 18245 4777 18279 4811
rect 20361 4777 20395 4811
rect 3341 4709 3375 4743
rect 5457 4709 5491 4743
rect 8769 4709 8803 4743
rect 20085 4709 20119 4743
rect 20453 4709 20487 4743
rect 20729 4709 20763 4743
rect 3157 4641 3191 4675
rect 4445 4641 4479 4675
rect 4905 4641 4939 4675
rect 4997 4641 5031 4675
rect 6009 4641 6043 4675
rect 6101 4641 6135 4675
rect 7021 4641 7055 4675
rect 7205 4641 7239 4675
rect 8033 4641 8067 4675
rect 8493 4641 8527 4675
rect 9505 4641 9539 4675
rect 10425 4641 10459 4675
rect 11253 4641 11287 4675
rect 12909 4641 12943 4675
rect 13645 4641 13679 4675
rect 14565 4641 14599 4675
rect 15669 4641 15703 4675
rect 15853 4641 15887 4675
rect 16221 4641 16255 4675
rect 16865 4641 16899 4675
rect 18981 4641 19015 4675
rect 19809 4641 19843 4675
rect 9321 4573 9355 4607
rect 9413 4573 9447 4607
rect 10241 4573 10275 4607
rect 10333 4573 10367 4607
rect 11437 4573 11471 4607
rect 12633 4573 12667 4607
rect 13553 4573 13587 4607
rect 14749 4573 14783 4607
rect 15577 4573 15611 4607
rect 16405 4573 16439 4607
rect 19625 4573 19659 4607
rect 2912 4505 2946 4539
rect 4353 4505 4387 4539
rect 5917 4505 5951 4539
rect 6929 4505 6963 4539
rect 12081 4505 12115 4539
rect 13461 4505 13495 4539
rect 14105 4505 14139 4539
rect 17132 4505 17166 4539
rect 18797 4505 18831 4539
rect 21373 4505 21407 4539
rect 1593 4437 1627 4471
rect 3433 4437 3467 4471
rect 4261 4437 4295 4471
rect 5089 4437 5123 4471
rect 5549 4437 5583 4471
rect 6561 4437 6595 4471
rect 7389 4437 7423 4471
rect 7757 4437 7791 4471
rect 7849 4437 7883 4471
rect 10885 4437 10919 4471
rect 11345 4437 11379 4471
rect 11989 4437 12023 4471
rect 12725 4437 12759 4471
rect 13093 4437 13127 4471
rect 14657 4437 14691 4471
rect 15117 4437 15151 4471
rect 15209 4437 15243 4471
rect 16313 4437 16347 4471
rect 18337 4437 18371 4471
rect 18705 4437 18739 4471
rect 19257 4437 19291 4471
rect 19717 4437 19751 4471
rect 21189 4437 21223 4471
rect 21557 4437 21591 4471
rect 2697 4233 2731 4267
rect 2973 4233 3007 4267
rect 6009 4233 6043 4267
rect 8585 4233 8619 4267
rect 9137 4233 9171 4267
rect 9781 4233 9815 4267
rect 13093 4233 13127 4267
rect 14657 4233 14691 4267
rect 17601 4233 17635 4267
rect 18429 4233 18463 4267
rect 18521 4233 18555 4267
rect 19349 4233 19383 4267
rect 2329 4165 2363 4199
rect 5672 4165 5706 4199
rect 7104 4165 7138 4199
rect 9965 4165 9999 4199
rect 10977 4165 11011 4199
rect 16865 4165 16899 4199
rect 2881 4097 2915 4131
rect 4097 4097 4131 4131
rect 5917 4097 5951 4131
rect 6837 4097 6871 4131
rect 8677 4097 8711 4131
rect 9321 4097 9355 4131
rect 10057 4097 10091 4131
rect 12357 4097 12391 4131
rect 13185 4097 13219 4131
rect 15117 4097 15151 4131
rect 15384 4097 15418 4131
rect 17049 4097 17083 4131
rect 17693 4097 17727 4131
rect 19441 4097 19475 4131
rect 2145 4029 2179 4063
rect 2237 4029 2271 4063
rect 4353 4029 4387 4063
rect 6561 4029 6595 4063
rect 8401 4029 8435 4063
rect 10333 4029 10367 4063
rect 11069 4029 11103 4063
rect 11253 4029 11287 4063
rect 11621 4029 11655 4063
rect 12081 4029 12115 4063
rect 12265 4029 12299 4063
rect 13001 4029 13035 4063
rect 14197 4029 14231 4063
rect 14749 4029 14783 4063
rect 14933 4029 14967 4063
rect 16773 4029 16807 4063
rect 17509 4029 17543 4063
rect 18245 4029 18279 4063
rect 19533 4029 19567 4063
rect 6469 3961 6503 3995
rect 9045 3961 9079 3995
rect 16497 3961 16531 3995
rect 18061 3961 18095 3995
rect 18889 3961 18923 3995
rect 19901 3961 19935 3995
rect 1777 3893 1811 3927
rect 4537 3893 4571 3927
rect 8217 3893 8251 3927
rect 9505 3893 9539 3927
rect 10609 3893 10643 3927
rect 11805 3893 11839 3927
rect 12725 3893 12759 3927
rect 13553 3893 13587 3927
rect 13829 3893 13863 3927
rect 14289 3893 14323 3927
rect 18981 3893 19015 3927
rect 20085 3893 20119 3927
rect 2053 3689 2087 3723
rect 4077 3689 4111 3723
rect 5181 3689 5215 3723
rect 6009 3689 6043 3723
rect 8677 3689 8711 3723
rect 14105 3689 14139 3723
rect 15761 3689 15795 3723
rect 17325 3689 17359 3723
rect 18153 3689 18187 3723
rect 19257 3689 19291 3723
rect 4997 3621 5031 3655
rect 10425 3621 10459 3655
rect 12357 3621 12391 3655
rect 17233 3621 17267 3655
rect 2513 3553 2547 3587
rect 2605 3553 2639 3587
rect 3525 3553 3559 3587
rect 4721 3553 4755 3587
rect 5641 3553 5675 3587
rect 5825 3553 5859 3587
rect 8125 3553 8159 3587
rect 11989 3553 12023 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15485 3553 15519 3587
rect 16313 3553 16347 3587
rect 17785 3553 17819 3587
rect 17877 3553 17911 3587
rect 18705 3553 18739 3587
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 5549 3485 5583 3519
rect 6193 3485 6227 3519
rect 7665 3485 7699 3519
rect 8953 3485 8987 3519
rect 12173 3485 12207 3519
rect 13921 3485 13955 3519
rect 15301 3485 15335 3519
rect 15393 3485 15427 3519
rect 16129 3485 16163 3519
rect 16957 3485 16991 3519
rect 18613 3485 18647 3519
rect 3341 3417 3375 3451
rect 4537 3417 4571 3451
rect 6460 3417 6494 3451
rect 8217 3417 8251 3451
rect 9198 3417 9232 3451
rect 11744 3417 11778 3451
rect 13676 3417 13710 3451
rect 16773 3417 16807 3451
rect 17693 3417 17727 3451
rect 18521 3417 18555 3451
rect 18981 3417 19015 3451
rect 2421 3349 2455 3383
rect 2881 3349 2915 3383
rect 4445 3349 4479 3383
rect 7573 3349 7607 3383
rect 8309 3349 8343 3383
rect 10333 3349 10367 3383
rect 10609 3349 10643 3383
rect 12541 3349 12575 3383
rect 14473 3349 14507 3383
rect 14933 3349 14967 3383
rect 16221 3349 16255 3383
rect 16681 3349 16715 3383
rect 2697 3145 2731 3179
rect 3157 3145 3191 3179
rect 3709 3145 3743 3179
rect 7297 3145 7331 3179
rect 8585 3145 8619 3179
rect 8953 3145 8987 3179
rect 11345 3145 11379 3179
rect 13645 3145 13679 3179
rect 14013 3145 14047 3179
rect 16405 3145 16439 3179
rect 8217 3077 8251 3111
rect 10210 3077 10244 3111
rect 11805 3077 11839 3111
rect 13286 3077 13320 3111
rect 14105 3077 14139 3111
rect 3065 3009 3099 3043
rect 5733 3009 5767 3043
rect 6377 3009 6411 3043
rect 7389 3009 7423 3043
rect 9045 3009 9079 3043
rect 9873 3009 9907 3043
rect 11529 3009 11563 3043
rect 14749 3009 14783 3043
rect 15117 3009 15151 3043
rect 15301 3009 15335 3043
rect 15853 3009 15887 3043
rect 16681 3009 16715 3043
rect 17325 3009 17359 3043
rect 17417 3009 17451 3043
rect 17785 3009 17819 3043
rect 18153 3009 18187 3043
rect 18521 3009 18555 3043
rect 18889 3009 18923 3043
rect 19257 3009 19291 3043
rect 3249 2941 3283 2975
rect 6653 2941 6687 2975
rect 6929 2941 6963 2975
rect 7113 2941 7147 2975
rect 7941 2941 7975 2975
rect 8125 2941 8159 2975
rect 8861 2941 8895 2975
rect 9965 2941 9999 2975
rect 13553 2941 13587 2975
rect 14197 2941 14231 2975
rect 15577 2941 15611 2975
rect 16129 2941 16163 2975
rect 7757 2873 7791 2907
rect 14933 2873 14967 2907
rect 17141 2873 17175 2907
rect 18337 2873 18371 2907
rect 19073 2873 19107 2907
rect 3893 2805 3927 2839
rect 4997 2805 5031 2839
rect 9413 2805 9447 2839
rect 9689 2805 9723 2839
rect 12173 2805 12207 2839
rect 14565 2805 14599 2839
rect 16865 2805 16899 2839
rect 17601 2805 17635 2839
rect 17969 2805 18003 2839
rect 18705 2805 18739 2839
rect 3801 2601 3835 2635
rect 6193 2601 6227 2635
rect 7573 2601 7607 2635
rect 7665 2601 7699 2635
rect 8953 2601 8987 2635
rect 11253 2601 11287 2635
rect 11897 2601 11931 2635
rect 14565 2601 14599 2635
rect 16681 2601 16715 2635
rect 17325 2601 17359 2635
rect 17693 2601 17727 2635
rect 18061 2601 18095 2635
rect 18429 2601 18463 2635
rect 3341 2533 3375 2567
rect 9781 2533 9815 2567
rect 11713 2533 11747 2567
rect 13645 2533 13679 2567
rect 14933 2533 14967 2567
rect 16221 2533 16255 2567
rect 3617 2465 3651 2499
rect 4261 2465 4295 2499
rect 4445 2465 4479 2499
rect 7021 2465 7055 2499
rect 8309 2465 8343 2499
rect 9505 2465 9539 2499
rect 10793 2465 10827 2499
rect 12725 2465 12759 2499
rect 14289 2465 14323 2499
rect 15853 2465 15887 2499
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 5080 2397 5114 2431
rect 8033 2397 8067 2431
rect 9321 2397 9355 2431
rect 10057 2397 10091 2431
rect 10609 2397 10643 2431
rect 11529 2397 11563 2431
rect 12909 2397 12943 2431
rect 13001 2397 13035 2431
rect 14749 2397 14783 2431
rect 15393 2397 15427 2431
rect 15485 2397 15519 2431
rect 16037 2397 16071 2431
rect 16865 2397 16899 2431
rect 6469 2329 6503 2363
rect 6745 2329 6779 2363
rect 8125 2329 8159 2363
rect 10333 2329 10367 2363
rect 4721 2261 4755 2295
rect 7113 2261 7147 2295
rect 7205 2261 7239 2295
rect 8493 2261 8527 2295
rect 8677 2261 8711 2295
rect 9413 2261 9447 2295
rect 13185 2261 13219 2295
rect 15209 2261 15243 2295
rect 15669 2261 15703 2295
rect 17049 2261 17083 2295
<< metal1 >>
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 10962 20992 10968 21004
rect 3936 20964 10968 20992
rect 3936 20952 3942 20964
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 20530 20788 20536 20800
rect 4120 20760 20536 20788
rect 4120 20748 4126 20760
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 4709 20587 4767 20593
rect 4709 20584 4721 20587
rect 992 20556 4721 20584
rect 992 20544 998 20556
rect 4709 20553 4721 20556
rect 4755 20584 4767 20587
rect 5169 20587 5227 20593
rect 5169 20584 5181 20587
rect 4755 20556 5181 20584
rect 4755 20553 4767 20556
rect 4709 20547 4767 20553
rect 5169 20553 5181 20556
rect 5215 20584 5227 20587
rect 5810 20584 5816 20596
rect 5215 20556 5816 20584
rect 5215 20553 5227 20556
rect 5169 20547 5227 20553
rect 5810 20544 5816 20556
rect 5868 20544 5874 20596
rect 6181 20587 6239 20593
rect 6181 20553 6193 20587
rect 6227 20584 6239 20587
rect 6917 20587 6975 20593
rect 6917 20584 6929 20587
rect 6227 20556 6929 20584
rect 6227 20553 6239 20556
rect 6181 20547 6239 20553
rect 6917 20553 6929 20556
rect 6963 20553 6975 20587
rect 6917 20547 6975 20553
rect 10689 20587 10747 20593
rect 10689 20553 10701 20587
rect 10735 20584 10747 20587
rect 10870 20584 10876 20596
rect 10735 20556 10876 20584
rect 10735 20553 10747 20556
rect 10689 20547 10747 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20584 11759 20587
rect 12342 20584 12348 20596
rect 11747 20556 12348 20584
rect 11747 20553 11759 20556
rect 11701 20547 11759 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 14921 20587 14979 20593
rect 14921 20553 14933 20587
rect 14967 20584 14979 20587
rect 15286 20584 15292 20596
rect 14967 20556 15292 20584
rect 14967 20553 14979 20556
rect 14921 20547 14979 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 16853 20587 16911 20593
rect 16853 20553 16865 20587
rect 16899 20584 16911 20587
rect 17126 20584 17132 20596
rect 16899 20556 17132 20584
rect 16899 20553 16911 20556
rect 16853 20547 16911 20553
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 18693 20587 18751 20593
rect 18693 20553 18705 20587
rect 18739 20584 18751 20587
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 18739 20556 20085 20584
rect 18739 20553 18751 20556
rect 18693 20547 18751 20553
rect 20073 20553 20085 20556
rect 20119 20584 20131 20587
rect 20438 20584 20444 20596
rect 20119 20556 20444 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20438 20544 20444 20556
rect 20496 20544 20502 20596
rect 5074 20476 5080 20528
rect 5132 20516 5138 20528
rect 18877 20519 18935 20525
rect 5132 20488 11376 20516
rect 5132 20476 5138 20488
rect 4985 20451 5043 20457
rect 4985 20417 4997 20451
rect 5031 20448 5043 20451
rect 5534 20448 5540 20460
rect 5031 20420 5540 20448
rect 5031 20417 5043 20420
rect 4985 20411 5043 20417
rect 5534 20408 5540 20420
rect 5592 20448 5598 20460
rect 5721 20451 5779 20457
rect 5721 20448 5733 20451
rect 5592 20420 5733 20448
rect 5592 20408 5598 20420
rect 5721 20417 5733 20420
rect 5767 20417 5779 20451
rect 7009 20451 7067 20457
rect 7009 20448 7021 20451
rect 5721 20411 5779 20417
rect 5828 20420 7021 20448
rect 5626 20380 5632 20392
rect 5587 20352 5632 20380
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 5828 20380 5856 20420
rect 7009 20417 7021 20420
rect 7055 20448 7067 20451
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 7055 20420 7665 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 7653 20417 7665 20420
rect 7699 20448 7711 20451
rect 8294 20448 8300 20460
rect 7699 20420 8300 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 10410 20448 10416 20460
rect 10371 20420 10416 20448
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 10502 20408 10508 20460
rect 10560 20448 10566 20460
rect 10873 20451 10931 20457
rect 10560 20420 10605 20448
rect 10560 20408 10566 20420
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 5736 20352 5856 20380
rect 6825 20383 6883 20389
rect 1302 20272 1308 20324
rect 1360 20312 1366 20324
rect 5736 20312 5764 20352
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 7098 20380 7104 20392
rect 6871 20352 7104 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7098 20340 7104 20352
rect 7156 20340 7162 20392
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10888 20380 10916 20411
rect 10275 20352 10916 20380
rect 11348 20380 11376 20488
rect 18877 20485 18889 20519
rect 18923 20516 18935 20519
rect 20990 20516 20996 20528
rect 18923 20488 19748 20516
rect 20951 20488 20996 20516
rect 18923 20485 18935 20488
rect 18877 20479 18935 20485
rect 11514 20448 11520 20460
rect 11475 20420 11520 20448
rect 11514 20408 11520 20420
rect 11572 20408 11578 20460
rect 14185 20451 14243 20457
rect 14185 20417 14197 20451
rect 14231 20448 14243 20451
rect 14366 20448 14372 20460
rect 14231 20420 14372 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 14737 20451 14795 20457
rect 14737 20448 14749 20451
rect 14516 20420 14749 20448
rect 14516 20408 14522 20420
rect 14737 20417 14749 20420
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17218 20448 17224 20460
rect 16715 20420 17224 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 18506 20448 18512 20460
rect 17359 20420 18512 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 18506 20408 18512 20420
rect 18564 20448 18570 20460
rect 18966 20448 18972 20460
rect 18564 20420 18972 20448
rect 18564 20408 18570 20420
rect 18966 20408 18972 20420
rect 19024 20408 19030 20460
rect 19426 20448 19432 20460
rect 19387 20420 19432 20448
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 19720 20457 19748 20488
rect 20990 20476 20996 20488
rect 21048 20476 21054 20528
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20448 19763 20451
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 19751 20420 19901 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 19889 20417 19901 20420
rect 19935 20448 19947 20451
rect 20070 20448 20076 20460
rect 19935 20420 20076 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 20717 20451 20775 20457
rect 20717 20448 20729 20451
rect 20220 20420 20265 20448
rect 20364 20420 20729 20448
rect 20220 20408 20226 20420
rect 11348 20352 12020 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 1360 20284 5764 20312
rect 1360 20272 1366 20284
rect 5902 20272 5908 20324
rect 5960 20312 5966 20324
rect 10594 20312 10600 20324
rect 5960 20284 10600 20312
rect 5960 20272 5966 20284
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 11057 20315 11115 20321
rect 11057 20281 11069 20315
rect 11103 20312 11115 20315
rect 11698 20312 11704 20324
rect 11103 20284 11704 20312
rect 11103 20281 11115 20284
rect 11057 20275 11115 20281
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 11992 20312 12020 20352
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 18414 20380 18420 20392
rect 12124 20352 18420 20380
rect 12124 20340 12130 20352
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 18984 20380 19012 20408
rect 20364 20380 20392 20420
rect 20717 20417 20729 20420
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 18984 20352 20392 20380
rect 20441 20383 20499 20389
rect 20441 20349 20453 20383
rect 20487 20380 20499 20383
rect 21542 20380 21548 20392
rect 20487 20352 21548 20380
rect 20487 20349 20499 20352
rect 20441 20343 20499 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 16758 20312 16764 20324
rect 11992 20284 16764 20312
rect 16758 20272 16764 20284
rect 16816 20272 16822 20324
rect 17586 20272 17592 20324
rect 17644 20312 17650 20324
rect 17773 20315 17831 20321
rect 17773 20312 17785 20315
rect 17644 20284 17785 20312
rect 17644 20272 17650 20284
rect 17773 20281 17785 20284
rect 17819 20312 17831 20315
rect 19061 20315 19119 20321
rect 19061 20312 19073 20315
rect 17819 20284 19073 20312
rect 17819 20281 17831 20284
rect 17773 20275 17831 20281
rect 19061 20281 19073 20284
rect 19107 20312 19119 20315
rect 19334 20312 19340 20324
rect 19107 20284 19340 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 19702 20272 19708 20324
rect 19760 20312 19766 20324
rect 21453 20315 21511 20321
rect 21453 20312 21465 20315
rect 19760 20284 21465 20312
rect 19760 20272 19766 20284
rect 21453 20281 21465 20284
rect 21499 20281 21511 20315
rect 21453 20275 21511 20281
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 4706 20244 4712 20256
rect 3752 20216 4712 20244
rect 3752 20204 3758 20216
rect 4706 20204 4712 20216
rect 4764 20204 4770 20256
rect 5258 20244 5264 20256
rect 5219 20216 5264 20244
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5442 20204 5448 20256
rect 5500 20244 5506 20256
rect 6365 20247 6423 20253
rect 6365 20244 6377 20247
rect 5500 20216 6377 20244
rect 5500 20204 5506 20216
rect 6365 20213 6377 20216
rect 6411 20213 6423 20247
rect 7374 20244 7380 20256
rect 7335 20216 7380 20244
rect 6365 20207 6423 20213
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 7524 20216 7569 20244
rect 7524 20204 7530 20216
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 11204 20216 11253 20244
rect 11204 20204 11210 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11241 20207 11299 20213
rect 12897 20247 12955 20253
rect 12897 20213 12909 20247
rect 12943 20244 12955 20247
rect 12986 20244 12992 20256
rect 12943 20216 12992 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 12986 20204 12992 20216
rect 13044 20204 13050 20256
rect 14369 20247 14427 20253
rect 14369 20213 14381 20247
rect 14415 20244 14427 20247
rect 14734 20244 14740 20256
rect 14415 20216 14740 20244
rect 14415 20213 14427 20216
rect 14369 20207 14427 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 15102 20244 15108 20256
rect 15063 20216 15108 20244
rect 15102 20204 15108 20216
rect 15160 20204 15166 20256
rect 15470 20244 15476 20256
rect 15431 20216 15476 20244
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 17129 20247 17187 20253
rect 17129 20213 17141 20247
rect 17175 20244 17187 20247
rect 17218 20244 17224 20256
rect 17175 20216 17224 20244
rect 17175 20213 17187 20216
rect 17129 20207 17187 20213
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 19352 20244 19380 20272
rect 19886 20244 19892 20256
rect 19352 20216 19892 20244
rect 19886 20204 19892 20216
rect 19944 20244 19950 20256
rect 20162 20244 20168 20256
rect 19944 20216 20168 20244
rect 19944 20204 19950 20216
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1670 20000 1676 20052
rect 1728 20040 1734 20052
rect 4065 20043 4123 20049
rect 4065 20040 4077 20043
rect 1728 20012 4077 20040
rect 1728 20000 1734 20012
rect 4065 20009 4077 20012
rect 4111 20040 4123 20043
rect 5442 20040 5448 20052
rect 4111 20012 5448 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 7098 20040 7104 20052
rect 7059 20012 7104 20040
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7650 20000 7656 20052
rect 7708 20040 7714 20052
rect 11790 20040 11796 20052
rect 7708 20012 11796 20040
rect 7708 20000 7714 20012
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 11974 20040 11980 20052
rect 11935 20012 11980 20040
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13173 20043 13231 20049
rect 13173 20040 13185 20043
rect 13136 20012 13185 20040
rect 13136 20000 13142 20012
rect 13173 20009 13185 20012
rect 13219 20009 13231 20043
rect 13173 20003 13231 20009
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13596 20012 14197 20040
rect 13596 20000 13602 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14553 20043 14611 20049
rect 14553 20040 14565 20043
rect 14332 20012 14565 20040
rect 14332 20000 14338 20012
rect 14553 20009 14565 20012
rect 14599 20009 14611 20043
rect 14553 20003 14611 20009
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14700 20012 14933 20040
rect 14700 20000 14706 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15381 20043 15439 20049
rect 15381 20040 15393 20043
rect 15252 20012 15393 20040
rect 15252 20000 15258 20012
rect 15381 20009 15393 20012
rect 15427 20009 15439 20043
rect 15381 20003 15439 20009
rect 15654 20000 15660 20052
rect 15712 20040 15718 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15712 20012 15761 20040
rect 15712 20000 15718 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 16942 20040 16948 20052
rect 16163 20012 16948 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18656 20012 18797 20040
rect 18656 20000 18662 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 19061 20043 19119 20049
rect 19061 20009 19073 20043
rect 19107 20040 19119 20043
rect 20806 20040 20812 20052
rect 19107 20012 20812 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 5644 19904 5672 20000
rect 7006 19932 7012 19984
rect 7064 19972 7070 19984
rect 9585 19975 9643 19981
rect 9585 19972 9597 19975
rect 7064 19944 9597 19972
rect 7064 19932 7070 19944
rect 9585 19941 9597 19944
rect 9631 19941 9643 19975
rect 9585 19935 9643 19941
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 11112 19944 12434 19972
rect 11112 19932 11118 19944
rect 7282 19904 7288 19916
rect 5644 19876 5856 19904
rect 7243 19876 7288 19904
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4212 19808 4261 19836
rect 4212 19796 4218 19808
rect 4249 19805 4261 19808
rect 4295 19836 4307 19839
rect 5258 19836 5264 19848
rect 4295 19808 5264 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 5258 19796 5264 19808
rect 5316 19836 5322 19848
rect 5626 19836 5632 19848
rect 5316 19808 5632 19836
rect 5316 19796 5322 19808
rect 5626 19796 5632 19808
rect 5684 19836 5690 19848
rect 5721 19839 5779 19845
rect 5721 19836 5733 19839
rect 5684 19808 5733 19836
rect 5684 19796 5690 19808
rect 5721 19805 5733 19808
rect 5767 19805 5779 19839
rect 5828 19836 5856 19876
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 7469 19907 7527 19913
rect 7469 19904 7481 19907
rect 7432 19876 7481 19904
rect 7432 19864 7438 19876
rect 7469 19873 7481 19876
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8662 19904 8668 19916
rect 8251 19876 8668 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 11146 19904 11152 19916
rect 10980 19876 11152 19904
rect 5977 19839 6035 19845
rect 5977 19836 5989 19839
rect 5828 19808 5989 19836
rect 5721 19799 5779 19805
rect 5977 19805 5989 19808
rect 6023 19805 6035 19839
rect 7300 19836 7328 19864
rect 7742 19836 7748 19848
rect 7300 19808 7748 19836
rect 5977 19799 6035 19805
rect 7742 19796 7748 19808
rect 7800 19796 7806 19848
rect 9030 19836 9036 19848
rect 8991 19808 9036 19836
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 10980 19845 11008 19876
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19873 11299 19907
rect 12406 19904 12434 19944
rect 12710 19932 12716 19984
rect 12768 19972 12774 19984
rect 13449 19975 13507 19981
rect 13449 19972 13461 19975
rect 12768 19944 13461 19972
rect 12768 19932 12774 19944
rect 13449 19941 13461 19944
rect 13495 19941 13507 19975
rect 13449 19935 13507 19941
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 12406 19876 17325 19904
rect 11241 19867 11299 19873
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10612 19808 10977 19836
rect 10612 19780 10640 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11054 19796 11060 19848
rect 11112 19845 11118 19848
rect 11112 19839 11125 19845
rect 11113 19836 11125 19839
rect 11256 19836 11284 19867
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 17865 19907 17923 19913
rect 17865 19904 17877 19907
rect 17828 19876 17877 19904
rect 17828 19864 17834 19876
rect 17865 19873 17877 19876
rect 17911 19873 17923 19907
rect 18414 19904 18420 19916
rect 18375 19876 18420 19904
rect 17865 19867 17923 19873
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 11514 19836 11520 19848
rect 11113 19808 11157 19836
rect 11256 19808 11520 19836
rect 11113 19805 11125 19808
rect 11112 19799 11125 19805
rect 11112 19796 11118 19799
rect 11514 19796 11520 19808
rect 11572 19796 11578 19848
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11756 19808 11805 19836
rect 11756 19796 11762 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 12894 19836 12900 19848
rect 12855 19808 12900 19836
rect 11793 19799 11851 19805
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 12986 19796 12992 19848
rect 13044 19836 13050 19848
rect 13633 19839 13691 19845
rect 13044 19808 13089 19836
rect 13044 19796 13050 19808
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13679 19808 13713 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 4494 19771 4552 19777
rect 4494 19768 4506 19771
rect 3936 19740 4506 19768
rect 3936 19728 3942 19740
rect 4494 19737 4506 19740
rect 4540 19737 4552 19771
rect 4494 19731 4552 19737
rect 4706 19728 4712 19780
rect 4764 19768 4770 19780
rect 9309 19771 9367 19777
rect 4764 19740 8892 19768
rect 4764 19728 4770 19740
rect 2222 19700 2228 19712
rect 2183 19672 2228 19700
rect 2222 19660 2228 19672
rect 2280 19660 2286 19712
rect 2590 19700 2596 19712
rect 2551 19672 2596 19700
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 2774 19660 2780 19712
rect 2832 19700 2838 19712
rect 2869 19703 2927 19709
rect 2869 19700 2881 19703
rect 2832 19672 2881 19700
rect 2832 19660 2838 19672
rect 2869 19669 2881 19672
rect 2915 19700 2927 19703
rect 3050 19700 3056 19712
rect 2915 19672 3056 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3200 19672 3801 19700
rect 3200 19660 3206 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 7248 19672 7573 19700
rect 7248 19660 7254 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7561 19663 7619 19669
rect 7929 19703 7987 19709
rect 7929 19669 7941 19703
rect 7975 19700 7987 19703
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7975 19672 8309 19700
rect 7975 19669 7987 19672
rect 7929 19663 7987 19669
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 8297 19663 8355 19669
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 8754 19700 8760 19712
rect 8444 19672 8489 19700
rect 8715 19672 8760 19700
rect 8444 19660 8450 19672
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 8864 19700 8892 19740
rect 9309 19737 9321 19771
rect 9355 19768 9367 19771
rect 10502 19768 10508 19780
rect 9355 19740 10508 19768
rect 9355 19737 9367 19740
rect 9309 19731 9367 19737
rect 10502 19728 10508 19740
rect 10560 19728 10566 19780
rect 10594 19728 10600 19780
rect 10652 19728 10658 19780
rect 10778 19777 10784 19780
rect 10720 19771 10784 19777
rect 10720 19737 10732 19771
rect 10766 19737 10784 19771
rect 10720 19731 10784 19737
rect 10778 19728 10784 19731
rect 10836 19728 10842 19780
rect 12066 19768 12072 19780
rect 10888 19740 12072 19768
rect 10888 19700 10916 19740
rect 12066 19728 12072 19740
rect 12124 19728 12130 19780
rect 12621 19771 12679 19777
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 13170 19768 13176 19780
rect 12667 19740 13176 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 13170 19728 13176 19740
rect 13228 19728 13234 19780
rect 13648 19768 13676 19799
rect 14274 19796 14280 19848
rect 14332 19836 14338 19848
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 14332 19808 14381 19836
rect 14332 19796 14338 19808
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14734 19836 14740 19848
rect 14695 19808 14740 19836
rect 14369 19799 14427 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 15102 19836 15108 19848
rect 15063 19808 15108 19836
rect 15102 19796 15108 19808
rect 15160 19796 15166 19848
rect 15194 19796 15200 19848
rect 15252 19836 15258 19848
rect 15252 19808 15297 19836
rect 15252 19796 15258 19808
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15565 19839 15623 19845
rect 15565 19836 15577 19839
rect 15528 19808 15577 19836
rect 15528 19796 15534 19808
rect 15565 19805 15577 19808
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 13725 19771 13783 19777
rect 13725 19768 13737 19771
rect 13280 19740 13737 19768
rect 11698 19700 11704 19712
rect 8864 19672 10916 19700
rect 11659 19672 11704 19700
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 13280 19700 13308 19740
rect 13725 19737 13737 19740
rect 13771 19737 13783 19771
rect 15580 19768 15608 19799
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15712 19808 15945 19836
rect 15712 19796 15718 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 16758 19836 16764 19848
rect 16719 19808 16764 19836
rect 15933 19799 15991 19805
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17586 19836 17592 19848
rect 17547 19808 17592 19836
rect 17037 19799 17095 19805
rect 17052 19768 17080 19799
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 18598 19836 18604 19848
rect 18187 19808 18604 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 18598 19796 18604 19808
rect 18656 19796 18662 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18966 19836 18972 19848
rect 18739 19808 18972 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18966 19796 18972 19808
rect 19024 19836 19030 19848
rect 19076 19836 19104 20003
rect 20806 20000 20812 20012
rect 20864 20040 20870 20052
rect 21453 20043 21511 20049
rect 21453 20040 21465 20043
rect 20864 20012 21465 20040
rect 20864 20000 20870 20012
rect 21453 20009 21465 20012
rect 21499 20040 21511 20043
rect 21542 20040 21548 20052
rect 21499 20012 21548 20040
rect 21499 20009 21511 20012
rect 21453 20003 21511 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 19610 19904 19616 19916
rect 19571 19876 19616 19904
rect 19610 19864 19616 19876
rect 19668 19864 19674 19916
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 21085 19907 21143 19913
rect 21085 19904 21097 19907
rect 20680 19876 21097 19904
rect 20680 19864 20686 19876
rect 21085 19873 21097 19876
rect 21131 19873 21143 19907
rect 21085 19867 21143 19873
rect 19024 19808 19104 19836
rect 19024 19796 19030 19808
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19852 19808 20085 19836
rect 19852 19796 19858 19808
rect 20073 19805 20085 19808
rect 20119 19805 20131 19839
rect 20073 19799 20131 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20438 19836 20444 19848
rect 20395 19808 20444 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 18506 19768 18512 19780
rect 15580 19740 15976 19768
rect 17052 19740 18512 19768
rect 13725 19731 13783 19737
rect 15948 19712 15976 19740
rect 18506 19728 18512 19740
rect 18564 19728 18570 19780
rect 20162 19728 20168 19780
rect 20220 19768 20226 19780
rect 20916 19768 20944 19799
rect 20220 19740 20944 19768
rect 20220 19728 20226 19740
rect 11848 19672 13308 19700
rect 11848 19660 11854 19672
rect 15930 19660 15936 19712
rect 15988 19660 15994 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 3326 19496 3332 19508
rect 2700 19468 3332 19496
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 2700 19437 2728 19468
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 3878 19496 3884 19508
rect 3839 19468 3884 19496
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 4706 19456 4712 19508
rect 4764 19496 4770 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 4764 19468 5365 19496
rect 4764 19456 4770 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5810 19496 5816 19508
rect 5771 19468 5816 19496
rect 5353 19459 5411 19465
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6512 19468 6837 19496
rect 6512 19456 6518 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 7190 19496 7196 19508
rect 7151 19468 7196 19496
rect 6825 19459 6883 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 7466 19456 7472 19508
rect 7524 19456 7530 19508
rect 8662 19496 8668 19508
rect 8623 19468 8668 19496
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 10229 19499 10287 19505
rect 10229 19465 10241 19499
rect 10275 19496 10287 19499
rect 10410 19496 10416 19508
rect 10275 19468 10416 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 11238 19496 11244 19508
rect 11199 19468 11244 19496
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 13814 19496 13820 19508
rect 13403 19468 13820 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15289 19499 15347 19505
rect 15289 19496 15301 19499
rect 15252 19468 15301 19496
rect 15252 19456 15258 19468
rect 15289 19465 15301 19468
rect 15335 19465 15347 19499
rect 15289 19459 15347 19465
rect 15933 19499 15991 19505
rect 15933 19465 15945 19499
rect 15979 19496 15991 19499
rect 16022 19496 16028 19508
rect 15979 19468 16028 19496
rect 15979 19465 15991 19468
rect 15933 19459 15991 19465
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 16390 19456 16396 19508
rect 16448 19496 16454 19508
rect 16761 19499 16819 19505
rect 16761 19496 16773 19499
rect 16448 19468 16773 19496
rect 16448 19456 16454 19468
rect 16761 19465 16773 19468
rect 16807 19465 16819 19499
rect 16761 19459 16819 19465
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 17494 19496 17500 19508
rect 17267 19468 17500 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 17862 19496 17868 19508
rect 17823 19468 17868 19496
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18156 19468 18337 19496
rect 2685 19431 2743 19437
rect 2685 19428 2697 19431
rect 2096 19400 2697 19428
rect 2096 19388 2102 19400
rect 2685 19397 2697 19400
rect 2731 19397 2743 19431
rect 2685 19391 2743 19397
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 3200 19400 3464 19428
rect 3200 19388 3206 19400
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 2222 19360 2228 19372
rect 2179 19332 2228 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 2590 19360 2596 19372
rect 2547 19332 2596 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 2590 19320 2596 19332
rect 2648 19360 2654 19372
rect 2866 19360 2872 19372
rect 2648 19332 2872 19360
rect 2648 19320 2654 19332
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 3050 19320 3056 19372
rect 3108 19360 3114 19372
rect 3237 19363 3295 19369
rect 3237 19360 3249 19363
rect 3108 19332 3249 19360
rect 3108 19320 3114 19332
rect 3237 19329 3249 19332
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3436 19301 3464 19400
rect 6564 19400 6776 19428
rect 4154 19360 4160 19372
rect 4080 19332 4160 19360
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19261 3479 19295
rect 3421 19255 3479 19261
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 4080 19292 4108 19332
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 5005 19363 5063 19369
rect 5005 19329 5017 19363
rect 5051 19360 5063 19363
rect 5166 19360 5172 19372
rect 5051 19332 5172 19360
rect 5051 19329 5063 19332
rect 5005 19323 5063 19329
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 5258 19320 5264 19372
rect 5316 19369 5322 19372
rect 5316 19363 5330 19369
rect 5318 19360 5330 19363
rect 5318 19332 5361 19360
rect 5318 19329 5330 19332
rect 5316 19323 5330 19329
rect 5316 19320 5322 19323
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 5721 19363 5779 19369
rect 5721 19360 5733 19363
rect 5500 19332 5733 19360
rect 5500 19320 5506 19332
rect 5721 19329 5733 19332
rect 5767 19360 5779 19363
rect 6564 19360 6592 19400
rect 5767 19332 6592 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 5902 19292 5908 19304
rect 3835 19264 4108 19292
rect 5863 19264 5908 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6748 19301 6776 19400
rect 7190 19320 7196 19372
rect 7248 19360 7254 19372
rect 7484 19360 7512 19456
rect 7552 19431 7610 19437
rect 7552 19397 7564 19431
rect 7598 19428 7610 19431
rect 7742 19428 7748 19440
rect 7598 19400 7748 19428
rect 7598 19397 7610 19400
rect 7552 19391 7610 19397
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 8680 19360 8708 19456
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 10689 19431 10747 19437
rect 10689 19428 10701 19431
rect 8812 19400 10701 19428
rect 8812 19388 8818 19400
rect 10689 19397 10701 19400
rect 10735 19397 10747 19431
rect 10689 19391 10747 19397
rect 10962 19388 10968 19440
rect 11020 19428 11026 19440
rect 11762 19431 11820 19437
rect 11762 19428 11774 19431
rect 11020 19400 11774 19428
rect 11020 19388 11026 19400
rect 11762 19397 11774 19400
rect 11808 19397 11820 19431
rect 11762 19391 11820 19397
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 14458 19428 14464 19440
rect 13780 19400 14320 19428
rect 14419 19400 14464 19428
rect 13780 19388 13786 19400
rect 9013 19363 9071 19369
rect 9013 19360 9025 19363
rect 7248 19332 8524 19360
rect 8680 19332 9025 19360
rect 7248 19320 7254 19332
rect 7300 19301 7328 19332
rect 8496 19304 8524 19332
rect 9013 19329 9025 19332
rect 9059 19329 9071 19363
rect 10594 19360 10600 19372
rect 10555 19332 10600 19360
rect 9013 19323 9071 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 10870 19320 10876 19372
rect 10928 19360 10934 19372
rect 11057 19363 11115 19369
rect 11057 19360 11069 19363
rect 10928 19332 11069 19360
rect 10928 19320 10934 19332
rect 11057 19329 11069 19332
rect 11103 19329 11115 19363
rect 11057 19323 11115 19329
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11296 19332 11529 19360
rect 11296 19320 11302 19332
rect 11517 19329 11529 19332
rect 11563 19360 11575 19363
rect 13170 19360 13176 19372
rect 11563 19332 12572 19360
rect 13131 19332 13176 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 6641 19255 6699 19261
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 7285 19295 7343 19301
rect 6779 19264 7236 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 2406 19184 2412 19236
rect 2464 19224 2470 19236
rect 2464 19196 3197 19224
rect 2464 19184 2470 19196
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3169 19156 3197 19196
rect 3234 19184 3240 19236
rect 3292 19224 3298 19236
rect 5534 19224 5540 19236
rect 3292 19196 4384 19224
rect 3292 19184 3298 19196
rect 4154 19156 4160 19168
rect 2924 19128 2969 19156
rect 3169 19128 4160 19156
rect 2924 19116 2930 19128
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 4356 19156 4384 19196
rect 5276 19196 5540 19224
rect 5276 19156 5304 19196
rect 5534 19184 5540 19196
rect 5592 19224 5598 19236
rect 5994 19224 6000 19236
rect 5592 19196 6000 19224
rect 5592 19184 5598 19196
rect 5994 19184 6000 19196
rect 6052 19224 6058 19236
rect 6362 19224 6368 19236
rect 6052 19196 6368 19224
rect 6052 19184 6058 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 6656 19224 6684 19255
rect 7098 19224 7104 19236
rect 6656 19196 7104 19224
rect 7098 19184 7104 19196
rect 7156 19184 7162 19236
rect 4356 19128 5304 19156
rect 7208 19156 7236 19264
rect 7285 19261 7297 19295
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 8536 19264 8769 19292
rect 8536 19252 8542 19264
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 12544 19292 12572 19332
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14185 19363 14243 19369
rect 14185 19360 14197 19363
rect 13872 19332 14197 19360
rect 13872 19320 13878 19332
rect 14185 19329 14197 19332
rect 14231 19329 14243 19363
rect 14292 19360 14320 19400
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15013 19431 15071 19437
rect 15013 19397 15025 19431
rect 15059 19428 15071 19431
rect 15654 19428 15660 19440
rect 15059 19400 15660 19428
rect 15059 19397 15071 19400
rect 15013 19391 15071 19397
rect 15654 19388 15660 19400
rect 15712 19388 15718 19440
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 18156 19428 18184 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18506 19496 18512 19508
rect 18467 19468 18512 19496
rect 18325 19459 18383 19465
rect 18506 19456 18512 19468
rect 18564 19496 18570 19508
rect 18564 19468 20576 19496
rect 18564 19456 18570 19468
rect 17644 19400 18184 19428
rect 17644 19388 17650 19400
rect 18230 19388 18236 19440
rect 18288 19428 18294 19440
rect 19061 19431 19119 19437
rect 19061 19428 19073 19431
rect 18288 19400 19073 19428
rect 18288 19388 18294 19400
rect 19061 19397 19073 19400
rect 19107 19397 19119 19431
rect 19702 19428 19708 19440
rect 19663 19400 19708 19428
rect 19061 19391 19119 19397
rect 19702 19388 19708 19400
rect 19760 19388 19766 19440
rect 20254 19428 20260 19440
rect 20215 19400 20260 19428
rect 20254 19388 20260 19400
rect 20312 19388 20318 19440
rect 20548 19372 20576 19468
rect 20809 19431 20867 19437
rect 20809 19397 20821 19431
rect 20855 19428 20867 19431
rect 21174 19428 21180 19440
rect 20855 19400 21180 19428
rect 20855 19397 20867 19400
rect 20809 19391 20867 19397
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 21361 19431 21419 19437
rect 21361 19397 21373 19431
rect 21407 19428 21419 19431
rect 21450 19428 21456 19440
rect 21407 19400 21456 19428
rect 21407 19397 21419 19400
rect 21361 19391 21419 19397
rect 21450 19388 21456 19400
rect 21508 19388 21514 19440
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14292 19332 14749 19360
rect 14185 19323 14243 19329
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 15749 19363 15807 19369
rect 15749 19360 15761 19363
rect 14737 19323 14795 19329
rect 15672 19332 15761 19360
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 10836 19264 10929 19292
rect 12544 19264 13001 19292
rect 10836 19252 10842 19264
rect 12989 19261 13001 19264
rect 13035 19292 13047 19295
rect 13078 19292 13084 19304
rect 13035 19264 13084 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 10137 19227 10195 19233
rect 10137 19193 10149 19227
rect 10183 19224 10195 19227
rect 10796 19224 10824 19252
rect 10183 19196 10824 19224
rect 12897 19227 12955 19233
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 12897 19193 12909 19227
rect 12943 19224 12955 19227
rect 13538 19224 13544 19236
rect 12943 19196 13544 19224
rect 12943 19193 12955 19196
rect 12897 19187 12955 19193
rect 13538 19184 13544 19196
rect 13596 19184 13602 19236
rect 15672 19168 15700 19332
rect 15749 19329 15761 19332
rect 15795 19329 15807 19363
rect 16942 19360 16948 19372
rect 16903 19332 16948 19360
rect 15749 19323 15807 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 17405 19363 17463 19369
rect 17405 19360 17417 19363
rect 17092 19332 17417 19360
rect 17092 19320 17098 19332
rect 17405 19329 17417 19332
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 19334 19360 19340 19372
rect 19295 19332 19340 19360
rect 18049 19323 18107 19329
rect 16482 19292 16488 19304
rect 16395 19264 16488 19292
rect 16482 19252 16488 19264
rect 16540 19292 16546 19304
rect 16960 19292 16988 19320
rect 18064 19292 18092 19323
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 20438 19360 20444 19372
rect 20027 19332 20444 19360
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 16540 19264 16988 19292
rect 17604 19264 18092 19292
rect 16540 19252 16546 19264
rect 17604 19168 17632 19264
rect 18598 19252 18604 19304
rect 18656 19292 18662 19304
rect 19058 19292 19064 19304
rect 18656 19264 19064 19292
rect 18656 19252 18662 19264
rect 19058 19252 19064 19264
rect 19116 19292 19122 19304
rect 19444 19292 19472 19323
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20588 19332 20681 19360
rect 20732 19332 21097 19360
rect 20588 19320 20594 19332
rect 19116 19264 19472 19292
rect 19116 19252 19122 19264
rect 19886 19252 19892 19304
rect 19944 19292 19950 19304
rect 20732 19292 20760 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 19944 19264 20760 19292
rect 19944 19252 19950 19264
rect 8018 19156 8024 19168
rect 7208 19128 8024 19156
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 12802 19156 12808 19168
rect 8352 19128 12808 19156
rect 8352 19116 8358 19128
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 13688 19128 13921 19156
rect 13688 19116 13694 19128
rect 13909 19125 13921 19128
rect 13955 19156 13967 19159
rect 14366 19156 14372 19168
rect 13955 19128 14372 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 15654 19156 15660 19168
rect 15615 19128 15660 19156
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 17586 19156 17592 19168
rect 17547 19128 17592 19156
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 18782 19156 18788 19168
rect 18743 19128 18788 19156
rect 18782 19116 18788 19128
rect 18840 19156 18846 19168
rect 19334 19156 19340 19168
rect 18840 19128 19340 19156
rect 18840 19116 18846 19128
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 4249 18955 4307 18961
rect 4249 18952 4261 18955
rect 3384 18924 4261 18952
rect 3384 18912 3390 18924
rect 4249 18921 4261 18924
rect 4295 18952 4307 18955
rect 4798 18952 4804 18964
rect 4295 18924 4804 18952
rect 4295 18921 4307 18924
rect 4249 18915 4307 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 5169 18955 5227 18961
rect 5169 18952 5181 18955
rect 5092 18924 5181 18952
rect 3142 18884 3148 18896
rect 2056 18856 3148 18884
rect 2056 18825 2084 18856
rect 3142 18844 3148 18856
rect 3200 18884 3206 18896
rect 3602 18884 3608 18896
rect 3200 18856 3608 18884
rect 3200 18844 3206 18856
rect 3602 18844 3608 18856
rect 3660 18844 3666 18896
rect 4154 18884 4160 18896
rect 4115 18856 4160 18884
rect 4154 18844 4160 18856
rect 4212 18844 4218 18896
rect 4890 18844 4896 18896
rect 4948 18884 4954 18896
rect 5092 18884 5120 18924
rect 5169 18921 5181 18924
rect 5215 18921 5227 18955
rect 7190 18952 7196 18964
rect 5169 18915 5227 18921
rect 6932 18924 7196 18952
rect 4948 18856 5120 18884
rect 4948 18844 4954 18856
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 2832 18788 2877 18816
rect 2832 18776 2838 18788
rect 2958 18776 2964 18828
rect 3016 18816 3022 18828
rect 3881 18819 3939 18825
rect 3881 18816 3893 18819
rect 3016 18788 3893 18816
rect 3016 18776 3022 18788
rect 3881 18785 3893 18788
rect 3927 18816 3939 18819
rect 4522 18816 4528 18828
rect 3927 18788 4528 18816
rect 3927 18785 3939 18788
rect 3881 18779 3939 18785
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 2130 18748 2136 18760
rect 1811 18720 2136 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2866 18708 2872 18760
rect 2924 18748 2930 18760
rect 3053 18751 3111 18757
rect 3053 18748 3065 18751
rect 2924 18720 3065 18748
rect 2924 18708 2930 18720
rect 3053 18717 3065 18720
rect 3099 18717 3111 18751
rect 4632 18748 4660 18779
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 5534 18816 5540 18828
rect 4764 18788 4809 18816
rect 5184 18788 5540 18816
rect 4764 18776 4770 18788
rect 5184 18748 5212 18788
rect 5534 18776 5540 18788
rect 5592 18776 5598 18828
rect 5718 18816 5724 18828
rect 5679 18788 5724 18816
rect 5718 18776 5724 18788
rect 5776 18776 5782 18828
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 5902 18816 5908 18828
rect 5859 18788 5908 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 4632 18720 5212 18748
rect 3053 18711 3111 18717
rect 3234 18680 3240 18692
rect 2148 18652 3240 18680
rect 2148 18621 2176 18652
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 4801 18683 4859 18689
rect 4801 18649 4813 18683
rect 4847 18680 4859 18683
rect 4847 18652 5304 18680
rect 4847 18649 4859 18652
rect 4801 18643 4859 18649
rect 2133 18615 2191 18621
rect 2133 18612 2145 18615
rect 1044 18584 2145 18612
rect 566 18368 572 18420
rect 624 18408 630 18420
rect 1044 18408 1072 18584
rect 2133 18581 2145 18584
rect 2179 18581 2191 18615
rect 2133 18575 2191 18581
rect 2225 18615 2283 18621
rect 2225 18581 2237 18615
rect 2271 18612 2283 18615
rect 2314 18612 2320 18624
rect 2271 18584 2320 18612
rect 2271 18581 2283 18584
rect 2225 18575 2283 18581
rect 2314 18572 2320 18584
rect 2372 18572 2378 18624
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2639 18584 2973 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2961 18581 2973 18584
rect 3007 18581 3019 18615
rect 2961 18575 3019 18581
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3421 18615 3479 18621
rect 3421 18612 3433 18615
rect 3384 18584 3433 18612
rect 3384 18572 3390 18584
rect 3421 18581 3433 18584
rect 3467 18581 3479 18615
rect 3602 18612 3608 18624
rect 3563 18584 3608 18612
rect 3421 18575 3479 18581
rect 3602 18572 3608 18584
rect 3660 18572 3666 18624
rect 5276 18621 5304 18652
rect 5350 18640 5356 18692
rect 5408 18680 5414 18692
rect 5828 18680 5856 18779
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6362 18816 6368 18828
rect 6323 18788 6368 18816
rect 6181 18779 6239 18785
rect 6196 18748 6224 18779
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 6932 18825 6960 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 7340 18924 8309 18952
rect 7340 18912 7346 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 8297 18915 8355 18921
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 8536 18924 8769 18952
rect 8536 18912 8542 18924
rect 8757 18921 8769 18924
rect 8803 18952 8815 18955
rect 9582 18952 9588 18964
rect 8803 18924 9588 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 10594 18952 10600 18964
rect 9723 18924 10600 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 10689 18955 10747 18961
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 10962 18952 10968 18964
rect 10735 18924 10968 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11790 18952 11796 18964
rect 11072 18924 11796 18952
rect 8018 18844 8024 18896
rect 8076 18884 8082 18896
rect 11072 18884 11100 18924
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 12894 18912 12900 18964
rect 12952 18952 12958 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12952 18924 13001 18952
rect 12952 18912 12958 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 18966 18952 18972 18964
rect 18927 18924 18972 18952
rect 12989 18915 13047 18921
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 19058 18912 19064 18964
rect 19116 18952 19122 18964
rect 19337 18955 19395 18961
rect 19337 18952 19349 18955
rect 19116 18924 19349 18952
rect 19116 18912 19122 18924
rect 19337 18921 19349 18924
rect 19383 18921 19395 18955
rect 21358 18952 21364 18964
rect 21319 18924 21364 18952
rect 19337 18915 19395 18921
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 13078 18884 13084 18896
rect 8076 18856 11100 18884
rect 12084 18856 13084 18884
rect 8076 18844 8082 18856
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18785 6975 18819
rect 6917 18779 6975 18785
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8720 18788 9045 18816
rect 8720 18776 8726 18788
rect 9033 18785 9045 18788
rect 9079 18785 9091 18819
rect 9033 18779 9091 18785
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 10870 18816 10876 18828
rect 10091 18788 10876 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 12084 18825 12112 18856
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 20714 18884 20720 18896
rect 16592 18856 20720 18884
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18785 12127 18819
rect 12802 18816 12808 18828
rect 12763 18788 12808 18816
rect 12069 18779 12127 18785
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 13538 18816 13544 18828
rect 13499 18788 13544 18816
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 14182 18816 14188 18828
rect 14143 18788 14188 18816
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14366 18816 14372 18828
rect 14327 18788 14372 18816
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 16592 18816 16620 18856
rect 20714 18844 20720 18856
rect 20772 18884 20778 18896
rect 20772 18856 21220 18884
rect 20772 18844 20778 18856
rect 15620 18788 16620 18816
rect 18877 18819 18935 18825
rect 15620 18776 15626 18788
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 18923 18788 20484 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 20456 18760 20484 18788
rect 7006 18748 7012 18760
rect 6196 18720 7012 18748
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7184 18751 7242 18757
rect 7184 18717 7196 18751
rect 7230 18717 7242 18751
rect 7184 18711 7242 18717
rect 6454 18680 6460 18692
rect 5408 18652 5856 18680
rect 6415 18652 6460 18680
rect 5408 18640 5414 18652
rect 6454 18640 6460 18652
rect 6512 18640 6518 18692
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18581 5319 18615
rect 5261 18575 5319 18581
rect 5629 18615 5687 18621
rect 5629 18581 5641 18615
rect 5675 18612 5687 18615
rect 5718 18612 5724 18624
rect 5675 18584 5724 18612
rect 5675 18581 5687 18584
rect 5629 18575 5687 18581
rect 5718 18572 5724 18584
rect 5776 18612 5782 18624
rect 5902 18612 5908 18624
rect 5776 18584 5908 18612
rect 5776 18572 5782 18584
rect 5902 18572 5908 18584
rect 5960 18572 5966 18624
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7024 18612 7052 18708
rect 7098 18640 7104 18692
rect 7156 18680 7162 18692
rect 7208 18680 7236 18711
rect 8018 18708 8024 18760
rect 8076 18748 8082 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 8076 18720 9781 18748
rect 8076 18708 8082 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 13817 18751 13875 18757
rect 13817 18748 13829 18751
rect 9769 18711 9827 18717
rect 9876 18720 13829 18748
rect 7156 18652 7236 18680
rect 7156 18640 7162 18652
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 9876 18680 9904 18720
rect 13817 18717 13829 18720
rect 13863 18748 13875 18751
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 13863 18720 14473 18748
rect 13863 18717 13875 18720
rect 13817 18711 13875 18717
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19024 18720 19533 18748
rect 19024 18708 19030 18720
rect 19521 18717 19533 18720
rect 19567 18748 19579 18751
rect 20073 18751 20131 18757
rect 20073 18748 20085 18751
rect 19567 18720 20085 18748
rect 19567 18717 19579 18720
rect 19521 18711 19579 18717
rect 20073 18717 20085 18720
rect 20119 18717 20131 18751
rect 20346 18748 20352 18760
rect 20307 18720 20352 18748
rect 20073 18711 20131 18717
rect 20346 18708 20352 18720
rect 20404 18708 20410 18760
rect 20438 18708 20444 18760
rect 20496 18748 20502 18760
rect 21192 18757 21220 18856
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20496 18720 20637 18748
rect 20496 18708 20502 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 21177 18751 21235 18757
rect 21177 18717 21189 18751
rect 21223 18748 21235 18751
rect 21266 18748 21272 18760
rect 21223 18720 21272 18748
rect 21223 18717 21235 18720
rect 21177 18711 21235 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 7524 18652 9904 18680
rect 7524 18640 7530 18652
rect 11698 18640 11704 18692
rect 11756 18680 11762 18692
rect 11802 18683 11860 18689
rect 11802 18680 11814 18683
rect 11756 18652 11814 18680
rect 11756 18640 11762 18652
rect 11802 18649 11814 18652
rect 11848 18649 11860 18683
rect 11802 18643 11860 18649
rect 11974 18640 11980 18692
rect 12032 18680 12038 18692
rect 13449 18683 13507 18689
rect 13449 18680 13461 18683
rect 12032 18652 13461 18680
rect 12032 18640 12038 18652
rect 13449 18649 13461 18652
rect 13495 18649 13507 18683
rect 13449 18643 13507 18649
rect 19797 18683 19855 18689
rect 19797 18649 19809 18683
rect 19843 18649 19855 18683
rect 19797 18643 19855 18649
rect 20901 18683 20959 18689
rect 20901 18649 20913 18683
rect 20947 18680 20959 18683
rect 20990 18680 20996 18692
rect 20947 18652 20996 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 7374 18612 7380 18624
rect 7024 18584 7380 18612
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 9088 18584 9229 18612
rect 9088 18572 9094 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9364 18584 9409 18612
rect 9364 18572 9370 18584
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 10321 18615 10379 18621
rect 10321 18612 10333 18615
rect 9732 18584 10333 18612
rect 9732 18572 9738 18584
rect 10321 18581 10333 18584
rect 10367 18612 10379 18615
rect 10686 18612 10692 18624
rect 10367 18584 10692 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 12161 18615 12219 18621
rect 12161 18612 12173 18615
rect 10928 18584 12173 18612
rect 10928 18572 10934 18584
rect 12161 18581 12173 18584
rect 12207 18581 12219 18615
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12161 18575 12219 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13354 18612 13360 18624
rect 12676 18584 12721 18612
rect 13315 18584 13360 18612
rect 12676 18572 12682 18584
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 14829 18615 14887 18621
rect 14829 18581 14841 18615
rect 14875 18612 14887 18615
rect 15746 18612 15752 18624
rect 14875 18584 15752 18612
rect 14875 18581 14887 18584
rect 14829 18575 14887 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 19812 18612 19840 18643
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 22278 18612 22284 18624
rect 19812 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1673 18411 1731 18417
rect 1673 18408 1685 18411
rect 624 18380 1685 18408
rect 624 18368 630 18380
rect 1673 18377 1685 18380
rect 1719 18377 1731 18411
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1673 18371 1731 18377
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2314 18368 2320 18420
rect 2372 18368 2378 18420
rect 4341 18411 4399 18417
rect 4341 18377 4353 18411
rect 4387 18408 4399 18411
rect 7377 18411 7435 18417
rect 4387 18380 7144 18408
rect 4387 18377 4399 18380
rect 4341 18371 4399 18377
rect 1302 18300 1308 18352
rect 1360 18340 1366 18352
rect 1489 18343 1547 18349
rect 1489 18340 1501 18343
rect 1360 18312 1501 18340
rect 1360 18300 1366 18312
rect 1489 18309 1501 18312
rect 1535 18340 1547 18343
rect 2332 18340 2360 18368
rect 1535 18312 2360 18340
rect 1535 18309 1547 18312
rect 1489 18303 1547 18309
rect 3050 18300 3056 18352
rect 3108 18340 3114 18352
rect 3108 18312 5396 18340
rect 3108 18300 3114 18312
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2314 18272 2320 18284
rect 2179 18244 2320 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 3142 18272 3148 18284
rect 3103 18244 3148 18272
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 3973 18275 4031 18281
rect 3973 18241 3985 18275
rect 4019 18272 4031 18275
rect 5258 18272 5264 18284
rect 4019 18244 5264 18272
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 5368 18272 5396 18312
rect 5534 18300 5540 18352
rect 5592 18349 5598 18352
rect 5592 18340 5604 18349
rect 6181 18343 6239 18349
rect 6181 18340 6193 18343
rect 5592 18312 5637 18340
rect 5828 18312 6193 18340
rect 5592 18303 5604 18312
rect 5592 18300 5598 18303
rect 5828 18272 5856 18312
rect 6181 18309 6193 18312
rect 6227 18340 6239 18343
rect 7116 18340 7144 18380
rect 7377 18377 7389 18411
rect 7423 18408 7435 18411
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7423 18380 7757 18408
rect 7423 18377 7435 18380
rect 7377 18371 7435 18377
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8386 18408 8392 18420
rect 8251 18380 8392 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8386 18368 8392 18380
rect 8444 18368 8450 18420
rect 8665 18411 8723 18417
rect 8665 18377 8677 18411
rect 8711 18408 8723 18411
rect 9125 18411 9183 18417
rect 9125 18408 9137 18411
rect 8711 18380 9137 18408
rect 8711 18377 8723 18380
rect 8665 18371 8723 18377
rect 9125 18377 9137 18380
rect 9171 18377 9183 18411
rect 10042 18408 10048 18420
rect 9125 18371 9183 18377
rect 9646 18380 10048 18408
rect 8018 18340 8024 18352
rect 6227 18312 7052 18340
rect 7116 18312 8024 18340
rect 6227 18309 6239 18312
rect 6181 18303 6239 18309
rect 5368 18244 5856 18272
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 5960 18244 6500 18272
rect 5960 18232 5966 18244
rect 2866 18204 2872 18216
rect 2827 18176 2872 18204
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 3050 18204 3056 18216
rect 3011 18176 3056 18204
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3786 18204 3792 18216
rect 3747 18176 3792 18204
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 4522 18204 4528 18216
rect 3927 18176 4528 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 5859 18176 6040 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 3513 18139 3571 18145
rect 3513 18105 3525 18139
rect 3559 18136 3571 18139
rect 3970 18136 3976 18148
rect 3559 18108 3976 18136
rect 3559 18105 3571 18108
rect 3513 18099 3571 18105
rect 3970 18096 3976 18108
rect 4028 18096 4034 18148
rect 4706 18136 4712 18148
rect 4080 18108 4712 18136
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2225 18071 2283 18077
rect 2225 18068 2237 18071
rect 2188 18040 2237 18068
rect 2188 18028 2194 18040
rect 2225 18037 2237 18040
rect 2271 18037 2283 18071
rect 2225 18031 2283 18037
rect 3602 18028 3608 18080
rect 3660 18068 3666 18080
rect 4080 18068 4108 18108
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 3660 18040 4108 18068
rect 4433 18071 4491 18077
rect 3660 18028 3666 18040
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 5166 18068 5172 18080
rect 4479 18040 5172 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 6012 18077 6040 18176
rect 6472 18136 6500 18244
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6730 18272 6736 18284
rect 6604 18244 6736 18272
rect 6604 18232 6610 18244
rect 6730 18232 6736 18244
rect 6788 18272 6794 18284
rect 7024 18281 7052 18312
rect 8018 18300 8024 18312
rect 8076 18300 8082 18352
rect 9493 18343 9551 18349
rect 9493 18309 9505 18343
rect 9539 18340 9551 18343
rect 9646 18340 9674 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 10870 18408 10876 18420
rect 10831 18380 10876 18408
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 10965 18411 11023 18417
rect 10965 18377 10977 18411
rect 11011 18408 11023 18411
rect 11885 18411 11943 18417
rect 11885 18408 11897 18411
rect 11011 18380 11897 18408
rect 11011 18377 11023 18380
rect 10965 18371 11023 18377
rect 11885 18377 11897 18380
rect 11931 18377 11943 18411
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 11885 18371 11943 18377
rect 12250 18368 12256 18380
rect 12308 18408 12314 18420
rect 12308 18380 14136 18408
rect 12308 18368 12314 18380
rect 9539 18312 9674 18340
rect 9539 18309 9551 18312
rect 9493 18303 9551 18309
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 13078 18340 13084 18352
rect 11756 18312 12572 18340
rect 13039 18312 13084 18340
rect 11756 18300 11762 18312
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6788 18244 6929 18272
rect 6788 18232 6794 18244
rect 6917 18241 6929 18244
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7466 18272 7472 18284
rect 7055 18244 7472 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18272 7895 18275
rect 8478 18272 8484 18284
rect 7883 18244 8484 18272
rect 7883 18241 7895 18244
rect 7837 18235 7895 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9600 18244 10149 18272
rect 9600 18216 9628 18244
rect 10137 18241 10149 18244
rect 10183 18272 10195 18275
rect 12158 18272 12164 18284
rect 10183 18244 12164 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12544 18272 12572 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 13440 18343 13498 18349
rect 13440 18309 13452 18343
rect 13486 18340 13498 18343
rect 13538 18340 13544 18352
rect 13486 18312 13544 18340
rect 13486 18309 13498 18312
rect 13440 18303 13498 18309
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 14108 18340 14136 18380
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14458 18408 14464 18420
rect 14240 18380 14464 18408
rect 14240 18368 14246 18380
rect 14458 18368 14464 18380
rect 14516 18408 14522 18420
rect 14553 18411 14611 18417
rect 14553 18408 14565 18411
rect 14516 18380 14565 18408
rect 14516 18368 14522 18380
rect 14553 18377 14565 18380
rect 14599 18377 14611 18411
rect 15562 18408 15568 18420
rect 15523 18380 15568 18408
rect 14553 18371 14611 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 19794 18408 19800 18420
rect 19755 18380 19800 18408
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 20530 18408 20536 18420
rect 20491 18380 20536 18408
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 21450 18408 21456 18420
rect 21411 18380 21456 18408
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 17034 18340 17040 18352
rect 14108 18312 17040 18340
rect 17034 18300 17040 18312
rect 17092 18340 17098 18352
rect 18322 18340 18328 18352
rect 17092 18312 18328 18340
rect 17092 18300 17098 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 20548 18340 20576 18368
rect 19996 18312 20576 18340
rect 20993 18343 21051 18349
rect 12802 18272 12808 18284
rect 12544 18244 12808 18272
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7098 18204 7104 18216
rect 6871 18176 7104 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 7340 18176 7573 18204
rect 7340 18164 7346 18176
rect 7561 18173 7573 18176
rect 7607 18204 7619 18207
rect 8294 18204 8300 18216
rect 7607 18176 8300 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 8294 18164 8300 18176
rect 8352 18204 8358 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 8352 18176 8401 18204
rect 8352 18164 8358 18176
rect 8389 18173 8401 18176
rect 8435 18173 8447 18207
rect 8389 18167 8447 18173
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8662 18204 8668 18216
rect 8619 18176 8668 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18173 9735 18207
rect 9677 18167 9735 18173
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 10962 18204 10968 18216
rect 10827 18176 10968 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 6730 18136 6736 18148
rect 6472 18108 6736 18136
rect 6730 18096 6736 18108
rect 6788 18096 6794 18148
rect 5997 18071 6055 18077
rect 5997 18037 6009 18071
rect 6043 18068 6055 18071
rect 7006 18068 7012 18080
rect 6043 18040 7012 18068
rect 6043 18037 6055 18040
rect 5997 18031 6055 18037
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 7116 18068 7144 18164
rect 9030 18136 9036 18148
rect 8991 18108 9036 18136
rect 9030 18096 9036 18108
rect 9088 18096 9094 18148
rect 9490 18096 9496 18148
rect 9548 18136 9554 18148
rect 9692 18136 9720 18167
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 11609 18207 11667 18213
rect 11609 18173 11621 18207
rect 11655 18204 11667 18207
rect 11882 18204 11888 18216
rect 11655 18176 11888 18204
rect 11655 18173 11667 18176
rect 11609 18167 11667 18173
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 12342 18204 12348 18216
rect 12303 18176 12348 18204
rect 12342 18164 12348 18176
rect 12400 18164 12406 18216
rect 12544 18213 12572 18244
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13096 18272 13124 18300
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 13096 18244 14657 18272
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18173 12587 18207
rect 12710 18204 12716 18216
rect 12671 18176 12716 18204
rect 12529 18167 12587 18173
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 13096 18204 13124 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 19518 18232 19524 18284
rect 19576 18272 19582 18284
rect 19996 18281 20024 18312
rect 20993 18309 21005 18343
rect 21039 18340 21051 18343
rect 21634 18340 21640 18352
rect 21039 18312 21640 18340
rect 21039 18309 21051 18312
rect 20993 18303 21051 18309
rect 21634 18300 21640 18312
rect 21692 18300 21698 18352
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19576 18244 19625 18272
rect 19576 18232 19582 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20717 18275 20775 18281
rect 20717 18272 20729 18275
rect 20496 18244 20729 18272
rect 20496 18232 20502 18244
rect 20717 18241 20729 18244
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 13096 18176 13185 18204
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20165 18207 20223 18213
rect 20165 18204 20177 18207
rect 20128 18176 20177 18204
rect 20128 18164 20134 18176
rect 20165 18173 20177 18176
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 9548 18108 9720 18136
rect 11333 18139 11391 18145
rect 9548 18096 9554 18108
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 11974 18136 11980 18148
rect 11379 18108 11980 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 11974 18096 11980 18108
rect 12032 18096 12038 18148
rect 19337 18139 19395 18145
rect 19337 18105 19349 18139
rect 19383 18136 19395 18139
rect 19794 18136 19800 18148
rect 19383 18108 19800 18136
rect 19383 18105 19395 18108
rect 19337 18099 19395 18105
rect 19794 18096 19800 18108
rect 19852 18136 19858 18148
rect 21284 18136 21312 18235
rect 19852 18108 21312 18136
rect 19852 18096 19858 18108
rect 8386 18068 8392 18080
rect 7116 18040 8392 18068
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11664 18040 11713 18068
rect 11664 18028 11670 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 11701 18031 11759 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1762 17864 1768 17876
rect 1723 17836 1768 17864
rect 1762 17824 1768 17836
rect 1820 17824 1826 17876
rect 4522 17864 4528 17876
rect 4483 17836 4528 17864
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 5258 17824 5264 17876
rect 5316 17864 5322 17876
rect 5353 17867 5411 17873
rect 5353 17864 5365 17867
rect 5316 17836 5365 17864
rect 5316 17824 5322 17836
rect 5353 17833 5365 17836
rect 5399 17833 5411 17867
rect 5353 17827 5411 17833
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5902 17864 5908 17876
rect 5592 17836 5908 17864
rect 5592 17824 5598 17836
rect 5902 17824 5908 17836
rect 5960 17824 5966 17876
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 6181 17867 6239 17873
rect 6181 17864 6193 17867
rect 6052 17836 6193 17864
rect 6052 17824 6058 17836
rect 6181 17833 6193 17836
rect 6227 17833 6239 17867
rect 6546 17864 6552 17876
rect 6507 17836 6552 17864
rect 6181 17827 6239 17833
rect 6546 17824 6552 17836
rect 6604 17824 6610 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 6788 17836 7849 17864
rect 6788 17824 6794 17836
rect 5810 17756 5816 17808
rect 5868 17796 5874 17808
rect 6454 17796 6460 17808
rect 5868 17768 6040 17796
rect 6415 17768 6460 17796
rect 5868 17756 5874 17768
rect 4890 17688 4896 17740
rect 4948 17728 4954 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4948 17700 4997 17728
rect 4948 17688 4954 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 5905 17731 5963 17737
rect 5905 17728 5917 17731
rect 5224 17700 5917 17728
rect 5224 17688 5230 17700
rect 5905 17697 5917 17700
rect 5951 17697 5963 17731
rect 6012 17728 6040 17768
rect 6454 17756 6460 17768
rect 6512 17756 6518 17808
rect 6748 17768 7236 17796
rect 6748 17737 6776 17768
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6012 17700 6745 17728
rect 5905 17691 5963 17697
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 7098 17728 7104 17740
rect 7059 17700 7104 17728
rect 6733 17691 6791 17697
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 7208 17737 7236 17768
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 1946 17660 1952 17672
rect 1627 17632 1952 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 3154 17663 3212 17669
rect 3154 17660 3166 17663
rect 2832 17632 3166 17660
rect 2832 17620 2838 17632
rect 3154 17629 3166 17632
rect 3200 17629 3212 17663
rect 3154 17623 3212 17629
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3510 17660 3516 17672
rect 3467 17632 3516 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3510 17620 3516 17632
rect 3568 17660 3574 17672
rect 3605 17663 3663 17669
rect 3605 17660 3617 17663
rect 3568 17632 3617 17660
rect 3568 17620 3574 17632
rect 3605 17629 3617 17632
rect 3651 17660 3663 17663
rect 3881 17663 3939 17669
rect 3881 17660 3893 17663
rect 3651 17632 3893 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 3881 17629 3893 17632
rect 3927 17660 3939 17663
rect 4522 17660 4528 17672
rect 3927 17632 4528 17660
rect 3927 17629 3939 17632
rect 3881 17623 3939 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 4614 17620 4620 17672
rect 4672 17660 4678 17672
rect 4672 17632 6500 17660
rect 4672 17620 4678 17632
rect 4893 17595 4951 17601
rect 4893 17561 4905 17595
rect 4939 17592 4951 17595
rect 5994 17592 6000 17604
rect 4939 17564 6000 17592
rect 4939 17561 4951 17564
rect 4893 17555 4951 17561
rect 5994 17552 6000 17564
rect 6052 17552 6058 17604
rect 2038 17524 2044 17536
rect 1999 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 5258 17524 5264 17536
rect 4304 17496 5264 17524
rect 4304 17484 4310 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5721 17527 5779 17533
rect 5721 17524 5733 17527
rect 5592 17496 5733 17524
rect 5592 17484 5598 17496
rect 5721 17493 5733 17496
rect 5767 17493 5779 17527
rect 5721 17487 5779 17493
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 6472 17524 6500 17632
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 7285 17663 7343 17669
rect 7285 17660 7297 17663
rect 6604 17632 7297 17660
rect 6604 17620 6610 17632
rect 7285 17629 7297 17632
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 7576 17592 7604 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 8757 17867 8815 17873
rect 8757 17833 8769 17867
rect 8803 17864 8815 17867
rect 9306 17864 9312 17876
rect 8803 17836 9312 17864
rect 8803 17833 8815 17836
rect 8757 17827 8815 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 12066 17864 12072 17876
rect 9456 17836 12072 17864
rect 9456 17824 9462 17836
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 12342 17864 12348 17876
rect 12299 17836 12348 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 20073 17867 20131 17873
rect 20073 17833 20085 17867
rect 20119 17864 20131 17867
rect 20438 17864 20444 17876
rect 20119 17836 20444 17864
rect 20119 17833 20131 17836
rect 20073 17827 20131 17833
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 21542 17864 21548 17876
rect 21503 17836 21548 17864
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17765 7711 17799
rect 7653 17759 7711 17765
rect 7668 17660 7696 17759
rect 8478 17756 8484 17808
rect 8536 17796 8542 17808
rect 8941 17799 8999 17805
rect 8941 17796 8953 17799
rect 8536 17768 8953 17796
rect 8536 17756 8542 17768
rect 8941 17765 8953 17768
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 9122 17756 9128 17808
rect 9180 17796 9186 17808
rect 9861 17799 9919 17805
rect 9861 17796 9873 17799
rect 9180 17768 9873 17796
rect 9180 17756 9186 17768
rect 9861 17765 9873 17768
rect 9907 17765 9919 17799
rect 9861 17759 9919 17765
rect 11333 17799 11391 17805
rect 11333 17765 11345 17799
rect 11379 17796 11391 17799
rect 13354 17796 13360 17808
rect 11379 17768 13360 17796
rect 11379 17765 11391 17768
rect 11333 17759 11391 17765
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 19886 17756 19892 17808
rect 19944 17796 19950 17808
rect 20165 17799 20223 17805
rect 20165 17796 20177 17799
rect 19944 17768 20177 17796
rect 19944 17756 19950 17768
rect 20165 17765 20177 17768
rect 20211 17765 20223 17799
rect 20165 17759 20223 17765
rect 8205 17731 8263 17737
rect 8205 17697 8217 17731
rect 8251 17728 8263 17731
rect 8294 17728 8300 17740
rect 8251 17700 8300 17728
rect 8251 17697 8263 17700
rect 8205 17691 8263 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 9490 17728 9496 17740
rect 9451 17700 9496 17728
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10226 17728 10232 17740
rect 10183 17700 10232 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10962 17728 10968 17740
rect 10827 17700 10968 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11756 17700 11989 17728
rect 11756 17688 11762 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 12802 17728 12808 17740
rect 12763 17700 12808 17728
rect 11977 17691 12035 17697
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15580 17700 16221 17728
rect 11793 17663 11851 17669
rect 7668 17632 11560 17660
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 7576 17564 9413 17592
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 10686 17592 10692 17604
rect 9447 17564 10692 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 10686 17552 10692 17564
rect 10744 17552 10750 17604
rect 10965 17595 11023 17601
rect 10965 17561 10977 17595
rect 11011 17592 11023 17595
rect 11532 17592 11560 17632
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 12710 17660 12716 17672
rect 11839 17632 12716 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 14458 17669 14464 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13136 17632 14197 17660
rect 13136 17620 13142 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14452 17660 14464 17669
rect 14419 17632 14464 17660
rect 14185 17623 14243 17629
rect 14452 17623 14464 17632
rect 14516 17660 14522 17672
rect 15470 17660 15476 17672
rect 14516 17632 15476 17660
rect 14458 17620 14464 17623
rect 14516 17620 14522 17632
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 12526 17592 12532 17604
rect 11011 17564 11468 17592
rect 11532 17564 12532 17592
rect 11011 17561 11023 17564
rect 10965 17555 11023 17561
rect 8018 17524 8024 17536
rect 5868 17496 5913 17524
rect 6472 17496 8024 17524
rect 5868 17484 5874 17496
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 8260 17496 8309 17524
rect 8260 17484 8266 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 8570 17524 8576 17536
rect 8435 17496 8576 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 8812 17496 9321 17524
rect 8812 17484 8818 17496
rect 9309 17493 9321 17496
rect 9355 17524 9367 17527
rect 10229 17527 10287 17533
rect 10229 17524 10241 17527
rect 9355 17496 10241 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 10229 17493 10241 17496
rect 10275 17493 10287 17527
rect 10229 17487 10287 17493
rect 10873 17527 10931 17533
rect 10873 17493 10885 17527
rect 10919 17524 10931 17527
rect 11054 17524 11060 17536
rect 10919 17496 11060 17524
rect 10919 17493 10931 17496
rect 10873 17487 10931 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11440 17533 11468 17564
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 12621 17595 12679 17601
rect 12621 17561 12633 17595
rect 12667 17592 12679 17595
rect 12986 17592 12992 17604
rect 12667 17564 12992 17592
rect 12667 17561 12679 17564
rect 12621 17555 12679 17561
rect 12986 17552 12992 17564
rect 13044 17592 13050 17604
rect 14734 17592 14740 17604
rect 13044 17564 14740 17592
rect 13044 17552 13050 17564
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 11425 17527 11483 17533
rect 11425 17493 11437 17527
rect 11471 17493 11483 17527
rect 11882 17524 11888 17536
rect 11843 17496 11888 17524
rect 11425 17487 11483 17493
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 12768 17496 13093 17524
rect 12768 17484 12774 17496
rect 13081 17493 13093 17496
rect 13127 17493 13139 17527
rect 13081 17487 13139 17493
rect 15378 17484 15384 17536
rect 15436 17524 15442 17536
rect 15580 17533 15608 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16209 17691 16267 17697
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15712 17632 16129 17660
rect 15712 17620 15718 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 20180 17660 20208 17759
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 20180 17632 20361 17660
rect 16117 17623 16175 17629
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17660 20959 17663
rect 21560 17660 21588 17824
rect 20947 17632 21588 17660
rect 20947 17629 20959 17632
rect 20901 17623 20959 17629
rect 16025 17595 16083 17601
rect 16025 17561 16037 17595
rect 16071 17592 16083 17595
rect 16206 17592 16212 17604
rect 16071 17564 16212 17592
rect 16071 17561 16083 17564
rect 16025 17555 16083 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 20625 17595 20683 17601
rect 20625 17592 20637 17595
rect 20364 17564 20637 17592
rect 20364 17536 20392 17564
rect 20625 17561 20637 17564
rect 20671 17561 20683 17595
rect 20625 17555 20683 17561
rect 21177 17595 21235 17601
rect 21177 17561 21189 17595
rect 21223 17592 21235 17595
rect 21542 17592 21548 17604
rect 21223 17564 21548 17592
rect 21223 17561 21235 17564
rect 21177 17555 21235 17561
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 15565 17527 15623 17533
rect 15565 17524 15577 17527
rect 15436 17496 15577 17524
rect 15436 17484 15442 17496
rect 15565 17493 15577 17496
rect 15611 17493 15623 17527
rect 15565 17487 15623 17493
rect 15654 17484 15660 17536
rect 15712 17524 15718 17536
rect 15712 17496 15757 17524
rect 15712 17484 15718 17496
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 16448 17496 16589 17524
rect 16448 17484 16454 17496
rect 16577 17493 16589 17496
rect 16623 17524 16635 17527
rect 19610 17524 19616 17536
rect 16623 17496 19616 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 20346 17484 20352 17536
rect 20404 17484 20410 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 3421 17323 3479 17329
rect 3421 17320 3433 17323
rect 2924 17292 3433 17320
rect 2924 17280 2930 17292
rect 3421 17289 3433 17292
rect 3467 17320 3479 17323
rect 5445 17323 5503 17329
rect 3467 17292 3801 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 2038 17212 2044 17264
rect 2096 17252 2102 17264
rect 2286 17255 2344 17261
rect 2286 17252 2298 17255
rect 2096 17224 2298 17252
rect 2096 17212 2102 17224
rect 2286 17221 2298 17224
rect 2332 17221 2344 17255
rect 3602 17252 3608 17264
rect 2286 17215 2344 17221
rect 3436 17224 3608 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 1949 17187 2007 17193
rect 1949 17184 1961 17187
rect 1627 17156 1961 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 1949 17153 1961 17156
rect 1995 17184 2007 17187
rect 3436 17184 3464 17224
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 3773 17261 3801 17292
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5718 17320 5724 17332
rect 5491 17292 5724 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 5828 17292 7021 17320
rect 3758 17255 3816 17261
rect 3758 17221 3770 17255
rect 3804 17221 3816 17255
rect 3758 17215 3816 17221
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 5828 17252 5856 17292
rect 7009 17289 7021 17292
rect 7055 17320 7067 17323
rect 7282 17320 7288 17332
rect 7055 17292 7288 17320
rect 7055 17289 7067 17292
rect 7009 17283 7067 17289
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 8202 17320 8208 17332
rect 8163 17292 8208 17320
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8720 17292 9045 17320
rect 8720 17280 8726 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9180 17292 9413 17320
rect 9180 17280 9186 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 10226 17320 10232 17332
rect 9539 17292 10232 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11606 17320 11612 17332
rect 11287 17292 11612 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 11790 17320 11796 17332
rect 11703 17292 11796 17320
rect 11790 17280 11796 17292
rect 11848 17320 11854 17332
rect 12437 17323 12495 17329
rect 11848 17292 12112 17320
rect 11848 17280 11854 17292
rect 3936 17224 5856 17252
rect 3936 17212 3942 17224
rect 5902 17212 5908 17264
rect 5960 17212 5966 17264
rect 7098 17212 7104 17264
rect 7156 17252 7162 17264
rect 7156 17224 12020 17252
rect 7156 17212 7162 17224
rect 1995 17156 3464 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 5224 17156 5273 17184
rect 5224 17144 5230 17156
rect 5261 17153 5273 17156
rect 5307 17184 5319 17187
rect 5813 17187 5871 17193
rect 5813 17184 5825 17187
rect 5307 17156 5825 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 5813 17153 5825 17156
rect 5859 17153 5871 17187
rect 5920 17184 5948 17212
rect 6914 17184 6920 17196
rect 5920 17156 6040 17184
rect 6875 17156 6920 17184
rect 5813 17147 5871 17153
rect 2041 17119 2099 17125
rect 2041 17085 2053 17119
rect 2087 17085 2099 17119
rect 3510 17116 3516 17128
rect 3471 17088 3516 17116
rect 2041 17079 2099 17085
rect 2056 16980 2084 17079
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 5902 17116 5908 17128
rect 5863 17088 5908 17116
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 6012 17125 6040 17156
rect 6914 17144 6920 17156
rect 6972 17184 6978 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 6972 17156 7389 17184
rect 6972 17144 6978 17156
rect 7377 17153 7389 17156
rect 7423 17184 7435 17187
rect 7650 17184 7656 17196
rect 7423 17156 7656 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 7760 17156 8585 17184
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17116 6055 17119
rect 6086 17116 6092 17128
rect 6043 17088 6092 17116
rect 6043 17085 6055 17088
rect 5997 17079 6055 17085
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 6457 17119 6515 17125
rect 6457 17085 6469 17119
rect 6503 17116 6515 17119
rect 7006 17116 7012 17128
rect 6503 17088 7012 17116
rect 6503 17085 6515 17088
rect 6457 17079 6515 17085
rect 3528 16980 3556 17076
rect 4893 17051 4951 17057
rect 4893 17017 4905 17051
rect 4939 17048 4951 17051
rect 4982 17048 4988 17060
rect 4939 17020 4988 17048
rect 4939 17017 4951 17020
rect 4893 17011 4951 17017
rect 4982 17008 4988 17020
rect 5040 17048 5046 17060
rect 5350 17048 5356 17060
rect 5040 17020 5356 17048
rect 5040 17008 5046 17020
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 6472 17048 6500 17079
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17085 7159 17119
rect 7101 17079 7159 17085
rect 5460 17020 6500 17048
rect 7116 17048 7144 17079
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7760 17125 7788 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 10060 17184 10088 17224
rect 10117 17187 10175 17193
rect 10117 17184 10129 17187
rect 10060 17156 10129 17184
rect 8573 17147 8631 17153
rect 10117 17153 10129 17156
rect 10163 17153 10175 17187
rect 10117 17147 10175 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 11885 17187 11943 17193
rect 11885 17184 11897 17187
rect 10744 17156 11897 17184
rect 10744 17144 10750 17156
rect 11885 17153 11897 17156
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7248 17088 7757 17116
rect 7248 17076 7254 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17116 8171 17119
rect 8386 17116 8392 17128
rect 8159 17088 8392 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17085 8723 17119
rect 8665 17079 8723 17085
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17116 8815 17119
rect 9490 17116 9496 17128
rect 8803 17088 9496 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 7466 17048 7472 17060
rect 7116 17020 7472 17048
rect 2056 16952 3556 16980
rect 4614 16940 4620 16992
rect 4672 16980 4678 16992
rect 5077 16983 5135 16989
rect 5077 16980 5089 16983
rect 4672 16952 5089 16980
rect 4672 16940 4678 16952
rect 5077 16949 5089 16952
rect 5123 16980 5135 16983
rect 5460 16980 5488 17020
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 8680 17048 8708 17079
rect 7668 17020 8708 17048
rect 7668 16992 7696 17020
rect 6546 16980 6552 16992
rect 5123 16952 5488 16980
rect 6507 16952 6552 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 7650 16980 7656 16992
rect 7611 16952 7656 16980
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8772 16980 8800 17079
rect 9490 17076 9496 17088
rect 9548 17116 9554 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9548 17088 9597 17116
rect 9548 17076 9554 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9732 17088 9873 17116
rect 9732 17076 9738 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17116 11759 17119
rect 11790 17116 11796 17128
rect 11747 17088 11796 17116
rect 11747 17085 11759 17088
rect 11701 17079 11759 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11900 17048 11928 17147
rect 11992 17116 12020 17224
rect 12084 17184 12112 17292
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12986 17320 12992 17332
rect 12483 17292 12992 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13814 17320 13820 17332
rect 13775 17292 13820 17320
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 14231 17292 14657 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 15013 17323 15071 17329
rect 15013 17289 15025 17323
rect 15059 17320 15071 17323
rect 15654 17320 15660 17332
rect 15059 17292 15660 17320
rect 15059 17289 15071 17292
rect 15013 17283 15071 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 16390 17320 16396 17332
rect 15804 17292 15849 17320
rect 16351 17292 16396 17320
rect 15804 17280 15810 17292
rect 16390 17280 16396 17292
rect 16448 17280 16454 17332
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21082 17320 21088 17332
rect 21039 17292 21088 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 21358 17320 21364 17332
rect 21319 17292 21364 17320
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 12897 17255 12955 17261
rect 12897 17252 12909 17255
rect 12216 17224 12909 17252
rect 12216 17212 12222 17224
rect 12897 17221 12909 17224
rect 12943 17221 12955 17255
rect 12897 17215 12955 17221
rect 14277 17255 14335 17261
rect 14277 17221 14289 17255
rect 14323 17252 14335 17255
rect 14323 17224 15700 17252
rect 14323 17221 14335 17224
rect 14277 17215 14335 17221
rect 15672 17196 15700 17224
rect 12713 17187 12771 17193
rect 12713 17184 12725 17187
rect 12084 17156 12725 17184
rect 12713 17153 12725 17156
rect 12759 17153 12771 17187
rect 12713 17147 12771 17153
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15286 17184 15292 17196
rect 15151 17156 15292 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 15838 17184 15844 17196
rect 15799 17156 15844 17184
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 19978 17184 19984 17196
rect 19939 17156 19984 17184
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 12342 17116 12348 17128
rect 11992 17088 12348 17116
rect 12342 17076 12348 17088
rect 12400 17116 12406 17128
rect 12802 17116 12808 17128
rect 12400 17088 12808 17116
rect 12400 17076 12406 17088
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 13228 17088 14381 17116
rect 13228 17076 13234 17088
rect 14369 17085 14381 17088
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 15197 17119 15255 17125
rect 15197 17085 15209 17119
rect 15243 17085 15255 17119
rect 15197 17079 15255 17085
rect 12066 17048 12072 17060
rect 11900 17020 12072 17048
rect 12066 17008 12072 17020
rect 12124 17008 12130 17060
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12526 17048 12532 17060
rect 12299 17020 12532 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17048 12679 17051
rect 13078 17048 13084 17060
rect 12667 17020 13084 17048
rect 12667 17017 12679 17020
rect 12621 17011 12679 17017
rect 13078 17008 13084 17020
rect 13136 17048 13142 17060
rect 13262 17048 13268 17060
rect 13136 17020 13268 17048
rect 13136 17008 13142 17020
rect 13262 17008 13268 17020
rect 13320 17008 13326 17060
rect 14274 17008 14280 17060
rect 14332 17048 14338 17060
rect 15212 17048 15240 17079
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 15565 17119 15623 17125
rect 15565 17116 15577 17119
rect 15436 17088 15577 17116
rect 15436 17076 15442 17088
rect 15565 17085 15577 17088
rect 15611 17085 15623 17119
rect 21192 17116 21220 17147
rect 15565 17079 15623 17085
rect 20456 17088 21220 17116
rect 16114 17048 16120 17060
rect 14332 17020 16120 17048
rect 14332 17008 14338 17020
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 8352 16952 8800 16980
rect 8352 16940 8358 16952
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 12986 16980 12992 16992
rect 12216 16952 12992 16980
rect 12216 16940 12222 16952
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16209 16983 16267 16989
rect 16209 16980 16221 16983
rect 16080 16952 16221 16980
rect 16080 16940 16086 16952
rect 16209 16949 16221 16952
rect 16255 16949 16267 16983
rect 16758 16980 16764 16992
rect 16719 16952 16764 16980
rect 16209 16943 16267 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20456 16989 20484 17088
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19944 16952 20453 16980
rect 19944 16940 19950 16952
rect 20441 16949 20453 16952
rect 20487 16949 20499 16983
rect 20441 16943 20499 16949
rect 20717 16983 20775 16989
rect 20717 16949 20729 16983
rect 20763 16980 20775 16983
rect 20806 16980 20812 16992
rect 20763 16952 20812 16980
rect 20763 16949 20775 16952
rect 20717 16943 20775 16949
rect 20806 16940 20812 16952
rect 20864 16980 20870 16992
rect 22462 16980 22468 16992
rect 20864 16952 22468 16980
rect 20864 16940 20870 16952
rect 22462 16940 22468 16952
rect 22520 16940 22526 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2777 16779 2835 16785
rect 2777 16776 2789 16779
rect 1964 16748 2789 16776
rect 1964 16572 1992 16748
rect 2777 16745 2789 16748
rect 2823 16776 2835 16779
rect 4890 16776 4896 16788
rect 2823 16748 4896 16776
rect 2823 16745 2835 16748
rect 2777 16739 2835 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 5960 16748 6561 16776
rect 5960 16736 5966 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 6549 16739 6607 16745
rect 7098 16736 7104 16788
rect 7156 16776 7162 16788
rect 7926 16776 7932 16788
rect 7156 16748 7932 16776
rect 7156 16736 7162 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8076 16748 8432 16776
rect 8076 16736 8082 16748
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2096 16680 3556 16708
rect 2096 16668 2102 16680
rect 3528 16649 3556 16680
rect 5718 16668 5724 16720
rect 5776 16708 5782 16720
rect 6086 16708 6092 16720
rect 5776 16680 6092 16708
rect 5776 16668 5782 16680
rect 6086 16668 6092 16680
rect 6144 16668 6150 16720
rect 7377 16711 7435 16717
rect 7377 16708 7389 16711
rect 7024 16680 7389 16708
rect 7024 16652 7052 16680
rect 7377 16677 7389 16680
rect 7423 16677 7435 16711
rect 7377 16671 7435 16677
rect 8036 16680 8340 16708
rect 8036 16652 8064 16680
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16640 3571 16643
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3559 16612 4353 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4672 16612 4721 16640
rect 4672 16600 4678 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 7006 16640 7012 16652
rect 4709 16603 4767 16609
rect 5736 16612 6868 16640
rect 6967 16612 7012 16640
rect 2041 16575 2099 16581
rect 2041 16572 2053 16575
rect 1964 16544 2053 16572
rect 2041 16541 2053 16544
rect 2087 16541 2099 16575
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2041 16535 2099 16541
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 2590 16572 2596 16584
rect 2551 16544 2596 16572
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 3326 16572 3332 16584
rect 3287 16544 3332 16572
rect 3326 16532 3332 16544
rect 3384 16532 3390 16584
rect 4982 16581 4988 16584
rect 4965 16575 4988 16581
rect 4965 16572 4977 16575
rect 4895 16544 4977 16572
rect 4965 16541 4977 16544
rect 5040 16572 5046 16584
rect 5736 16572 5764 16612
rect 5040 16544 5764 16572
rect 6840 16572 6868 16612
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7466 16640 7472 16652
rect 7239 16612 7472 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7208 16572 7236 16603
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8018 16640 8024 16652
rect 7975 16612 8024 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8312 16649 8340 16680
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16609 8355 16643
rect 8404 16640 8432 16748
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 8628 16748 8769 16776
rect 8628 16736 8634 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9398 16776 9404 16788
rect 9079 16748 9404 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 10873 16779 10931 16785
rect 10873 16776 10885 16779
rect 9876 16748 10885 16776
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 9876 16708 9904 16748
rect 10873 16745 10885 16748
rect 10919 16776 10931 16779
rect 10919 16748 11367 16776
rect 10919 16745 10931 16748
rect 10873 16739 10931 16745
rect 11238 16708 11244 16720
rect 8536 16680 9904 16708
rect 9968 16680 11244 16708
rect 8536 16668 8542 16680
rect 9968 16649 9996 16680
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 9953 16643 10011 16649
rect 8404 16612 9904 16640
rect 8297 16603 8355 16609
rect 6840 16544 7236 16572
rect 4965 16535 4988 16541
rect 4982 16532 4988 16535
rect 5040 16532 5046 16544
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7340 16544 7573 16572
rect 7340 16532 7346 16544
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 8386 16572 8392 16584
rect 8347 16544 8392 16572
rect 7561 16535 7619 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 9876 16572 9904 16612
rect 9953 16609 9965 16643
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 10042 16600 10048 16652
rect 10100 16640 10106 16652
rect 10781 16643 10839 16649
rect 10100 16612 10145 16640
rect 10100 16600 10106 16612
rect 10781 16609 10793 16643
rect 10827 16640 10839 16643
rect 11339 16640 11367 16748
rect 11698 16736 11704 16788
rect 11756 16776 11762 16788
rect 11882 16776 11888 16788
rect 11756 16748 11888 16776
rect 11756 16736 11762 16748
rect 11882 16736 11888 16748
rect 11940 16776 11946 16788
rect 14093 16779 14151 16785
rect 11940 16748 14044 16776
rect 11940 16736 11946 16748
rect 14016 16708 14044 16748
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14274 16776 14280 16788
rect 14139 16748 14280 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 15565 16779 15623 16785
rect 14568 16748 15516 16776
rect 14568 16708 14596 16748
rect 14016 16680 14596 16708
rect 15488 16708 15516 16748
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 15654 16776 15660 16788
rect 15611 16748 15660 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 15804 16748 17233 16776
rect 15804 16736 15810 16748
rect 17221 16745 17233 16748
rect 17267 16745 17279 16779
rect 19518 16776 19524 16788
rect 17221 16739 17279 16745
rect 17880 16748 19524 16776
rect 17880 16720 17908 16748
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 20993 16779 21051 16785
rect 20993 16745 21005 16779
rect 21039 16776 21051 16779
rect 21082 16776 21088 16788
rect 21039 16748 21088 16776
rect 21039 16745 21051 16748
rect 20993 16739 21051 16745
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 17405 16711 17463 16717
rect 17405 16708 17417 16711
rect 15488 16680 17417 16708
rect 17405 16677 17417 16680
rect 17451 16708 17463 16711
rect 17862 16708 17868 16720
rect 17451 16680 17868 16708
rect 17451 16677 17463 16680
rect 17405 16671 17463 16677
rect 17862 16668 17868 16680
rect 17920 16668 17926 16720
rect 11606 16640 11612 16652
rect 10827 16612 11100 16640
rect 11339 16612 11468 16640
rect 11567 16612 11612 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 11072 16584 11100 16612
rect 10134 16572 10140 16584
rect 9876 16544 10140 16572
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11440 16572 11468 16612
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 13262 16640 13268 16652
rect 13223 16612 13268 16640
rect 13262 16600 13268 16612
rect 13320 16640 13326 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13320 16612 13553 16640
rect 13320 16600 13326 16612
rect 13541 16609 13553 16612
rect 13587 16640 13599 16643
rect 14458 16640 14464 16652
rect 13587 16612 14464 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 16022 16640 16028 16652
rect 15983 16612 16028 16640
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16172 16612 16217 16640
rect 16316 16612 16957 16640
rect 16172 16600 16178 16612
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11112 16544 11376 16572
rect 11440 16544 11529 16572
rect 11112 16532 11118 16544
rect 3142 16464 3148 16516
rect 3200 16504 3206 16516
rect 3200 16476 3832 16504
rect 3200 16464 3206 16476
rect 2869 16439 2927 16445
rect 2869 16405 2881 16439
rect 2915 16436 2927 16439
rect 3050 16436 3056 16448
rect 2915 16408 3056 16436
rect 2915 16405 2927 16408
rect 2869 16399 2927 16405
rect 3050 16396 3056 16408
rect 3108 16396 3114 16448
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3694 16436 3700 16448
rect 3283 16408 3700 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 3804 16445 3832 16476
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 4120 16476 4261 16504
rect 4120 16464 4126 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 4249 16467 4307 16473
rect 5810 16464 5816 16516
rect 5868 16504 5874 16516
rect 6181 16507 6239 16513
rect 6181 16504 6193 16507
rect 5868 16476 6193 16504
rect 5868 16464 5874 16476
rect 6181 16473 6193 16476
rect 6227 16473 6239 16507
rect 6181 16467 6239 16473
rect 6454 16464 6460 16516
rect 6512 16504 6518 16516
rect 7006 16504 7012 16516
rect 6512 16476 7012 16504
rect 6512 16464 6518 16476
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11348 16504 11376 16544
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 13009 16575 13067 16581
rect 13009 16541 13021 16575
rect 13055 16572 13067 16575
rect 13170 16572 13176 16584
rect 13055 16544 13176 16572
rect 13055 16541 13067 16544
rect 13009 16535 13067 16541
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 14476 16572 14504 16600
rect 15473 16575 15531 16581
rect 15473 16572 15485 16575
rect 14476 16544 15485 16572
rect 15473 16541 15485 16544
rect 15519 16541 15531 16575
rect 16316 16572 16344 16612
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 19978 16640 19984 16652
rect 19567 16612 19984 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 15473 16535 15531 16541
rect 15856 16544 16344 16572
rect 13449 16507 13507 16513
rect 11020 16476 11100 16504
rect 11020 16464 11026 16476
rect 3789 16439 3847 16445
rect 3789 16405 3801 16439
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4157 16439 4215 16445
rect 4157 16436 4169 16439
rect 3936 16408 4169 16436
rect 3936 16396 3942 16408
rect 4157 16405 4169 16408
rect 4203 16405 4215 16439
rect 4157 16399 4215 16405
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 6917 16439 6975 16445
rect 6917 16436 6929 16439
rect 6880 16408 6929 16436
rect 6880 16396 6886 16408
rect 6917 16405 6929 16408
rect 6963 16405 6975 16439
rect 9490 16436 9496 16448
rect 9451 16408 9496 16436
rect 6917 16399 6975 16405
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 9858 16436 9864 16448
rect 9819 16408 9864 16436
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 11072 16445 11100 16476
rect 11348 16476 12434 16504
rect 11057 16439 11115 16445
rect 11057 16405 11069 16439
rect 11103 16405 11115 16439
rect 11348 16436 11376 16476
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 11348 16408 11437 16436
rect 11057 16399 11115 16405
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11425 16399 11483 16405
rect 11790 16396 11796 16448
rect 11848 16436 11854 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11848 16408 11897 16436
rect 11848 16396 11854 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 12406 16436 12434 16476
rect 13449 16473 13461 16507
rect 13495 16504 13507 16507
rect 13630 16504 13636 16516
rect 13495 16476 13636 16504
rect 13495 16473 13507 16476
rect 13449 16467 13507 16473
rect 13630 16464 13636 16476
rect 13688 16464 13694 16516
rect 15194 16464 15200 16516
rect 15252 16513 15258 16516
rect 15252 16504 15264 16513
rect 15378 16504 15384 16516
rect 15252 16476 15384 16504
rect 15252 16467 15264 16476
rect 15252 16464 15258 16467
rect 15378 16464 15384 16476
rect 15436 16504 15442 16516
rect 15856 16504 15884 16544
rect 17402 16532 17408 16584
rect 17460 16572 17466 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 17460 16544 19257 16572
rect 17460 16532 17466 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16572 20867 16575
rect 20855 16544 20889 16572
rect 20855 16541 20867 16544
rect 20809 16535 20867 16541
rect 15436 16476 15884 16504
rect 15933 16507 15991 16513
rect 15436 16464 15442 16476
rect 15933 16473 15945 16507
rect 15979 16504 15991 16507
rect 16758 16504 16764 16516
rect 15979 16476 16436 16504
rect 16671 16476 16764 16504
rect 15979 16473 15991 16476
rect 15933 16467 15991 16473
rect 16298 16436 16304 16448
rect 12406 16408 16304 16436
rect 11885 16399 11943 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16408 16445 16436 16476
rect 16758 16464 16764 16476
rect 16816 16504 16822 16516
rect 17586 16504 17592 16516
rect 16816 16476 17592 16504
rect 16816 16464 16822 16476
rect 17586 16464 17592 16476
rect 17644 16504 17650 16516
rect 20162 16504 20168 16516
rect 17644 16476 20168 16504
rect 17644 16464 17650 16476
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 20717 16507 20775 16513
rect 20717 16473 20729 16507
rect 20763 16504 20775 16507
rect 20824 16504 20852 16535
rect 22554 16504 22560 16516
rect 20763 16476 22560 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 16393 16439 16451 16445
rect 16393 16405 16405 16439
rect 16439 16405 16451 16439
rect 16393 16399 16451 16405
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 17034 16436 17040 16448
rect 16899 16408 17040 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 21174 16436 21180 16448
rect 21135 16408 21180 16436
rect 21174 16396 21180 16408
rect 21232 16396 21238 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3878 16232 3884 16244
rect 3743 16204 3884 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3878 16192 3884 16204
rect 3936 16192 3942 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 4203 16204 4629 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4617 16201 4629 16204
rect 4663 16201 4675 16235
rect 4617 16195 4675 16201
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 5534 16232 5540 16244
rect 5491 16204 5540 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 5810 16232 5816 16244
rect 5771 16204 5816 16232
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7282 16232 7288 16244
rect 7239 16204 7288 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7282 16192 7288 16204
rect 7340 16232 7346 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7340 16204 7849 16232
rect 7340 16192 7346 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 7837 16195 7895 16201
rect 8036 16204 8401 16232
rect 3068 16136 4384 16164
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2179 16068 2544 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2222 15892 2228 15904
rect 2183 15864 2228 15892
rect 2222 15852 2228 15864
rect 2280 15852 2286 15904
rect 2516 15901 2544 16068
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3068 16037 3096 16136
rect 3896 16108 3924 16136
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 3418 16096 3424 16108
rect 3375 16068 3424 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3878 16056 3884 16108
rect 3936 16056 3942 16108
rect 3053 16031 3111 16037
rect 3053 16028 3065 16031
rect 2924 16000 3065 16028
rect 2924 15988 2930 16000
rect 3053 15997 3065 16000
rect 3099 15997 3111 16031
rect 3053 15991 3111 15997
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 4246 16028 4252 16040
rect 4207 16000 4252 16028
rect 3237 15991 3295 15997
rect 2501 15895 2559 15901
rect 2501 15861 2513 15895
rect 2547 15892 2559 15895
rect 2682 15892 2688 15904
rect 2547 15864 2688 15892
rect 2547 15861 2559 15864
rect 2501 15855 2559 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 2958 15892 2964 15904
rect 2915 15864 2964 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 2958 15852 2964 15864
rect 3016 15892 3022 15904
rect 3252 15892 3280 15991
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 4356 16037 4384 16136
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 4764 16136 6561 16164
rect 4764 16124 4770 16136
rect 4982 16096 4988 16108
rect 4943 16068 4988 16096
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5184 16040 5212 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 6549 16127 6607 16133
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 8036 16173 8064 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 8389 16195 8447 16201
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 9490 16232 9496 16244
rect 8895 16204 9496 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 8021 16167 8079 16173
rect 8021 16164 8033 16167
rect 6972 16136 8033 16164
rect 6972 16124 6978 16136
rect 8021 16133 8033 16136
rect 8067 16133 8079 16167
rect 8404 16164 8432 16195
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 9582 16192 9588 16244
rect 9640 16232 9646 16244
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 9640 16204 10885 16232
rect 9640 16192 9646 16204
rect 10873 16201 10885 16204
rect 10919 16232 10931 16235
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10919 16204 11069 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 11057 16195 11115 16201
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 12584 16204 12909 16232
rect 12584 16192 12590 16204
rect 12897 16201 12909 16204
rect 12943 16201 12955 16235
rect 12897 16195 12955 16201
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13170 16232 13176 16244
rect 13127 16204 13176 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 15657 16235 15715 16241
rect 15657 16201 15669 16235
rect 15703 16232 15715 16235
rect 15746 16232 15752 16244
rect 15703 16204 15752 16232
rect 15703 16201 15715 16204
rect 15657 16195 15715 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 15896 16204 16129 16232
rect 15896 16192 15902 16204
rect 16117 16201 16129 16204
rect 16163 16201 16175 16235
rect 16117 16195 16175 16201
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 17037 16235 17095 16241
rect 16264 16204 16309 16232
rect 16264 16192 16270 16204
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17083 16204 17509 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17862 16192 17868 16244
rect 17920 16232 17926 16244
rect 17957 16235 18015 16241
rect 17957 16232 17969 16235
rect 17920 16204 17969 16232
rect 17920 16192 17926 16204
rect 17957 16201 17969 16204
rect 18003 16201 18015 16235
rect 20622 16232 20628 16244
rect 20583 16204 20628 16232
rect 17957 16195 18015 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20993 16235 21051 16241
rect 20993 16201 21005 16235
rect 21039 16232 21051 16235
rect 21082 16232 21088 16244
rect 21039 16204 21088 16232
rect 21039 16201 21051 16204
rect 20993 16195 21051 16201
rect 21082 16192 21088 16204
rect 21140 16192 21146 16244
rect 21358 16232 21364 16244
rect 21319 16204 21364 16232
rect 21358 16192 21364 16204
rect 21416 16192 21422 16244
rect 8404 16136 8892 16164
rect 8021 16127 8079 16133
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5776 16068 6040 16096
rect 5776 16056 5782 16068
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 15997 4399 16031
rect 4341 15991 4399 15997
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4948 16000 5089 16028
rect 4948 15988 4954 16000
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 5166 15988 5172 16040
rect 5224 16028 5230 16040
rect 6012 16037 6040 16068
rect 5905 16031 5963 16037
rect 5224 16000 5269 16028
rect 5224 15988 5230 16000
rect 5905 15997 5917 16031
rect 5951 15997 5963 16031
rect 5905 15991 5963 15997
rect 5997 16031 6055 16037
rect 5997 15997 6009 16031
rect 6043 15997 6055 16031
rect 6822 16028 6828 16040
rect 5997 15991 6055 15997
rect 6380 16000 6828 16028
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 3752 15932 3801 15960
rect 3752 15920 3758 15932
rect 3789 15929 3801 15932
rect 3835 15929 3847 15963
rect 3789 15923 3847 15929
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 5920 15960 5948 15991
rect 4856 15932 5948 15960
rect 4856 15920 4862 15932
rect 6380 15904 6408 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 15997 7343 16031
rect 7466 16028 7472 16040
rect 7427 16000 7472 16028
rect 7285 15991 7343 15997
rect 7300 15960 7328 15991
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8864 16028 8892 16136
rect 9214 16124 9220 16176
rect 9272 16164 9278 16176
rect 9668 16167 9726 16173
rect 9668 16164 9680 16167
rect 9272 16136 9680 16164
rect 9272 16124 9278 16136
rect 9668 16133 9680 16136
rect 9714 16164 9726 16167
rect 10042 16164 10048 16176
rect 9714 16136 10048 16164
rect 9714 16133 9726 16136
rect 9668 16127 9726 16133
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 12437 16167 12495 16173
rect 12437 16164 12449 16167
rect 10744 16136 12449 16164
rect 10744 16124 10750 16136
rect 12437 16133 12449 16136
rect 12483 16164 12495 16167
rect 13446 16164 13452 16176
rect 12483 16136 13452 16164
rect 12483 16133 12495 16136
rect 12437 16127 12495 16133
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 14274 16173 14280 16176
rect 14216 16167 14280 16173
rect 14216 16133 14228 16167
rect 14262 16133 14280 16167
rect 14216 16127 14280 16133
rect 14274 16124 14280 16127
rect 14332 16124 14338 16176
rect 15194 16164 15200 16176
rect 14660 16136 15200 16164
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9122 16096 9128 16108
rect 8987 16068 9128 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9390 16099 9448 16105
rect 9390 16096 9402 16099
rect 9232 16068 9402 16096
rect 9232 16028 9260 16068
rect 9390 16065 9402 16068
rect 9436 16065 9448 16099
rect 11146 16096 11152 16108
rect 9390 16059 9448 16065
rect 9508 16068 11152 16096
rect 9508 16028 9536 16068
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13630 16096 13636 16108
rect 12575 16068 13636 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14458 16096 14464 16108
rect 14419 16068 14464 16096
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 12342 16028 12348 16040
rect 8864 16000 9260 16028
rect 9324 16000 9536 16028
rect 12303 16000 12348 16028
rect 8757 15991 8815 15997
rect 7300 15932 7696 15960
rect 7668 15904 7696 15932
rect 6362 15892 6368 15904
rect 3016 15864 3280 15892
rect 6323 15864 6368 15892
rect 3016 15852 3022 15864
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7650 15892 7656 15904
rect 7611 15864 7656 15892
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 8772 15892 8800 15991
rect 9324 15969 9352 16000
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 14660 16037 14688 16136
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 16298 16124 16304 16176
rect 16356 16164 16362 16176
rect 18230 16164 18236 16176
rect 16356 16136 18236 16164
rect 16356 16124 16362 16136
rect 18230 16124 18236 16136
rect 18288 16164 18294 16176
rect 18325 16167 18383 16173
rect 18325 16164 18337 16167
rect 18288 16136 18337 16164
rect 18288 16124 18294 16136
rect 18325 16133 18337 16136
rect 18371 16133 18383 16167
rect 18325 16127 18383 16133
rect 18506 16124 18512 16176
rect 18564 16164 18570 16176
rect 20349 16167 20407 16173
rect 20349 16164 20361 16167
rect 18564 16136 20361 16164
rect 18564 16124 18570 16136
rect 20349 16133 20361 16136
rect 20395 16164 20407 16167
rect 20395 16136 20852 16164
rect 20395 16133 20407 16136
rect 20349 16127 20407 16133
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 16114 16096 16120 16108
rect 15795 16068 16120 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 17126 16056 17132 16108
rect 17184 16096 17190 16108
rect 17865 16099 17923 16105
rect 17865 16096 17877 16099
rect 17184 16068 17877 16096
rect 17184 16056 17190 16068
rect 17865 16065 17877 16068
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20824 16105 20852 16136
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 20036 16068 20453 16096
rect 20036 16056 20042 16068
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21174 16096 21180 16108
rect 20956 16068 21180 16096
rect 20956 16056 20962 16068
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 15997 14703 16031
rect 14826 16028 14832 16040
rect 14787 16000 14832 16028
rect 14645 15991 14703 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15470 16028 15476 16040
rect 15431 16000 15476 16028
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 16724 16000 16773 16028
rect 16724 15988 16730 16000
rect 16761 15997 16773 16000
rect 16807 15997 16819 16031
rect 16761 15991 16819 15997
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17770 16028 17776 16040
rect 16991 16000 17776 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18141 16031 18199 16037
rect 18141 15997 18153 16031
rect 18187 16028 18199 16031
rect 18414 16028 18420 16040
rect 18187 16000 18420 16028
rect 18187 15997 18199 16000
rect 18141 15991 18199 15997
rect 9309 15963 9367 15969
rect 9309 15929 9321 15963
rect 9355 15929 9367 15963
rect 9309 15923 9367 15929
rect 16390 15920 16396 15972
rect 16448 15960 16454 15972
rect 18156 15960 18184 15991
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 20622 16028 20628 16040
rect 18840 16000 20628 16028
rect 18840 15988 18846 16000
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 16448 15932 18184 15960
rect 16448 15920 16454 15932
rect 10778 15892 10784 15904
rect 8772 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 17862 15892 17868 15904
rect 17451 15864 17868 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 1949 15691 2007 15697
rect 1949 15688 1961 15691
rect 1912 15660 1961 15688
rect 1912 15648 1918 15660
rect 1949 15657 1961 15660
rect 1995 15657 2007 15691
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 1949 15651 2007 15657
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 4154 15688 4160 15700
rect 2832 15660 2877 15688
rect 4067 15660 4160 15688
rect 2832 15648 2838 15660
rect 4154 15648 4160 15660
rect 4212 15688 4218 15700
rect 4614 15688 4620 15700
rect 4212 15660 4620 15688
rect 4212 15648 4218 15660
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5994 15688 6000 15700
rect 5955 15660 6000 15688
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 7466 15688 7472 15700
rect 6380 15660 7472 15688
rect 6380 15620 6408 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 11885 15691 11943 15697
rect 7708 15660 11468 15688
rect 7708 15648 7714 15660
rect 6822 15620 6828 15632
rect 2976 15592 6408 15620
rect 6472 15592 6828 15620
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 2222 15484 2228 15496
rect 2179 15456 2228 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2516 15416 2544 15447
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 2648 15456 2693 15484
rect 2648 15444 2654 15456
rect 2976 15425 3004 15592
rect 3418 15552 3424 15564
rect 3379 15524 3424 15552
rect 3418 15512 3424 15524
rect 3476 15512 3482 15564
rect 6472 15561 6500 15592
rect 6822 15580 6828 15592
rect 6880 15580 6886 15632
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 8941 15623 8999 15629
rect 8941 15620 8953 15623
rect 8444 15592 8953 15620
rect 8444 15580 8450 15592
rect 8941 15589 8953 15592
rect 8987 15620 8999 15623
rect 9214 15620 9220 15632
rect 8987 15592 9220 15620
rect 8987 15589 8999 15592
rect 8941 15583 8999 15589
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 11440 15620 11468 15660
rect 11885 15657 11897 15691
rect 11931 15688 11943 15691
rect 12434 15688 12440 15700
rect 11931 15660 12440 15688
rect 11931 15657 11943 15660
rect 11885 15651 11943 15657
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 13446 15688 13452 15700
rect 13407 15660 13452 15688
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 14458 15648 14464 15700
rect 14516 15688 14522 15700
rect 14553 15691 14611 15697
rect 14553 15688 14565 15691
rect 14516 15660 14565 15688
rect 14516 15648 14522 15660
rect 14553 15657 14565 15660
rect 14599 15657 14611 15691
rect 14553 15651 14611 15657
rect 15841 15691 15899 15697
rect 15841 15657 15853 15691
rect 15887 15688 15899 15691
rect 17034 15688 17040 15700
rect 15887 15660 17040 15688
rect 15887 15657 15899 15660
rect 15841 15651 15899 15657
rect 12710 15620 12716 15632
rect 11440 15592 12716 15620
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 13357 15623 13415 15629
rect 13357 15589 13369 15623
rect 13403 15620 13415 15623
rect 13906 15620 13912 15632
rect 13403 15592 13912 15620
rect 13403 15589 13415 15592
rect 13357 15583 13415 15589
rect 13906 15580 13912 15592
rect 13964 15580 13970 15632
rect 14568 15620 14596 15651
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 17828 15660 17877 15688
rect 17828 15648 17834 15660
rect 17865 15657 17877 15660
rect 17911 15657 17923 15691
rect 21358 15688 21364 15700
rect 21319 15660 21364 15688
rect 17865 15651 17923 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 16298 15620 16304 15632
rect 14568 15592 16304 15620
rect 16298 15580 16304 15592
rect 16356 15620 16362 15632
rect 16356 15592 16436 15620
rect 16356 15580 16362 15592
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 6549 15555 6607 15561
rect 6549 15521 6561 15555
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 5166 15484 5172 15496
rect 4356 15456 5172 15484
rect 2961 15419 3019 15425
rect 2961 15416 2973 15419
rect 2516 15388 2973 15416
rect 2961 15385 2973 15388
rect 3007 15385 3019 15419
rect 2961 15379 3019 15385
rect 4356 15360 4384 15456
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 6564 15484 6592 15515
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7282 15552 7288 15564
rect 6972 15524 7288 15552
rect 6972 15512 6978 15524
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 12676 15524 12721 15552
rect 12676 15512 12682 15524
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 12952 15524 14381 15552
rect 12952 15512 12958 15524
rect 14369 15521 14381 15524
rect 14415 15552 14427 15555
rect 14826 15552 14832 15564
rect 14415 15524 14832 15552
rect 14415 15521 14427 15524
rect 14369 15515 14427 15521
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 15470 15552 15476 15564
rect 15335 15524 15476 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 16408 15561 16436 15592
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15521 16451 15555
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 16393 15515 16451 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 5776 15456 6592 15484
rect 5776 15444 5782 15456
rect 7374 15444 7380 15496
rect 7432 15484 7438 15496
rect 7541 15487 7599 15493
rect 7541 15484 7553 15487
rect 7432 15456 7553 15484
rect 7432 15444 7438 15456
rect 7541 15453 7553 15456
rect 7587 15453 7599 15487
rect 7541 15447 7599 15453
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10502 15484 10508 15496
rect 10367 15456 10508 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10778 15493 10784 15496
rect 10772 15484 10784 15493
rect 10739 15456 10784 15484
rect 10772 15447 10784 15456
rect 10778 15444 10784 15447
rect 10836 15444 10842 15496
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 14921 15487 14979 15493
rect 14921 15484 14933 15487
rect 12124 15456 14933 15484
rect 12124 15444 12130 15456
rect 14921 15453 14933 15456
rect 14967 15484 14979 15487
rect 15010 15484 15016 15496
rect 14967 15456 15016 15484
rect 14967 15453 14979 15456
rect 14921 15447 14979 15453
rect 4890 15376 4896 15428
rect 4948 15416 4954 15428
rect 5445 15419 5503 15425
rect 5445 15416 5457 15419
rect 4948 15388 5457 15416
rect 4948 15376 4954 15388
rect 5445 15385 5457 15388
rect 5491 15385 5503 15419
rect 5445 15379 5503 15385
rect 6365 15419 6423 15425
rect 6365 15385 6377 15419
rect 6411 15416 6423 15419
rect 6546 15416 6552 15428
rect 6411 15388 6552 15416
rect 6411 15385 6423 15388
rect 6365 15379 6423 15385
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 9214 15416 9220 15428
rect 8680 15388 9220 15416
rect 4338 15348 4344 15360
rect 4299 15320 4344 15348
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 5261 15351 5319 15357
rect 5261 15348 5273 15351
rect 4856 15320 5273 15348
rect 4856 15308 4862 15320
rect 5261 15317 5273 15320
rect 5307 15317 5319 15351
rect 5261 15311 5319 15317
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 8680 15357 8708 15388
rect 9214 15376 9220 15388
rect 9272 15416 9278 15428
rect 10054 15419 10112 15425
rect 10054 15416 10066 15419
rect 9272 15388 10066 15416
rect 9272 15376 9278 15388
rect 10054 15385 10066 15388
rect 10100 15416 10112 15419
rect 10594 15416 10600 15428
rect 10100 15388 10600 15416
rect 10100 15385 10112 15388
rect 10054 15379 10112 15385
rect 10594 15376 10600 15388
rect 10652 15376 10658 15428
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12713 15419 12771 15425
rect 12308 15388 12664 15416
rect 12308 15376 12314 15388
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5592 15320 5641 15348
rect 5592 15308 5598 15320
rect 5629 15317 5641 15320
rect 5675 15317 5687 15351
rect 5629 15311 5687 15317
rect 8665 15351 8723 15357
rect 8665 15317 8677 15351
rect 8711 15317 8723 15351
rect 8665 15311 8723 15317
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11882 15348 11888 15360
rect 10928 15320 11888 15348
rect 10928 15308 10934 15320
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12434 15348 12440 15360
rect 12115 15320 12440 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12636 15348 12664 15388
rect 12713 15385 12725 15419
rect 12759 15416 12771 15419
rect 14277 15419 14335 15425
rect 12759 15388 13400 15416
rect 12759 15385 12771 15388
rect 12713 15379 12771 15385
rect 12894 15348 12900 15360
rect 12636 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 13044 15320 13093 15348
rect 13044 15308 13050 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13372 15348 13400 15388
rect 14277 15385 14289 15419
rect 14323 15416 14335 15419
rect 14734 15416 14740 15428
rect 14323 15388 14740 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 13446 15348 13452 15360
rect 13372 15320 13452 15348
rect 13081 15311 13139 15317
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 14936 15348 14964 15447
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 16666 15493 16672 15496
rect 16660 15484 16672 15493
rect 16627 15456 16672 15484
rect 16660 15447 16672 15456
rect 16724 15484 16730 15496
rect 16942 15484 16948 15496
rect 16724 15456 16948 15484
rect 16666 15444 16672 15447
rect 16724 15444 16730 15456
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 18230 15484 18236 15496
rect 18191 15456 18236 15484
rect 18230 15444 18236 15456
rect 18288 15444 18294 15496
rect 18322 15444 18328 15496
rect 18380 15484 18386 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18380 15456 18705 15484
rect 18380 15444 18386 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 19610 15484 19616 15496
rect 19571 15456 19616 15484
rect 18693 15447 18751 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15484 19947 15487
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 19935 15456 20821 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 20809 15453 20821 15456
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 21177 15487 21235 15493
rect 21177 15453 21189 15487
rect 21223 15453 21235 15487
rect 21177 15447 21235 15453
rect 15378 15416 15384 15428
rect 15291 15388 15384 15416
rect 15378 15376 15384 15388
rect 15436 15416 15442 15428
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 15436 15388 15945 15416
rect 15436 15376 15442 15388
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 17494 15416 17500 15428
rect 15933 15379 15991 15385
rect 16040 15388 17500 15416
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 14936 15320 15485 15348
rect 15473 15317 15485 15320
rect 15519 15348 15531 15351
rect 16040 15348 16068 15388
rect 17494 15376 17500 15388
rect 17552 15376 17558 15428
rect 18248 15416 18276 15444
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 18248 15388 20729 15416
rect 20717 15385 20729 15388
rect 20763 15416 20775 15419
rect 21192 15416 21220 15447
rect 20763 15388 21220 15416
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 15519 15320 16068 15348
rect 15519 15317 15531 15320
rect 15473 15311 15531 15317
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16209 15351 16267 15357
rect 16209 15348 16221 15351
rect 16172 15320 16221 15348
rect 16172 15308 16178 15320
rect 16209 15317 16221 15320
rect 16255 15317 16267 15351
rect 17770 15348 17776 15360
rect 17731 15320 17776 15348
rect 16209 15311 16267 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 18874 15348 18880 15360
rect 18835 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 20993 15351 21051 15357
rect 20993 15317 21005 15351
rect 21039 15348 21051 15351
rect 21082 15348 21088 15360
rect 21039 15320 21088 15348
rect 21039 15317 21051 15320
rect 20993 15311 21051 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 5626 15104 5632 15156
rect 5684 15144 5690 15156
rect 6914 15144 6920 15156
rect 5684 15116 6920 15144
rect 5684 15104 5690 15116
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 7524 15116 7941 15144
rect 7524 15104 7530 15116
rect 7929 15113 7941 15116
rect 7975 15144 7987 15147
rect 8110 15144 8116 15156
rect 7975 15116 8116 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9122 15144 9128 15156
rect 9079 15116 9128 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9398 15104 9404 15156
rect 9456 15144 9462 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 9456 15116 9505 15144
rect 9456 15104 9462 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9493 15107 9551 15113
rect 9582 15104 9588 15156
rect 9640 15144 9646 15156
rect 9953 15147 10011 15153
rect 9640 15116 9685 15144
rect 9640 15104 9646 15116
rect 9953 15113 9965 15147
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 3050 15076 3056 15088
rect 2608 15048 3056 15076
rect 2608 15017 2636 15048
rect 3050 15036 3056 15048
rect 3108 15036 3114 15088
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 7742 15076 7748 15088
rect 3200 15048 7748 15076
rect 3200 15036 3206 15048
rect 7742 15036 7748 15048
rect 7800 15036 7806 15088
rect 8665 15079 8723 15085
rect 8665 15045 8677 15079
rect 8711 15076 8723 15079
rect 9968 15076 9996 15107
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11296 15116 11529 15144
rect 11296 15104 11302 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 11977 15147 12035 15153
rect 11977 15144 11989 15147
rect 11940 15116 11989 15144
rect 11940 15104 11946 15116
rect 11977 15113 11989 15116
rect 12023 15113 12035 15147
rect 11977 15107 12035 15113
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13035 15116 13461 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13906 15144 13912 15156
rect 13867 15116 13912 15144
rect 13449 15107 13507 15113
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 16485 15147 16543 15153
rect 16485 15113 16497 15147
rect 16531 15144 16543 15147
rect 16574 15144 16580 15156
rect 16531 15116 16580 15144
rect 16531 15113 16543 15116
rect 16485 15107 16543 15113
rect 16574 15104 16580 15116
rect 16632 15144 16638 15156
rect 16942 15144 16948 15156
rect 16632 15116 16948 15144
rect 16632 15104 16638 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17126 15144 17132 15156
rect 17087 15116 17132 15144
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 10410 15076 10416 15088
rect 8711 15048 9996 15076
rect 10323 15048 10416 15076
rect 8711 15045 8723 15048
rect 8665 15039 8723 15045
rect 10410 15036 10416 15048
rect 10468 15076 10474 15088
rect 11333 15079 11391 15085
rect 11333 15076 11345 15079
rect 10468 15048 11345 15076
rect 10468 15036 10474 15048
rect 11333 15045 11345 15048
rect 11379 15076 11391 15079
rect 16206 15076 16212 15088
rect 11379 15048 16212 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 16298 15036 16304 15088
rect 16356 15076 16362 15088
rect 16669 15079 16727 15085
rect 16669 15076 16681 15079
rect 16356 15048 16681 15076
rect 16356 15036 16362 15048
rect 16669 15045 16681 15048
rect 16715 15076 16727 15079
rect 17488 15079 17546 15085
rect 16715 15048 17264 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 1995 14980 2237 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 2860 15011 2918 15017
rect 2860 14977 2872 15011
rect 2906 15008 2918 15011
rect 2906 14980 3832 15008
rect 2906 14977 2918 14980
rect 2860 14971 2918 14977
rect 2516 14804 2544 14971
rect 3804 14872 3832 14980
rect 3970 14968 3976 15020
rect 4028 15008 4034 15020
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 4028 14980 4445 15008
rect 4028 14968 4034 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 5166 15008 5172 15020
rect 4571 14980 5172 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 15008 5411 15011
rect 5626 15008 5632 15020
rect 5399 14980 5632 15008
rect 5399 14977 5411 14980
rect 5353 14971 5411 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 6822 15008 6828 15020
rect 6779 14980 6828 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 6822 14968 6828 14980
rect 6880 15008 6886 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6880 14980 7389 15008
rect 6880 14968 6886 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 10321 15011 10379 15017
rect 7377 14971 7435 14977
rect 7484 14980 10180 15008
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 4617 14943 4675 14949
rect 4617 14940 4629 14943
rect 3936 14912 4629 14940
rect 3936 14900 3942 14912
rect 3988 14881 4016 14912
rect 4617 14909 4629 14912
rect 4663 14909 4675 14943
rect 5442 14940 5448 14952
rect 5403 14912 5448 14940
rect 4617 14903 4675 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 6917 14943 6975 14949
rect 5592 14912 5637 14940
rect 5592 14900 5598 14912
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7006 14940 7012 14952
rect 6963 14912 7012 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 7006 14900 7012 14912
rect 7064 14940 7070 14952
rect 7484 14949 7512 14980
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7064 14912 7481 14940
rect 7064 14900 7070 14912
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7834 14940 7840 14952
rect 7699 14912 7840 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 8386 14940 8392 14952
rect 8347 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14900 8450 14952
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14940 8631 14943
rect 9582 14940 9588 14952
rect 8619 14912 9588 14940
rect 8619 14909 8631 14912
rect 8573 14903 8631 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 3973 14875 4031 14881
rect 3804 14844 3924 14872
rect 2774 14804 2780 14816
rect 2516 14776 2780 14804
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 3896 14804 3924 14844
rect 3973 14841 3985 14875
rect 4019 14841 4031 14875
rect 3973 14835 4031 14841
rect 6362 14832 6368 14884
rect 6420 14872 6426 14884
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 6420 14844 6561 14872
rect 6420 14832 6426 14844
rect 6549 14841 6561 14844
rect 6595 14872 6607 14875
rect 7282 14872 7288 14884
rect 6595 14844 7288 14872
rect 6595 14841 6607 14844
rect 6549 14835 6607 14841
rect 7282 14832 7288 14844
rect 7340 14832 7346 14884
rect 7374 14832 7380 14884
rect 7432 14872 7438 14884
rect 9692 14872 9720 14903
rect 10042 14872 10048 14884
rect 7432 14844 10048 14872
rect 7432 14832 7438 14844
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 4338 14804 4344 14816
rect 3896 14776 4344 14804
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4985 14807 5043 14813
rect 4985 14804 4997 14807
rect 4580 14776 4997 14804
rect 4580 14764 4586 14776
rect 4985 14773 4997 14776
rect 5031 14773 5043 14807
rect 7006 14804 7012 14816
rect 6967 14776 7012 14804
rect 4985 14767 5043 14773
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 8662 14804 8668 14816
rect 8251 14776 8668 14804
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9398 14804 9404 14816
rect 9171 14776 9404 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 10152 14804 10180 14980
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10367 14980 10793 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 11882 15008 11888 15020
rect 11843 14980 11888 15008
rect 10781 14971 10839 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14918 15008 14924 15020
rect 14879 14980 14924 15008
rect 14918 14968 14924 14980
rect 14976 14968 14982 15020
rect 15372 15011 15430 15017
rect 15372 14977 15384 15011
rect 15418 15008 15430 15011
rect 16390 15008 16396 15020
rect 15418 14980 16396 15008
rect 15418 14977 15430 14980
rect 15372 14971 15430 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17236 15017 17264 15048
rect 17488 15045 17500 15079
rect 17534 15076 17546 15079
rect 17770 15076 17776 15088
rect 17534 15048 17776 15076
rect 17534 15045 17546 15048
rect 17488 15039 17546 15045
rect 17770 15036 17776 15048
rect 17828 15036 17834 15088
rect 19978 15076 19984 15088
rect 19939 15048 19984 15076
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17310 15008 17316 15020
rect 17267 14980 17316 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 17310 14968 17316 14980
rect 17368 15008 17374 15020
rect 18693 15011 18751 15017
rect 18693 15008 18705 15011
rect 17368 14980 18705 15008
rect 17368 14968 17374 14980
rect 18693 14977 18705 14980
rect 18739 15008 18751 15011
rect 18874 15008 18880 15020
rect 18739 14980 18880 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 19702 15008 19708 15020
rect 19663 14980 19708 15008
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 10594 14940 10600 14952
rect 10555 14912 10600 14940
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 11054 14940 11060 14952
rect 11015 14912 11060 14940
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 10612 14872 10640 14900
rect 12084 14872 12112 14903
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 12713 14943 12771 14949
rect 12713 14940 12725 14943
rect 12584 14912 12725 14940
rect 12584 14900 12590 14912
rect 12713 14909 12725 14912
rect 12759 14909 12771 14943
rect 12894 14940 12900 14952
rect 12855 14912 12900 14940
rect 12713 14903 12771 14909
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14274 14940 14280 14952
rect 14139 14912 14280 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14516 14912 15117 14940
rect 14516 14900 14522 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 14737 14875 14795 14881
rect 14737 14872 14749 14875
rect 10612 14844 12112 14872
rect 12176 14844 14749 14872
rect 12176 14804 12204 14844
rect 14737 14841 14749 14844
rect 14783 14841 14795 14875
rect 19794 14872 19800 14884
rect 14737 14835 14795 14841
rect 18156 14844 19800 14872
rect 12434 14804 12440 14816
rect 10152 14776 12204 14804
rect 12395 14776 12440 14804
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 13354 14804 13360 14816
rect 13315 14776 13360 14804
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 14752 14804 14780 14835
rect 15838 14804 15844 14816
rect 14752 14776 15844 14804
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 17218 14804 17224 14816
rect 16264 14776 17224 14804
rect 16264 14764 16270 14776
rect 17218 14764 17224 14776
rect 17276 14804 17282 14816
rect 18156 14804 18184 14844
rect 19794 14832 19800 14844
rect 19852 14832 19858 14884
rect 17276 14776 18184 14804
rect 17276 14764 17282 14776
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 18601 14807 18659 14813
rect 18601 14804 18613 14807
rect 18288 14776 18613 14804
rect 18288 14764 18294 14776
rect 18601 14773 18613 14776
rect 18647 14773 18659 14807
rect 18601 14767 18659 14773
rect 21085 14807 21143 14813
rect 21085 14773 21097 14807
rect 21131 14804 21143 14807
rect 21174 14804 21180 14816
rect 21131 14776 21180 14804
rect 21131 14773 21143 14776
rect 21085 14767 21143 14773
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 2866 14600 2872 14612
rect 2827 14572 2872 14600
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3252 14572 4169 14600
rect 1578 14532 1584 14544
rect 1539 14504 1584 14532
rect 1578 14492 1584 14504
rect 1636 14492 1642 14544
rect 2774 14492 2780 14544
rect 2832 14532 2838 14544
rect 3252 14532 3280 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 5718 14600 5724 14612
rect 4157 14563 4215 14569
rect 4632 14572 5724 14600
rect 2832 14504 3280 14532
rect 2832 14492 2838 14504
rect 3326 14492 3332 14544
rect 3384 14532 3390 14544
rect 3605 14535 3663 14541
rect 3605 14532 3617 14535
rect 3384 14504 3617 14532
rect 3384 14492 3390 14504
rect 3605 14501 3617 14504
rect 3651 14532 3663 14535
rect 4062 14532 4068 14544
rect 3651 14504 4068 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2590 14464 2596 14476
rect 2179 14436 2596 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 4632 14473 4660 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 9858 14600 9864 14612
rect 7800 14572 9720 14600
rect 9819 14572 9864 14600
rect 7800 14560 7806 14572
rect 9582 14492 9588 14544
rect 9640 14492 9646 14544
rect 9692 14532 9720 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 11882 14600 11888 14612
rect 10735 14572 11888 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12526 14600 12532 14612
rect 12207 14572 12532 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 15194 14600 15200 14612
rect 14056 14572 15200 14600
rect 14056 14560 14062 14572
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 19337 14603 19395 14609
rect 19337 14569 19349 14603
rect 19383 14600 19395 14603
rect 19978 14600 19984 14612
rect 19383 14572 19984 14600
rect 19383 14569 19395 14572
rect 19337 14563 19395 14569
rect 19978 14560 19984 14572
rect 20036 14600 20042 14612
rect 20898 14600 20904 14612
rect 20036 14572 20904 14600
rect 20036 14560 20042 14572
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21358 14600 21364 14612
rect 21319 14572 21364 14600
rect 21358 14560 21364 14572
rect 21416 14560 21422 14612
rect 15473 14535 15531 14541
rect 9692 14504 10272 14532
rect 4617 14467 4675 14473
rect 2700 14436 3464 14464
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14365 1823 14399
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 1765 14359 1823 14365
rect 1780 14328 1808 14359
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2700 14405 2728 14436
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3142 14396 3148 14408
rect 3099 14368 3148 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3436 14340 3464 14436
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 4617 14427 4675 14433
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 4982 14464 4988 14476
rect 4847 14436 4988 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 6362 14464 6368 14476
rect 6323 14436 6368 14464
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8036 14436 8585 14464
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6098 14399 6156 14405
rect 6098 14396 6110 14399
rect 5592 14368 6110 14396
rect 5592 14356 5598 14368
rect 6098 14365 6110 14368
rect 6144 14365 6156 14399
rect 6098 14359 6156 14365
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7929 14399 7987 14405
rect 7929 14396 7941 14399
rect 7340 14368 7941 14396
rect 7340 14356 7346 14368
rect 7929 14365 7941 14368
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 3326 14328 3332 14340
rect 1780 14300 3332 14328
rect 3326 14288 3332 14300
rect 3384 14288 3390 14340
rect 3418 14288 3424 14340
rect 3476 14328 3482 14340
rect 7684 14331 7742 14337
rect 3476 14300 3521 14328
rect 3476 14288 3482 14300
rect 7684 14297 7696 14331
rect 7730 14328 7742 14331
rect 7834 14328 7840 14340
rect 7730 14300 7840 14328
rect 7730 14297 7742 14300
rect 7684 14291 7742 14297
rect 7834 14288 7840 14300
rect 7892 14328 7898 14340
rect 8036 14328 8064 14436
rect 8573 14433 8585 14436
rect 8619 14433 8631 14467
rect 9214 14464 9220 14476
rect 9175 14436 9220 14464
rect 8573 14427 8631 14433
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9398 14464 9404 14476
rect 9359 14436 9404 14464
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 9600 14464 9628 14492
rect 9858 14464 9864 14476
rect 9600 14436 9864 14464
rect 9858 14424 9864 14436
rect 9916 14424 9922 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10244 14473 10272 14504
rect 15473 14501 15485 14535
rect 15519 14532 15531 14535
rect 20993 14535 21051 14541
rect 15519 14504 17264 14532
rect 15519 14501 15531 14504
rect 15473 14495 15531 14501
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 10318 14464 10324 14476
rect 10275 14436 10324 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 13872 14436 13921 14464
rect 13872 14424 13878 14436
rect 13909 14433 13921 14436
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14433 15715 14467
rect 15838 14464 15844 14476
rect 15799 14436 15844 14464
rect 15657 14427 15715 14433
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8168 14368 8401 14396
rect 8168 14356 8174 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14396 8539 14399
rect 8662 14396 8668 14408
rect 8527 14368 8668 14396
rect 8527 14365 8539 14368
rect 8481 14359 8539 14365
rect 7892 14300 8064 14328
rect 8404 14328 8432 14359
rect 8662 14356 8668 14368
rect 8720 14396 8726 14408
rect 9582 14396 9588 14408
rect 8720 14368 9588 14396
rect 8720 14356 8726 14368
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 12526 14405 12532 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 10560 14368 10793 14396
rect 10560 14356 10566 14368
rect 10781 14365 10793 14368
rect 10827 14396 10839 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 10827 14368 12265 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12520 14396 12532 14405
rect 12487 14368 12532 14396
rect 12253 14359 12311 14365
rect 12520 14359 12532 14368
rect 10686 14328 10692 14340
rect 8404 14300 10692 14328
rect 7892 14288 7898 14300
rect 9646 14272 9674 14300
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 11054 14337 11060 14340
rect 11048 14291 11060 14337
rect 11112 14328 11118 14340
rect 12268 14328 12296 14359
rect 12526 14356 12532 14359
rect 12584 14356 12590 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 12636 14368 14105 14396
rect 12434 14328 12440 14340
rect 11112 14300 11148 14328
rect 12268 14300 12440 14328
rect 11054 14288 11060 14291
rect 11112 14288 11118 14300
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 12636 14328 12664 14368
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14642 14396 14648 14408
rect 14139 14368 14648 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15672 14396 15700 14427
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 16574 14464 16580 14476
rect 16535 14436 16580 14464
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 15930 14396 15936 14408
rect 15672 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 14338 14331 14396 14337
rect 14338 14328 14350 14331
rect 12492 14300 12664 14328
rect 13648 14300 14350 14328
rect 12492 14288 12498 14300
rect 2498 14260 2504 14272
rect 2459 14232 2504 14260
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 3970 14260 3976 14272
rect 3931 14232 3976 14260
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 4982 14260 4988 14272
rect 4943 14232 4988 14260
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 5868 14232 6561 14260
rect 5868 14220 5874 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6549 14223 6607 14229
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 6788 14232 8033 14260
rect 6788 14220 6794 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8938 14260 8944 14272
rect 8899 14232 8944 14260
rect 8021 14223 8079 14229
rect 8938 14220 8944 14232
rect 8996 14260 9002 14272
rect 9493 14263 9551 14269
rect 9493 14260 9505 14263
rect 8996 14232 9505 14260
rect 8996 14220 9002 14232
rect 9493 14229 9505 14232
rect 9539 14229 9551 14263
rect 9646 14232 9680 14272
rect 9493 14223 9551 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10321 14263 10379 14269
rect 10321 14229 10333 14263
rect 10367 14260 10379 14263
rect 10870 14260 10876 14272
rect 10367 14232 10876 14260
rect 10367 14229 10379 14232
rect 10321 14223 10379 14229
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13648 14269 13676 14300
rect 14338 14297 14350 14300
rect 14384 14297 14396 14331
rect 14338 14291 14396 14297
rect 16669 14331 16727 14337
rect 16669 14297 16681 14331
rect 16715 14328 16727 14331
rect 17034 14328 17040 14340
rect 16715 14300 17040 14328
rect 16715 14297 16727 14300
rect 16669 14291 16727 14297
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 17236 14328 17264 14504
rect 20993 14501 21005 14535
rect 21039 14532 21051 14535
rect 21082 14532 21088 14544
rect 21039 14504 21088 14532
rect 21039 14501 21051 14504
rect 20993 14495 21051 14501
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 17310 14424 17316 14476
rect 17368 14464 17374 14476
rect 17586 14464 17592 14476
rect 17368 14436 17592 14464
rect 17368 14424 17374 14436
rect 17586 14424 17592 14436
rect 17644 14464 17650 14476
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 17644 14436 17693 14464
rect 17644 14424 17650 14436
rect 17681 14433 17693 14436
rect 17727 14433 17739 14467
rect 17681 14427 17739 14433
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 20717 14399 20775 14405
rect 20717 14396 20729 14399
rect 18472 14368 20729 14396
rect 18472 14356 18478 14368
rect 20717 14365 20729 14368
rect 20763 14396 20775 14399
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20763 14368 20821 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 21174 14396 21180 14408
rect 21135 14368 21180 14396
rect 20809 14359 20867 14365
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 17310 14328 17316 14340
rect 17236 14300 17316 14328
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17948 14331 18006 14337
rect 17948 14297 17960 14331
rect 17994 14328 18006 14331
rect 18138 14328 18144 14340
rect 17994 14300 18144 14328
rect 17994 14297 18006 14300
rect 17948 14291 18006 14297
rect 18138 14288 18144 14300
rect 18196 14288 18202 14340
rect 18690 14288 18696 14340
rect 18748 14328 18754 14340
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 18748 14300 19441 14328
rect 18748 14288 18754 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 12860 14232 13645 14260
rect 12860 14220 12866 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15654 14260 15660 14272
rect 14976 14232 15660 14260
rect 14976 14220 14982 14232
rect 15654 14220 15660 14232
rect 15712 14260 15718 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15712 14232 15945 14260
rect 15712 14220 15718 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 16298 14260 16304 14272
rect 16259 14232 16304 14260
rect 15933 14223 15991 14229
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 16761 14263 16819 14269
rect 16761 14229 16773 14263
rect 16807 14260 16819 14263
rect 16942 14260 16948 14272
rect 16807 14232 16948 14260
rect 16807 14229 16819 14232
rect 16761 14223 16819 14229
rect 16942 14220 16948 14232
rect 17000 14220 17006 14272
rect 17129 14263 17187 14269
rect 17129 14229 17141 14263
rect 17175 14260 17187 14263
rect 17770 14260 17776 14272
rect 17175 14232 17776 14260
rect 17175 14229 17187 14232
rect 17129 14223 17187 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 18840 14232 19073 14260
rect 18840 14220 18846 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 19061 14223 19119 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 1728 14028 3617 14056
rect 1728 14016 1734 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5592 14028 5917 14056
rect 5592 14016 5598 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 6546 14056 6552 14068
rect 5951 14028 6552 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6730 14056 6736 14068
rect 6691 14028 6736 14056
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7006 14056 7012 14068
rect 6871 14028 7012 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9858 14056 9864 14068
rect 9447 14028 9711 14056
rect 9819 14028 9864 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 2808 13991 2866 13997
rect 2808 13957 2820 13991
rect 2854 13988 2866 13991
rect 3050 13988 3056 14000
rect 2854 13960 3056 13988
rect 2854 13957 2866 13960
rect 2808 13951 2866 13957
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 3200 13960 3249 13988
rect 3200 13948 3206 13960
rect 3237 13957 3249 13960
rect 3283 13988 3295 13991
rect 3513 13991 3571 13997
rect 3513 13988 3525 13991
rect 3283 13960 3525 13988
rect 3283 13957 3295 13960
rect 3237 13951 3295 13957
rect 3513 13957 3525 13960
rect 3559 13988 3571 13991
rect 4154 13988 4160 14000
rect 3559 13960 4160 13988
rect 3559 13957 3571 13960
rect 3513 13951 3571 13957
rect 3053 13855 3111 13861
rect 3053 13821 3065 13855
rect 3099 13852 3111 13855
rect 3252 13852 3280 13951
rect 4154 13948 4160 13960
rect 4212 13988 4218 14000
rect 4212 13960 4568 13988
rect 4212 13948 4218 13960
rect 4540 13929 4568 13960
rect 4982 13948 4988 14000
rect 5040 13988 5046 14000
rect 7438 13991 7496 13997
rect 7438 13988 7450 13991
rect 5040 13960 7450 13988
rect 5040 13948 5046 13960
rect 7438 13957 7450 13960
rect 7484 13957 7496 13991
rect 7438 13951 7496 13957
rect 8941 13991 8999 13997
rect 8941 13957 8953 13991
rect 8987 13988 8999 13991
rect 9214 13988 9220 14000
rect 8987 13960 9220 13988
rect 8987 13957 8999 13960
rect 8941 13951 8999 13957
rect 9214 13948 9220 13960
rect 9272 13948 9278 14000
rect 9493 13991 9551 13997
rect 9493 13988 9505 13991
rect 9416 13960 9505 13988
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 4525 13923 4583 13929
rect 4019 13892 4476 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 4062 13852 4068 13864
rect 3099 13824 3280 13852
rect 4023 13824 4068 13852
rect 3099 13821 3111 13824
rect 3053 13815 3111 13821
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4172 13784 4200 13815
rect 4028 13756 4200 13784
rect 4028 13744 4034 13756
rect 1673 13719 1731 13725
rect 1673 13685 1685 13719
rect 1719 13716 1731 13719
rect 1946 13716 1952 13728
rect 1719 13688 1952 13716
rect 1719 13685 1731 13688
rect 1673 13679 1731 13685
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 4448 13716 4476 13892
rect 4525 13889 4537 13923
rect 4571 13889 4583 13923
rect 4525 13883 4583 13889
rect 4792 13923 4850 13929
rect 4792 13889 4804 13923
rect 4838 13920 4850 13923
rect 5810 13920 5816 13932
rect 4838 13892 5816 13920
rect 4838 13889 4850 13892
rect 4792 13883 4850 13889
rect 5810 13880 5816 13892
rect 5868 13920 5874 13932
rect 7193 13923 7251 13929
rect 5868 13892 6132 13920
rect 5868 13880 5874 13892
rect 5994 13852 6000 13864
rect 5955 13824 6000 13852
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6104 13852 6132 13892
rect 7193 13889 7205 13923
rect 7239 13920 7251 13923
rect 7282 13920 7288 13932
rect 7239 13892 7288 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 6822 13852 6828 13864
rect 6104 13824 6828 13852
rect 6822 13812 6828 13824
rect 6880 13852 6886 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6880 13824 6929 13852
rect 6880 13812 6886 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 9416 13852 9444 13960
rect 9493 13957 9505 13960
rect 9539 13957 9551 13991
rect 9493 13951 9551 13957
rect 9683 13920 9711 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10376 14028 10977 14056
rect 10376 14016 10382 14028
rect 10965 14025 10977 14028
rect 11011 14056 11023 14059
rect 11330 14056 11336 14068
rect 11011 14028 11336 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 12952 14028 13369 14056
rect 12952 14016 12958 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 16669 14059 16727 14065
rect 13504 14028 13549 14056
rect 13504 14016 13510 14028
rect 16669 14025 16681 14059
rect 16715 14056 16727 14059
rect 17034 14056 17040 14068
rect 16715 14028 17040 14056
rect 16715 14025 16727 14028
rect 16669 14019 16727 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17770 14056 17776 14068
rect 17731 14028 17776 14056
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 18233 14059 18291 14065
rect 17920 14028 17965 14056
rect 17920 14016 17926 14028
rect 18233 14025 18245 14059
rect 18279 14025 18291 14059
rect 18233 14019 18291 14025
rect 19337 14059 19395 14065
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19797 14059 19855 14065
rect 19797 14056 19809 14059
rect 19383 14028 19809 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19797 14025 19809 14028
rect 19843 14025 19855 14059
rect 19797 14019 19855 14025
rect 20993 14059 21051 14065
rect 20993 14025 21005 14059
rect 21039 14056 21051 14059
rect 21082 14056 21088 14068
rect 21039 14028 21088 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 10042 13948 10048 14000
rect 10100 13988 10106 14000
rect 10229 13991 10287 13997
rect 10229 13988 10241 13991
rect 10100 13960 10241 13988
rect 10100 13948 10106 13960
rect 10229 13957 10241 13960
rect 10275 13957 10287 13991
rect 10229 13951 10287 13957
rect 12345 13991 12403 13997
rect 12345 13957 12357 13991
rect 12391 13988 12403 13991
rect 13817 13991 13875 13997
rect 12391 13960 13124 13988
rect 12391 13957 12403 13960
rect 12345 13951 12403 13957
rect 11514 13920 11520 13932
rect 9683 13892 11520 13920
rect 11514 13880 11520 13892
rect 11572 13920 11578 13932
rect 12066 13920 12072 13932
rect 11572 13892 12072 13920
rect 11572 13880 11578 13892
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12452 13892 13001 13920
rect 12452 13864 12480 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 9490 13852 9496 13864
rect 9416 13824 9496 13852
rect 6917 13815 6975 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9640 13824 9689 13852
rect 9640 13812 9646 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 10321 13855 10379 13861
rect 10321 13852 10333 13855
rect 9916 13824 10333 13852
rect 9916 13812 9922 13824
rect 10321 13821 10333 13824
rect 10367 13821 10379 13855
rect 10321 13815 10379 13821
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10594 13852 10600 13864
rect 10551 13824 10600 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10870 13852 10876 13864
rect 10831 13824 10876 13852
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11790 13852 11796 13864
rect 11112 13824 11796 13852
rect 11112 13812 11118 13824
rect 11790 13812 11796 13824
rect 11848 13852 11854 13864
rect 11848 13824 12388 13852
rect 11848 13812 11854 13824
rect 7006 13784 7012 13796
rect 6196 13756 7012 13784
rect 6196 13716 6224 13756
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 8573 13787 8631 13793
rect 8573 13753 8585 13787
rect 8619 13784 8631 13787
rect 8619 13756 9260 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 9232 13728 9260 13756
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 11606 13784 11612 13796
rect 11296 13756 11612 13784
rect 11296 13744 11302 13756
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 12360 13784 12388 13824
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12805 13855 12863 13861
rect 12492 13824 12537 13852
rect 12492 13812 12498 13824
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13096 13852 13124 13960
rect 13817 13957 13829 13991
rect 13863 13988 13875 13991
rect 13863 13960 14780 13988
rect 13863 13957 13875 13960
rect 13817 13951 13875 13957
rect 14752 13929 14780 13960
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 17129 13991 17187 13997
rect 17129 13988 17141 13991
rect 16356 13960 17141 13988
rect 16356 13948 16362 13960
rect 17129 13957 17141 13960
rect 17175 13957 17187 13991
rect 18248 13988 18276 14019
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 19610 13988 19616 14000
rect 18248 13960 19616 13988
rect 17129 13951 17187 13957
rect 19610 13948 19616 13960
rect 19668 13948 19674 14000
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14737 13923 14795 13929
rect 13955 13892 14596 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14568 13864 14596 13892
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 15378 13920 15384 13932
rect 14783 13892 15384 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15930 13880 15936 13932
rect 15988 13929 15994 13932
rect 15988 13920 16000 13929
rect 15988 13892 16033 13920
rect 15988 13883 16000 13892
rect 15988 13880 15994 13883
rect 16850 13880 16856 13932
rect 16908 13920 16914 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16908 13892 17049 13920
rect 16908 13880 16914 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 18966 13920 18972 13932
rect 18927 13892 18972 13920
rect 17037 13883 17095 13889
rect 18966 13880 18972 13892
rect 19024 13880 19030 13932
rect 19518 13880 19524 13932
rect 19576 13920 19582 13932
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 19576 13892 19901 13920
rect 19576 13880 19582 13892
rect 19889 13889 19901 13892
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 13998 13852 14004 13864
rect 12943 13824 14004 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 12820 13784 12848 13815
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13852 14151 13855
rect 14274 13852 14280 13864
rect 14139 13824 14280 13852
rect 14139 13821 14151 13824
rect 14093 13815 14151 13821
rect 14108 13784 14136 13815
rect 14274 13812 14280 13824
rect 14332 13812 14338 13864
rect 14550 13852 14556 13864
rect 14511 13824 14556 13852
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 15194 13852 15200 13864
rect 14844 13824 15200 13852
rect 12360 13756 14136 13784
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13784 14427 13787
rect 14642 13784 14648 13796
rect 14415 13756 14648 13784
rect 14415 13753 14427 13756
rect 14369 13747 14427 13753
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 14844 13793 14872 13824
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 16209 13855 16267 13861
rect 16209 13821 16221 13855
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 17221 13855 17279 13861
rect 17221 13821 17233 13855
rect 17267 13821 17279 13855
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 17221 13815 17279 13821
rect 14829 13787 14887 13793
rect 14829 13753 14841 13787
rect 14875 13753 14887 13787
rect 14829 13747 14887 13753
rect 16224 13728 16252 13815
rect 16390 13744 16396 13796
rect 16448 13784 16454 13796
rect 17236 13784 17264 13815
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 17828 13824 18337 13852
rect 17828 13812 17834 13824
rect 18325 13821 18337 13824
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 18693 13855 18751 13861
rect 18693 13821 18705 13855
rect 18739 13821 18751 13855
rect 18874 13852 18880 13864
rect 18835 13824 18880 13852
rect 18693 13815 18751 13821
rect 16448 13756 17264 13784
rect 18708 13784 18736 13815
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 19702 13852 19708 13864
rect 19444 13824 19708 13852
rect 19058 13784 19064 13796
rect 18708 13756 19064 13784
rect 16448 13744 16454 13756
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 19444 13793 19472 13824
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13821 20039 13855
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 19981 13815 20039 13821
rect 20088 13824 20729 13852
rect 19429 13787 19487 13793
rect 19429 13753 19441 13787
rect 19475 13753 19487 13787
rect 19429 13747 19487 13753
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 19996 13784 20024 13815
rect 19852 13756 20024 13784
rect 19852 13744 19858 13756
rect 6362 13716 6368 13728
rect 4448 13688 6224 13716
rect 6323 13688 6368 13716
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8665 13719 8723 13725
rect 8665 13716 8677 13719
rect 8444 13688 8677 13716
rect 8444 13676 8450 13688
rect 8665 13685 8677 13688
rect 8711 13685 8723 13719
rect 8665 13679 8723 13685
rect 9033 13719 9091 13725
rect 9033 13685 9045 13719
rect 9079 13716 9091 13719
rect 9122 13716 9128 13728
rect 9079 13688 9128 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9214 13676 9220 13728
rect 9272 13676 9278 13728
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 11020 13688 11161 13716
rect 11020 13676 11026 13688
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 11149 13679 11207 13685
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 15838 13716 15844 13728
rect 12216 13688 15844 13716
rect 12216 13676 12222 13688
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 16264 13688 16313 13716
rect 16264 13676 16270 13688
rect 16301 13685 16313 13688
rect 16347 13685 16359 13719
rect 16301 13679 16359 13685
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 20088 13716 20116 13824
rect 20717 13821 20729 13824
rect 20763 13852 20775 13855
rect 20824 13852 20852 13883
rect 20763 13824 20852 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 18564 13688 20116 13716
rect 18564 13676 18570 13688
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 2314 13512 2320 13524
rect 2179 13484 2320 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 2314 13472 2320 13484
rect 2372 13472 2378 13524
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4341 13515 4399 13521
rect 4341 13512 4353 13515
rect 4304 13484 4353 13512
rect 4304 13472 4310 13484
rect 4341 13481 4353 13484
rect 4387 13481 4399 13515
rect 4341 13475 4399 13481
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5442 13512 5448 13524
rect 5215 13484 5448 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5776 13484 6009 13512
rect 5776 13472 5782 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7374 13512 7380 13524
rect 6963 13484 7380 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7374 13472 7380 13484
rect 7432 13512 7438 13524
rect 12158 13512 12164 13524
rect 7432 13484 12164 13512
rect 7432 13472 7438 13484
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 13722 13512 13728 13524
rect 13495 13484 13728 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 16390 13512 16396 13524
rect 15252 13484 16068 13512
rect 15252 13472 15258 13484
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 8021 13447 8079 13453
rect 8021 13444 8033 13447
rect 4120 13416 8033 13444
rect 4120 13404 4126 13416
rect 8021 13413 8033 13416
rect 8067 13413 8079 13447
rect 8021 13407 8079 13413
rect 8941 13447 8999 13453
rect 8941 13413 8953 13447
rect 8987 13413 8999 13447
rect 8941 13407 8999 13413
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13376 1639 13379
rect 1946 13376 1952 13388
rect 1627 13348 1952 13376
rect 1627 13345 1639 13348
rect 1581 13339 1639 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 3605 13379 3663 13385
rect 3605 13345 3617 13379
rect 3651 13376 3663 13379
rect 4154 13376 4160 13388
rect 3651 13348 4160 13376
rect 3651 13345 3663 13348
rect 3605 13339 3663 13345
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 3620 13308 3648 13339
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4893 13379 4951 13385
rect 4893 13376 4905 13379
rect 4396 13348 4905 13376
rect 4396 13336 4402 13348
rect 4893 13345 4905 13348
rect 4939 13345 4951 13379
rect 4893 13339 4951 13345
rect 5350 13336 5356 13388
rect 5408 13376 5414 13388
rect 5629 13379 5687 13385
rect 5629 13376 5641 13379
rect 5408 13348 5641 13376
rect 5408 13336 5414 13348
rect 5629 13345 5641 13348
rect 5675 13345 5687 13379
rect 5810 13376 5816 13388
rect 5771 13348 5816 13376
rect 5629 13339 5687 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 6420 13348 6469 13376
rect 6420 13336 6426 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6604 13348 6649 13376
rect 6604 13336 6610 13348
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7561 13379 7619 13385
rect 7561 13376 7573 13379
rect 6880 13348 7573 13376
rect 6880 13336 6886 13348
rect 7561 13345 7573 13348
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 8573 13379 8631 13385
rect 8573 13376 8585 13379
rect 7800 13348 8585 13376
rect 7800 13336 7806 13348
rect 8573 13345 8585 13348
rect 8619 13376 8631 13379
rect 8956 13376 8984 13407
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 15930 13444 15936 13456
rect 10376 13416 14596 13444
rect 15891 13416 15936 13444
rect 10376 13404 10382 13416
rect 9214 13376 9220 13388
rect 8619 13348 9220 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 9214 13336 9220 13348
rect 9272 13336 9278 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10235 13348 10977 13376
rect 2648 13280 3648 13308
rect 4172 13308 4200 13336
rect 4522 13308 4528 13320
rect 4172 13280 4528 13308
rect 2648 13268 2654 13280
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 7466 13308 7472 13320
rect 7427 13280 7472 13308
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13308 7987 13311
rect 8202 13308 8208 13320
rect 7975 13280 8208 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 9490 13308 9496 13320
rect 8435 13280 9496 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 10054 13311 10112 13317
rect 10054 13308 10066 13311
rect 9640 13280 10066 13308
rect 9640 13268 9646 13280
rect 10054 13277 10066 13280
rect 10100 13308 10112 13311
rect 10235 13308 10263 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 12802 13376 12808 13388
rect 12763 13348 12808 13376
rect 10965 13339 11023 13345
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 12986 13376 12992 13388
rect 12947 13348 12992 13376
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 13722 13376 13728 13388
rect 13679 13348 13728 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14568 13376 14596 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 16040 13444 16068 13484
rect 16224 13484 16396 13512
rect 16224 13444 16252 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16761 13515 16819 13521
rect 16761 13481 16773 13515
rect 16807 13512 16819 13515
rect 16942 13512 16948 13524
rect 16807 13484 16948 13512
rect 16807 13481 16819 13484
rect 16761 13475 16819 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 18932 13484 19257 13512
rect 18932 13472 18938 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 21450 13512 21456 13524
rect 21411 13484 21456 13512
rect 19245 13475 19303 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 16850 13444 16856 13456
rect 16040 13416 16252 13444
rect 16811 13416 16856 13444
rect 16224 13385 16252 13416
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 18966 13404 18972 13456
rect 19024 13444 19030 13456
rect 20073 13447 20131 13453
rect 20073 13444 20085 13447
rect 19024 13416 20085 13444
rect 19024 13404 19030 13416
rect 20073 13413 20085 13416
rect 20119 13413 20131 13447
rect 20073 13407 20131 13413
rect 16209 13379 16267 13385
rect 14568 13348 14688 13376
rect 10100 13280 10263 13308
rect 10321 13311 10379 13317
rect 10100 13277 10112 13280
rect 10054 13271 10112 13277
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 11146 13308 11152 13320
rect 10367 13280 11152 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13354 13308 13360 13320
rect 13127 13280 13360 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14660 13308 14688 13348
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 16209 13339 16267 13345
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16356 13348 16401 13376
rect 16356 13336 16362 13348
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17405 13379 17463 13385
rect 17405 13376 17417 13379
rect 17000 13348 17417 13376
rect 17000 13336 17006 13348
rect 17405 13345 17417 13348
rect 17451 13345 17463 13379
rect 17405 13339 17463 13345
rect 17586 13336 17592 13388
rect 17644 13376 17650 13388
rect 17681 13379 17739 13385
rect 17681 13376 17693 13379
rect 17644 13348 17693 13376
rect 17644 13336 17650 13348
rect 17681 13345 17693 13348
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 19797 13379 19855 13385
rect 19797 13345 19809 13379
rect 19843 13376 19855 13379
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 19843 13348 20637 13376
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 20625 13345 20637 13348
rect 20671 13345 20683 13379
rect 20625 13339 20683 13345
rect 17034 13308 17040 13320
rect 14660 13280 17040 13308
rect 14553 13271 14611 13277
rect 1765 13243 1823 13249
rect 1765 13209 1777 13243
rect 1811 13240 1823 13243
rect 3142 13240 3148 13252
rect 1811 13212 3148 13240
rect 1811 13209 1823 13212
rect 1765 13203 1823 13209
rect 3142 13200 3148 13212
rect 3200 13200 3206 13252
rect 3326 13240 3332 13252
rect 3384 13249 3390 13252
rect 3384 13243 3418 13249
rect 3270 13212 3332 13240
rect 3326 13200 3332 13212
rect 3406 13240 3418 13243
rect 4154 13240 4160 13252
rect 3406 13212 4160 13240
rect 3406 13209 3418 13212
rect 3384 13203 3418 13209
rect 3384 13200 3390 13203
rect 4154 13200 4160 13212
rect 4212 13200 4218 13252
rect 6365 13243 6423 13249
rect 6365 13209 6377 13243
rect 6411 13240 6423 13243
rect 7374 13240 7380 13252
rect 6411 13212 7052 13240
rect 7335 13212 7380 13240
rect 6411 13209 6423 13212
rect 6365 13203 6423 13209
rect 2225 13175 2283 13181
rect 2225 13141 2237 13175
rect 2271 13172 2283 13175
rect 3050 13172 3056 13184
rect 2271 13144 3056 13172
rect 2271 13141 2283 13144
rect 2225 13135 2283 13141
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3292 13144 3801 13172
rect 3292 13132 3298 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 4249 13175 4307 13181
rect 4249 13141 4261 13175
rect 4295 13172 4307 13175
rect 4338 13172 4344 13184
rect 4295 13144 4344 13172
rect 4295 13141 4307 13144
rect 4249 13135 4307 13141
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 4709 13175 4767 13181
rect 4709 13172 4721 13175
rect 4672 13144 4721 13172
rect 4672 13132 4678 13144
rect 4709 13141 4721 13144
rect 4755 13141 4767 13175
rect 4709 13135 4767 13141
rect 4801 13175 4859 13181
rect 4801 13141 4813 13175
rect 4847 13172 4859 13175
rect 5442 13172 5448 13184
rect 4847 13144 5448 13172
rect 4847 13141 4859 13144
rect 4801 13135 4859 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5592 13144 5637 13172
rect 5592 13132 5598 13144
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 6638 13172 6644 13184
rect 5868 13144 6644 13172
rect 5868 13132 5874 13144
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7024 13181 7052 13212
rect 7374 13200 7380 13212
rect 7432 13200 7438 13252
rect 8481 13243 8539 13249
rect 8481 13209 8493 13243
rect 8527 13240 8539 13243
rect 8527 13212 9260 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13141 7067 13175
rect 7009 13135 7067 13141
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 9030 13172 9036 13184
rect 7984 13144 9036 13172
rect 7984 13132 7990 13144
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 9232 13172 9260 13212
rect 10594 13200 10600 13252
rect 10652 13240 10658 13252
rect 10781 13243 10839 13249
rect 10781 13240 10793 13243
rect 10652 13212 10793 13240
rect 10652 13200 10658 13212
rect 10781 13209 10793 13212
rect 10827 13209 10839 13243
rect 13814 13240 13820 13252
rect 10781 13203 10839 13209
rect 11072 13212 13820 13240
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9232 13144 10425 13172
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13172 10931 13175
rect 11072 13172 11100 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14568 13240 14596 13271
rect 17034 13268 17040 13280
rect 17092 13308 17098 13320
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 17092 13280 17325 13308
rect 17092 13268 17098 13280
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17948 13311 18006 13317
rect 17948 13308 17960 13311
rect 17313 13271 17371 13277
rect 17880 13280 17960 13308
rect 17880 13252 17908 13280
rect 17948 13277 17960 13280
rect 17994 13308 18006 13311
rect 18782 13308 18788 13320
rect 17994 13280 18788 13308
rect 17994 13277 18006 13280
rect 17948 13271 18006 13277
rect 18782 13268 18788 13280
rect 18840 13308 18846 13320
rect 19812 13308 19840 13339
rect 20530 13308 20536 13320
rect 18840 13280 19840 13308
rect 20491 13280 20536 13308
rect 18840 13268 18846 13280
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 14642 13240 14648 13252
rect 14568 13212 14648 13240
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 14820 13243 14878 13249
rect 14820 13209 14832 13243
rect 14866 13240 14878 13243
rect 15194 13240 15200 13252
rect 14866 13212 15200 13240
rect 14866 13209 14878 13212
rect 14820 13203 14878 13209
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 15838 13200 15844 13252
rect 15896 13240 15902 13252
rect 16393 13243 16451 13249
rect 16393 13240 16405 13243
rect 15896 13212 16405 13240
rect 15896 13200 15902 13212
rect 16393 13209 16405 13212
rect 16439 13209 16451 13243
rect 16393 13203 16451 13209
rect 17221 13243 17279 13249
rect 17221 13209 17233 13243
rect 17267 13240 17279 13243
rect 17770 13240 17776 13252
rect 17267 13212 17776 13240
rect 17267 13209 17279 13212
rect 17221 13203 17279 13209
rect 17770 13200 17776 13212
rect 17828 13200 17834 13252
rect 17862 13200 17868 13252
rect 17920 13200 17926 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 18524 13212 19625 13240
rect 10919 13144 11100 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 11204 13144 11345 13172
rect 11204 13132 11210 13144
rect 11333 13141 11345 13144
rect 11379 13172 11391 13175
rect 12342 13172 12348 13184
rect 11379 13144 12348 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 18524 13172 18552 13212
rect 19613 13209 19625 13212
rect 19659 13240 19671 13243
rect 19978 13240 19984 13252
rect 19659 13212 19984 13240
rect 19659 13209 19671 13212
rect 19613 13203 19671 13209
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 14792 13144 18552 13172
rect 14792 13132 14798 13144
rect 18966 13132 18972 13184
rect 19024 13172 19030 13184
rect 19061 13175 19119 13181
rect 19061 13172 19073 13175
rect 19024 13144 19073 13172
rect 19024 13132 19030 13144
rect 19061 13141 19073 13144
rect 19107 13141 19119 13175
rect 19702 13172 19708 13184
rect 19663 13144 19708 13172
rect 19061 13135 19119 13141
rect 19702 13132 19708 13144
rect 19760 13172 19766 13184
rect 20162 13172 20168 13184
rect 19760 13144 20168 13172
rect 19760 13132 19766 13144
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 20438 13172 20444 13184
rect 20399 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3970 12968 3976 12980
rect 3108 12940 3976 12968
rect 3108 12928 3114 12940
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 5626 12968 5632 12980
rect 5587 12940 5632 12968
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 7282 12968 7288 12980
rect 6135 12940 7288 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 1946 12860 1952 12912
rect 2004 12900 2010 12912
rect 2838 12903 2896 12909
rect 2838 12900 2850 12903
rect 2004 12872 2850 12900
rect 2004 12860 2010 12872
rect 2838 12869 2850 12872
rect 2884 12869 2896 12903
rect 2838 12863 2896 12869
rect 4706 12860 4712 12912
rect 4764 12900 4770 12912
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 4764 12872 5181 12900
rect 4764 12860 4770 12872
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 5261 12903 5319 12909
rect 5261 12869 5273 12903
rect 5307 12900 5319 12903
rect 5994 12900 6000 12912
rect 5307 12872 6000 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 5994 12860 6000 12872
rect 6052 12860 6058 12912
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12832 1823 12835
rect 2041 12835 2099 12841
rect 2041 12832 2053 12835
rect 1811 12804 2053 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2041 12801 2053 12804
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2363 12804 3924 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3896 12696 3924 12804
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4120 12804 4445 12832
rect 4120 12792 4126 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 4890 12832 4896 12844
rect 4571 12804 4896 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5350 12792 5356 12844
rect 5408 12832 5414 12844
rect 6380 12841 6408 12940
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7524 12940 7849 12968
rect 7524 12928 7530 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 8294 12968 8300 12980
rect 8255 12940 8300 12968
rect 7837 12931 7895 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8665 12971 8723 12977
rect 8665 12937 8677 12971
rect 8711 12937 8723 12971
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 8665 12931 8723 12937
rect 6822 12900 6828 12912
rect 6472 12872 6828 12900
rect 5905 12835 5963 12841
rect 5905 12832 5917 12835
rect 5408 12804 5917 12832
rect 5408 12792 5414 12804
rect 5905 12801 5917 12804
rect 5951 12832 5963 12835
rect 6365 12835 6423 12841
rect 5951 12804 6316 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4304 12736 4629 12764
rect 4304 12724 4310 12736
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5718 12764 5724 12776
rect 5123 12736 5724 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 5994 12724 6000 12776
rect 6052 12724 6058 12776
rect 6288 12764 6316 12804
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6472 12764 6500 12872
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 8680 12900 8708 12931
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 9950 12928 9956 12940
rect 10008 12968 10014 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10008 12940 10701 12968
rect 10008 12928 10014 12940
rect 10689 12937 10701 12940
rect 10735 12968 10747 12971
rect 12526 12968 12532 12980
rect 10735 12940 12532 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 13722 12968 13728 12980
rect 13403 12940 13728 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 15838 12968 15844 12980
rect 15799 12940 15844 12968
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 17034 12968 17040 12980
rect 16807 12940 17040 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 17034 12928 17040 12940
rect 17092 12968 17098 12980
rect 17954 12968 17960 12980
rect 17092 12940 17960 12968
rect 17092 12928 17098 12940
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 19426 12968 19432 12980
rect 18279 12940 19432 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19576 12940 19717 12968
rect 19576 12928 19582 12940
rect 19705 12937 19717 12940
rect 19751 12968 19763 12971
rect 19794 12968 19800 12980
rect 19751 12940 19800 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20438 12968 20444 12980
rect 20027 12940 20444 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 7064 12872 8708 12900
rect 8772 12872 12756 12900
rect 7064 12860 7070 12872
rect 6638 12841 6644 12844
rect 6621 12835 6644 12841
rect 6621 12801 6633 12835
rect 6621 12795 6644 12801
rect 6638 12792 6644 12795
rect 6696 12792 6702 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7800 12804 8217 12832
rect 7800 12792 7806 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 7834 12764 7840 12776
rect 6288 12736 6500 12764
rect 7747 12736 7840 12764
rect 6012 12696 6040 12724
rect 7760 12705 7788 12736
rect 7834 12724 7840 12736
rect 7892 12764 7898 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 7892 12736 8401 12764
rect 7892 12724 7898 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 3896 12668 6040 12696
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12665 7803 12699
rect 7745 12659 7803 12665
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 3936 12600 3985 12628
rect 3936 12588 3942 12600
rect 3973 12597 3985 12600
rect 4019 12597 4031 12631
rect 3973 12591 4031 12597
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4246 12628 4252 12640
rect 4111 12600 4252 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 5442 12628 5448 12640
rect 5132 12600 5448 12628
rect 5132 12588 5138 12600
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 8772 12628 8800 12872
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9490 12832 9496 12844
rect 9079 12804 9496 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9858 12832 9864 12844
rect 9771 12804 9864 12832
rect 9858 12792 9864 12804
rect 9916 12832 9922 12844
rect 9916 12804 11008 12832
rect 9916 12792 9922 12804
rect 9214 12764 9220 12776
rect 9175 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9582 12724 9588 12776
rect 9640 12764 9646 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9640 12736 10057 12764
rect 9640 12724 9646 12736
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10192 12736 10333 12764
rect 10192 12724 10198 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 10336 12696 10364 12727
rect 10686 12696 10692 12708
rect 10336 12668 10692 12696
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 6788 12600 8800 12628
rect 6788 12588 6794 12600
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 10594 12628 10600 12640
rect 9088 12600 10600 12628
rect 9088 12588 9094 12600
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10980 12637 11008 12804
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11204 12804 11529 12832
rect 11204 12792 11210 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11784 12835 11842 12841
rect 11784 12801 11796 12835
rect 11830 12832 11842 12835
rect 12342 12832 12348 12844
rect 11830 12804 12348 12832
rect 11830 12801 11842 12804
rect 11784 12795 11842 12801
rect 12342 12792 12348 12804
rect 12400 12832 12406 12844
rect 12728 12832 12756 12872
rect 14642 12860 14648 12912
rect 14700 12900 14706 12912
rect 14700 12872 15424 12900
rect 14700 12860 14706 12872
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 12400 12804 12664 12832
rect 12728 12804 13921 12832
rect 12400 12792 12406 12804
rect 12636 12764 12664 12804
rect 13280 12773 13308 12804
rect 13909 12801 13921 12804
rect 13955 12832 13967 12835
rect 14734 12832 14740 12844
rect 13955 12804 14740 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 15396 12841 15424 12872
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 16942 12900 16948 12912
rect 15988 12872 16948 12900
rect 15988 12860 15994 12872
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 17126 12900 17132 12912
rect 17087 12872 17132 12900
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 17218 12860 17224 12912
rect 17276 12860 17282 12912
rect 18570 12903 18628 12909
rect 18570 12900 18582 12903
rect 17696 12872 18582 12900
rect 15114 12835 15172 12841
rect 15114 12832 15126 12835
rect 14884 12804 15126 12832
rect 14884 12792 14890 12804
rect 15114 12801 15126 12804
rect 15160 12801 15172 12835
rect 15114 12795 15172 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12832 15439 12835
rect 15427 12804 15516 12832
rect 15427 12801 15439 12804
rect 15381 12795 15439 12801
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12636 12736 13093 12764
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 13538 12696 13544 12708
rect 12943 12668 13544 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 13538 12656 13544 12668
rect 13596 12656 13602 12708
rect 15488 12705 15516 12804
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17236 12832 17264 12860
rect 17092 12804 17264 12832
rect 17092 12792 17098 12804
rect 17696 12773 17724 12872
rect 18570 12869 18582 12872
rect 18616 12900 18628 12903
rect 18966 12900 18972 12912
rect 18616 12872 18972 12900
rect 18616 12869 18628 12872
rect 18570 12863 18628 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 20165 12903 20223 12909
rect 20165 12869 20177 12903
rect 20211 12900 20223 12903
rect 20530 12900 20536 12912
rect 20211 12872 20536 12900
rect 20211 12869 20223 12872
rect 20165 12863 20223 12869
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 20717 12903 20775 12909
rect 20717 12869 20729 12903
rect 20763 12900 20775 12903
rect 21266 12900 21272 12912
rect 20763 12872 21272 12900
rect 20763 12869 20775 12872
rect 20717 12863 20775 12869
rect 21266 12860 21272 12872
rect 21324 12860 21330 12912
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18230 12832 18236 12844
rect 17911 12804 18236 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 20438 12832 20444 12844
rect 20399 12804 20444 12832
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 17681 12767 17739 12773
rect 17681 12733 17693 12767
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 18046 12764 18052 12776
rect 17819 12736 18052 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 15473 12699 15531 12705
rect 15473 12665 15485 12699
rect 15519 12696 15531 12699
rect 16117 12699 16175 12705
rect 16117 12696 16129 12699
rect 15519 12668 16129 12696
rect 15519 12665 15531 12668
rect 15473 12659 15531 12665
rect 16117 12665 16129 12668
rect 16163 12696 16175 12699
rect 16206 12696 16212 12708
rect 16163 12668 16212 12696
rect 16163 12665 16175 12668
rect 16117 12659 16175 12665
rect 16206 12656 16212 12668
rect 16264 12696 16270 12708
rect 16393 12699 16451 12705
rect 16393 12696 16405 12699
rect 16264 12668 16405 12696
rect 16264 12656 16270 12668
rect 16393 12665 16405 12668
rect 16439 12696 16451 12699
rect 18340 12696 18368 12727
rect 16439 12668 18368 12696
rect 16439 12665 16451 12668
rect 16393 12659 16451 12665
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12628 11023 12631
rect 12986 12628 12992 12640
rect 11011 12600 12992 12628
rect 11011 12597 11023 12600
rect 10965 12591 11023 12597
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 13725 12631 13783 12637
rect 13725 12628 13737 12631
rect 13504 12600 13737 12628
rect 13504 12588 13510 12600
rect 13725 12597 13737 12600
rect 13771 12597 13783 12631
rect 13725 12591 13783 12597
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 15194 12628 15200 12640
rect 14047 12600 15200 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 15620 12600 15669 12628
rect 15620 12588 15626 12600
rect 15657 12597 15669 12600
rect 15703 12597 15715 12631
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 15657 12591 15715 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 17276 12600 17325 12628
rect 17276 12588 17282 12600
rect 17313 12597 17325 12600
rect 17359 12628 17371 12631
rect 17586 12628 17592 12640
rect 17359 12600 17592 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18322 12628 18328 12640
rect 18012 12600 18328 12628
rect 18012 12588 18018 12600
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19058 12628 19064 12640
rect 18748 12600 19064 12628
rect 18748 12588 18754 12600
rect 19058 12588 19064 12600
rect 19116 12628 19122 12640
rect 20257 12631 20315 12637
rect 20257 12628 20269 12631
rect 19116 12600 20269 12628
rect 19116 12588 19122 12600
rect 20257 12597 20269 12600
rect 20303 12597 20315 12631
rect 20257 12591 20315 12597
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20956 12600 21097 12628
rect 20956 12588 20962 12600
rect 21085 12597 21097 12600
rect 21131 12628 21143 12631
rect 22370 12628 22376 12640
rect 21131 12600 22376 12628
rect 21131 12597 21143 12600
rect 21085 12591 21143 12597
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1912 12396 1961 12424
rect 1912 12384 1918 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 2406 12424 2412 12436
rect 2367 12396 2412 12424
rect 1949 12387 2007 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3200 12396 3801 12424
rect 3200 12384 3206 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 4798 12424 4804 12436
rect 3789 12387 3847 12393
rect 3896 12396 4804 12424
rect 3896 12368 3924 12396
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 6052 12396 6285 12424
rect 6052 12384 6058 12396
rect 6273 12393 6285 12396
rect 6319 12393 6331 12427
rect 7282 12424 7288 12436
rect 7243 12396 7288 12424
rect 6273 12387 6331 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 7708 12396 8217 12424
rect 7708 12384 7714 12396
rect 8205 12393 8217 12396
rect 8251 12424 8263 12427
rect 8251 12396 12296 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2556 12328 3832 12356
rect 2556 12316 2562 12328
rect 2516 12288 2544 12316
rect 2148 12260 2544 12288
rect 3053 12291 3111 12297
rect 2148 12229 2176 12260
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3326 12288 3332 12300
rect 3099 12260 3332 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 1780 12152 1808 12183
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 3234 12220 3240 12232
rect 2280 12192 2325 12220
rect 3195 12192 3240 12220
rect 2280 12180 2286 12192
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 3804 12220 3832 12328
rect 3878 12316 3884 12368
rect 3936 12316 3942 12368
rect 3970 12316 3976 12368
rect 4028 12356 4034 12368
rect 6181 12359 6239 12365
rect 4028 12328 4384 12356
rect 4028 12316 4034 12328
rect 4246 12288 4252 12300
rect 4207 12260 4252 12288
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4356 12297 4384 12328
rect 6181 12325 6193 12359
rect 6227 12356 6239 12359
rect 6638 12356 6644 12368
rect 6227 12328 6644 12356
rect 6227 12325 6239 12328
rect 6181 12319 6239 12325
rect 6638 12316 6644 12328
rect 6696 12356 6702 12368
rect 7300 12356 7328 12384
rect 7837 12359 7895 12365
rect 7837 12356 7849 12359
rect 6696 12328 6868 12356
rect 7300 12328 7849 12356
rect 6696 12316 6702 12328
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 4522 12248 4528 12300
rect 4580 12288 4586 12300
rect 6840 12297 6868 12328
rect 7837 12325 7849 12328
rect 7883 12356 7895 12359
rect 9950 12356 9956 12368
rect 7883 12328 9956 12356
rect 7883 12325 7895 12328
rect 7837 12319 7895 12325
rect 8220 12300 8248 12328
rect 9950 12316 9956 12328
rect 10008 12316 10014 12368
rect 12268 12356 12296 12396
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 12400 12396 12449 12424
rect 12400 12384 12406 12396
rect 12437 12393 12449 12396
rect 12483 12393 12495 12427
rect 12437 12387 12495 12393
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 14553 12427 14611 12433
rect 14553 12424 14565 12427
rect 13044 12396 14565 12424
rect 13044 12384 13050 12396
rect 14553 12393 14565 12396
rect 14599 12424 14611 12427
rect 15473 12427 15531 12433
rect 14599 12396 15415 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 15286 12356 15292 12368
rect 12268 12328 15292 12356
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 15387 12356 15415 12396
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15519 12396 16252 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15746 12356 15752 12368
rect 15387 12328 15752 12356
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 16224 12356 16252 12396
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16356 12396 16405 12424
rect 16356 12384 16362 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 18046 12424 18052 12436
rect 18007 12396 18052 12424
rect 16393 12387 16451 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 19337 12427 19395 12433
rect 19337 12393 19349 12427
rect 19383 12424 19395 12427
rect 19702 12424 19708 12436
rect 19383 12396 19708 12424
rect 19383 12393 19395 12396
rect 19337 12387 19395 12393
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 20622 12384 20628 12436
rect 20680 12424 20686 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20680 12396 21005 12424
rect 20680 12384 20686 12396
rect 20993 12393 21005 12396
rect 21039 12393 21051 12427
rect 20993 12387 21051 12393
rect 20438 12356 20444 12368
rect 16224 12328 20444 12356
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 4801 12291 4859 12297
rect 4801 12288 4813 12291
rect 4580 12260 4813 12288
rect 4580 12248 4586 12260
rect 4801 12257 4813 12260
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 6825 12251 6883 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 8665 12291 8723 12297
rect 8665 12288 8677 12291
rect 8352 12260 8677 12288
rect 8352 12248 8358 12260
rect 8665 12257 8677 12260
rect 8711 12257 8723 12291
rect 13170 12288 13176 12300
rect 13131 12260 13176 12288
rect 8665 12251 8723 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13780 12260 13829 12288
rect 13780 12248 13786 12260
rect 13817 12257 13829 12260
rect 13863 12288 13875 12291
rect 14182 12288 14188 12300
rect 13863 12260 14188 12288
rect 13863 12257 13875 12260
rect 13817 12251 13875 12257
rect 14182 12248 14188 12260
rect 14240 12288 14246 12300
rect 14642 12288 14648 12300
rect 14240 12260 14648 12288
rect 14240 12248 14246 12260
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15194 12288 15200 12300
rect 14967 12260 15200 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12257 16267 12291
rect 16942 12288 16948 12300
rect 16903 12260 16948 12288
rect 16209 12251 16267 12257
rect 3804 12192 4292 12220
rect 3326 12152 3332 12164
rect 1780 12124 3332 12152
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3620 12124 4169 12152
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 3620 12093 3648 12124
rect 4157 12121 4169 12124
rect 4203 12121 4215 12155
rect 4157 12115 4215 12121
rect 4264 12096 4292 12192
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 7282 12220 7288 12232
rect 6604 12192 7288 12220
rect 6604 12180 6610 12192
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 11146 12220 11152 12232
rect 11103 12192 11152 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14550 12220 14556 12232
rect 14415 12192 14556 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 5068 12155 5126 12161
rect 5068 12121 5080 12155
rect 5114 12152 5126 12155
rect 5534 12152 5540 12164
rect 5114 12124 5540 12152
rect 5114 12121 5126 12124
rect 5068 12115 5126 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6972 12124 7205 12152
rect 6972 12112 6978 12124
rect 7193 12121 7205 12124
rect 7239 12152 7251 12155
rect 7742 12152 7748 12164
rect 7239 12124 7748 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 11302 12155 11360 12161
rect 11302 12152 11314 12155
rect 11072 12124 11314 12152
rect 11072 12096 11100 12124
rect 11302 12121 11314 12124
rect 11348 12121 11360 12155
rect 11302 12115 11360 12121
rect 12158 12112 12164 12164
rect 12216 12152 12222 12164
rect 13449 12155 13507 12161
rect 13449 12152 13461 12155
rect 12216 12124 13461 12152
rect 12216 12112 12222 12124
rect 13449 12121 13461 12124
rect 13495 12121 13507 12155
rect 14384 12152 14412 12183
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 16224 12220 16252 12251
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 18138 12288 18144 12300
rect 17451 12260 18144 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 18782 12288 18788 12300
rect 18739 12260 18788 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 19978 12248 19984 12300
rect 20036 12288 20042 12300
rect 20714 12288 20720 12300
rect 20036 12260 20720 12288
rect 20036 12248 20042 12260
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 15804 12192 16252 12220
rect 15804 12180 15810 12192
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 16724 12192 17601 12220
rect 16724 12180 16730 12192
rect 17589 12189 17601 12192
rect 17635 12220 17647 12223
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 17635 12192 18889 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 18877 12189 18889 12192
rect 18923 12189 18935 12223
rect 20162 12220 20168 12232
rect 20123 12192 20168 12220
rect 18877 12183 18935 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 20809 12223 20867 12229
rect 20809 12220 20821 12223
rect 20487 12192 20821 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 20809 12189 20821 12192
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 13449 12115 13507 12121
rect 13648 12124 14412 12152
rect 15105 12155 15163 12161
rect 2777 12087 2835 12093
rect 2777 12084 2789 12087
rect 2464 12056 2789 12084
rect 2464 12044 2470 12056
rect 2777 12053 2789 12056
rect 2823 12084 2835 12087
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 2823 12056 3157 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4614 12084 4620 12096
rect 4304 12056 4620 12084
rect 4304 12044 4310 12056
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6788 12056 6833 12084
rect 6788 12044 6794 12056
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 9398 12084 9404 12096
rect 7064 12056 9404 12084
rect 7064 12044 7070 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9582 12084 9588 12096
rect 9543 12056 9588 12084
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 11054 12044 11060 12096
rect 11112 12044 11118 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 12250 12084 12256 12096
rect 11204 12056 12256 12084
rect 11204 12044 11210 12056
rect 12250 12044 12256 12056
rect 12308 12044 12314 12096
rect 12618 12084 12624 12096
rect 12579 12056 12624 12084
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13081 12087 13139 12093
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13648 12084 13676 12124
rect 15105 12121 15117 12155
rect 15151 12152 15163 12155
rect 16758 12152 16764 12164
rect 15151 12124 15608 12152
rect 16719 12124 16764 12152
rect 15151 12121 15163 12124
rect 15105 12115 15163 12121
rect 13127 12056 13676 12084
rect 15013 12087 15071 12093
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 15013 12053 15025 12087
rect 15059 12084 15071 12087
rect 15286 12084 15292 12096
rect 15059 12056 15292 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15580 12093 15608 12124
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 17218 12112 17224 12164
rect 17276 12152 17282 12164
rect 17497 12155 17555 12161
rect 17497 12152 17509 12155
rect 17276 12124 17509 12152
rect 17276 12112 17282 12124
rect 17497 12121 17509 12124
rect 17543 12121 17555 12155
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 17497 12115 17555 12121
rect 17972 12124 18521 12152
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12053 15623 12087
rect 15930 12084 15936 12096
rect 15891 12056 15936 12084
rect 15565 12047 15623 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16022 12044 16028 12096
rect 16080 12084 16086 12096
rect 16853 12087 16911 12093
rect 16080 12056 16125 12084
rect 16080 12044 16086 12056
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 17770 12084 17776 12096
rect 16899 12056 17776 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17972 12093 18000 12124
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 18417 12087 18475 12093
rect 18417 12053 18429 12087
rect 18463 12084 18475 12087
rect 18598 12084 18604 12096
rect 18463 12056 18604 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19429 12087 19487 12093
rect 19429 12084 19441 12087
rect 19116 12056 19441 12084
rect 19116 12044 19122 12056
rect 19429 12053 19441 12056
rect 19475 12053 19487 12087
rect 19429 12047 19487 12053
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 21453 12087 21511 12093
rect 21453 12084 21465 12087
rect 21416 12056 21465 12084
rect 21416 12044 21422 12056
rect 21453 12053 21465 12056
rect 21499 12053 21511 12087
rect 21453 12047 21511 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2222 11880 2228 11892
rect 1964 11852 2228 11880
rect 1964 11821 1992 11852
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 4706 11880 4712 11892
rect 2746 11852 4712 11880
rect 1949 11815 2007 11821
rect 1949 11781 1961 11815
rect 1995 11781 2007 11815
rect 1949 11775 2007 11781
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 2746 11812 2774 11852
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 4856 11852 5089 11880
rect 4856 11840 4862 11852
rect 5077 11849 5089 11852
rect 5123 11880 5135 11883
rect 5442 11880 5448 11892
rect 5123 11852 5448 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5767 11852 6469 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 6963 11852 7297 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7650 11880 7656 11892
rect 7611 11852 7656 11880
rect 7285 11843 7343 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11849 8171 11883
rect 8113 11843 8171 11849
rect 8481 11883 8539 11889
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 8662 11880 8668 11892
rect 8527 11852 8668 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 2556 11784 2774 11812
rect 2556 11772 2562 11784
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 3973 11815 4031 11821
rect 3973 11812 3985 11815
rect 3292 11784 3985 11812
rect 3292 11772 3298 11784
rect 3973 11781 3985 11784
rect 4019 11812 4031 11815
rect 4062 11812 4068 11824
rect 4019 11784 4068 11812
rect 4019 11781 4031 11784
rect 3973 11775 4031 11781
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 4246 11812 4252 11824
rect 4203 11784 4252 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 4246 11772 4252 11784
rect 4304 11812 4310 11824
rect 4522 11812 4528 11824
rect 4304 11784 4528 11812
rect 4304 11772 4310 11784
rect 4522 11772 4528 11784
rect 4580 11772 4586 11824
rect 4890 11812 4896 11824
rect 4851 11784 4896 11812
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 6825 11815 6883 11821
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 8128 11812 8156 11843
rect 8662 11840 8668 11852
rect 8720 11880 8726 11892
rect 11238 11880 11244 11892
rect 8720 11852 11244 11880
rect 8720 11840 8726 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11480 11852 11805 11880
rect 11480 11840 11486 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 12158 11880 12164 11892
rect 11793 11843 11851 11849
rect 11992 11852 12164 11880
rect 6871 11784 8156 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 8294 11772 8300 11824
rect 8352 11812 8358 11824
rect 11885 11815 11943 11821
rect 8352 11784 10732 11812
rect 8352 11772 8358 11784
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2682 11744 2688 11756
rect 2271 11716 2360 11744
rect 2643 11716 2688 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 2332 11617 2360 11716
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4982 11744 4988 11756
rect 4764 11716 4988 11744
rect 4764 11704 4770 11716
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9493 11747 9551 11753
rect 8628 11716 9076 11744
rect 8628 11704 8634 11716
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2958 11676 2964 11688
rect 2832 11648 2877 11676
rect 2919 11648 2964 11676
rect 2832 11636 2838 11648
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 5534 11676 5540 11688
rect 5495 11648 5540 11676
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6604 11648 7021 11676
rect 6604 11636 6610 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7742 11676 7748 11688
rect 7703 11648 7748 11676
rect 7009 11639 7067 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11577 2375 11611
rect 2317 11571 2375 11577
rect 3970 11568 3976 11620
rect 4028 11608 4034 11620
rect 6181 11611 6239 11617
rect 4028 11580 5304 11608
rect 4028 11568 4034 11580
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 5132 11512 5181 11540
rect 5132 11500 5138 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5276 11540 5304 11580
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 6730 11608 6736 11620
rect 6227 11580 6736 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7944 11608 7972 11639
rect 8680 11608 8708 11639
rect 6972 11580 8708 11608
rect 6972 11568 6978 11580
rect 7926 11540 7932 11552
rect 5276 11512 7932 11540
rect 5169 11503 5227 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 9048 11549 9076 11716
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9766 11744 9772 11756
rect 9539 11716 9772 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 10220 11747 10278 11753
rect 10220 11713 10232 11747
rect 10266 11744 10278 11747
rect 10502 11744 10508 11756
rect 10266 11716 10508 11744
rect 10266 11713 10278 11716
rect 10220 11707 10278 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10704 11744 10732 11784
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 11992 11812 12020 11852
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 12299 11852 13553 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 14792 11852 15577 11880
rect 14792 11840 14798 11852
rect 15565 11849 15577 11852
rect 15611 11880 15623 11883
rect 15746 11880 15752 11892
rect 15611 11852 15752 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16080 11852 16681 11880
rect 16080 11840 16086 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 16669 11843 16727 11849
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 18693 11883 18751 11889
rect 18693 11880 18705 11883
rect 17828 11852 18705 11880
rect 17828 11840 17834 11852
rect 18693 11849 18705 11852
rect 18739 11880 18751 11883
rect 18966 11880 18972 11892
rect 18739 11852 18972 11880
rect 18739 11849 18751 11852
rect 18693 11843 18751 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 12802 11812 12808 11824
rect 11931 11784 12020 11812
rect 12763 11784 12808 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13446 11772 13452 11824
rect 13504 11812 13510 11824
rect 13633 11815 13691 11821
rect 13633 11812 13645 11815
rect 13504 11784 13645 11812
rect 13504 11772 13510 11784
rect 13633 11781 13645 11784
rect 13679 11781 13691 11815
rect 13633 11775 13691 11781
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 16117 11815 16175 11821
rect 16117 11812 16129 11815
rect 13872 11784 16129 11812
rect 13872 11772 13878 11784
rect 16117 11781 16129 11784
rect 16163 11781 16175 11815
rect 16117 11775 16175 11781
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 17865 11815 17923 11821
rect 17865 11812 17877 11815
rect 17552 11784 17877 11812
rect 17552 11772 17558 11784
rect 17865 11781 17877 11784
rect 17911 11812 17923 11815
rect 17954 11812 17960 11824
rect 17911 11784 17960 11812
rect 17911 11781 17923 11784
rect 17865 11775 17923 11781
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 18064 11784 18613 11812
rect 11514 11744 11520 11756
rect 10704 11716 11520 11744
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 12250 11744 12256 11756
rect 11624 11716 12256 11744
rect 9214 11676 9220 11688
rect 9175 11648 9220 11676
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9398 11676 9404 11688
rect 9359 11648 9404 11676
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 11624 11685 11652 11716
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12584 11716 12725 11744
rect 12584 11704 12590 11716
rect 12713 11713 12725 11716
rect 12759 11744 12771 11747
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 12759 11716 14013 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14182 11744 14188 11756
rect 14143 11716 14188 11744
rect 14001 11707 14059 11713
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11676 13047 11679
rect 13170 11676 13176 11688
rect 13035 11648 13176 11676
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11330 11608 11336 11620
rect 11112 11580 11336 11608
rect 11112 11568 11118 11580
rect 11330 11568 11336 11580
rect 11388 11608 11394 11620
rect 13004 11608 13032 11639
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13504 11648 13737 11676
rect 13504 11636 13510 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 11388 11580 13032 11608
rect 11388 11568 11394 11580
rect 9033 11543 9091 11549
rect 9033 11509 9045 11543
rect 9079 11540 9091 11543
rect 9306 11540 9312 11552
rect 9079 11512 9312 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 12342 11540 12348 11552
rect 12303 11512 12348 11540
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 13170 11540 13176 11552
rect 13131 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 14016 11540 14044 11707
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14458 11753 14464 11756
rect 14452 11744 14464 11753
rect 14371 11716 14464 11744
rect 14452 11707 14464 11716
rect 14516 11744 14522 11756
rect 14516 11716 15516 11744
rect 14458 11704 14464 11707
rect 14516 11704 14522 11716
rect 15488 11676 15516 11716
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16025 11747 16083 11753
rect 16025 11744 16037 11747
rect 15620 11716 16037 11744
rect 15620 11704 15626 11716
rect 16025 11713 16037 11716
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16206 11704 16212 11756
rect 16264 11744 16270 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16264 11716 17049 11744
rect 16264 11704 16270 11716
rect 17037 11713 17049 11716
rect 17083 11744 17095 11747
rect 18064 11744 18092 11784
rect 18601 11781 18613 11784
rect 18647 11812 18659 11815
rect 21174 11812 21180 11824
rect 18647 11784 21180 11812
rect 18647 11781 18659 11784
rect 18601 11775 18659 11781
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 19058 11744 19064 11756
rect 17083 11716 18092 11744
rect 19019 11716 19064 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 19328 11747 19386 11753
rect 19328 11713 19340 11747
rect 19374 11744 19386 11747
rect 19610 11744 19616 11756
rect 19374 11716 19616 11744
rect 19374 11713 19386 11716
rect 19328 11707 19386 11713
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20180 11716 21005 11744
rect 16298 11676 16304 11688
rect 15488 11648 15700 11676
rect 16259 11648 16304 11676
rect 15672 11608 15700 11648
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 17126 11676 17132 11688
rect 17087 11648 17132 11676
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 17221 11679 17279 11685
rect 17221 11645 17233 11679
rect 17267 11645 17279 11679
rect 17221 11639 17279 11645
rect 17589 11679 17647 11685
rect 17589 11645 17601 11679
rect 17635 11645 17647 11679
rect 17770 11676 17776 11688
rect 17731 11648 17776 11676
rect 17589 11639 17647 11645
rect 16850 11608 16856 11620
rect 15672 11580 16856 11608
rect 16850 11568 16856 11580
rect 16908 11608 16914 11620
rect 17236 11608 17264 11639
rect 16908 11580 17264 11608
rect 17604 11608 17632 11639
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 19076 11676 19104 11704
rect 18463 11648 19104 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 17862 11608 17868 11620
rect 17604 11580 17868 11608
rect 16908 11568 16914 11580
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 18012 11580 18889 11608
rect 18012 11568 18018 11580
rect 18877 11577 18889 11580
rect 18923 11577 18935 11611
rect 18877 11571 18935 11577
rect 15562 11540 15568 11552
rect 14016 11512 15568 11540
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 15657 11543 15715 11549
rect 15657 11509 15669 11543
rect 15703 11540 15715 11543
rect 15838 11540 15844 11552
rect 15703 11512 15844 11540
rect 15703 11509 15715 11512
rect 15657 11503 15715 11509
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 18046 11540 18052 11552
rect 17368 11512 18052 11540
rect 17368 11500 17374 11512
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18230 11540 18236 11552
rect 18191 11512 18236 11540
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 20180 11540 20208 11716
rect 20993 11713 21005 11716
rect 21039 11744 21051 11747
rect 21358 11744 21364 11756
rect 21039 11716 21364 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 21358 11704 21364 11716
rect 21416 11744 21422 11756
rect 22094 11744 22100 11756
rect 21416 11716 22100 11744
rect 21416 11704 21422 11716
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21634 11676 21640 11688
rect 20947 11648 21640 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 20824 11608 20852 11639
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 21174 11608 21180 11620
rect 20824 11580 21180 11608
rect 21174 11568 21180 11580
rect 21232 11568 21238 11620
rect 21266 11568 21272 11620
rect 21324 11608 21330 11620
rect 21453 11611 21511 11617
rect 21453 11608 21465 11611
rect 21324 11580 21465 11608
rect 21324 11568 21330 11580
rect 21453 11577 21465 11580
rect 21499 11577 21511 11611
rect 21453 11571 21511 11577
rect 20438 11540 20444 11552
rect 19024 11512 20208 11540
rect 20399 11512 20444 11540
rect 19024 11500 19030 11512
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3053 11339 3111 11345
rect 3053 11336 3065 11339
rect 3016 11308 3065 11336
rect 3016 11296 3022 11308
rect 3053 11305 3065 11308
rect 3099 11305 3111 11339
rect 3053 11299 3111 11305
rect 3237 11339 3295 11345
rect 3237 11305 3249 11339
rect 3283 11336 3295 11339
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3283 11308 3433 11336
rect 3283 11305 3295 11308
rect 3237 11299 3295 11305
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 3510 11336 3516 11348
rect 3467 11308 3516 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3510 11296 3516 11308
rect 3568 11336 3574 11348
rect 4246 11336 4252 11348
rect 3568 11308 4252 11336
rect 3568 11296 3574 11308
rect 4246 11296 4252 11308
rect 4304 11336 4310 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 4304 11308 4353 11336
rect 4304 11296 4310 11308
rect 4341 11305 4353 11308
rect 4387 11305 4399 11339
rect 5258 11336 5264 11348
rect 4341 11299 4399 11305
rect 4632 11308 5264 11336
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 4632 11268 4660 11308
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 5868 11308 6745 11336
rect 5868 11296 5874 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8757 11339 8815 11345
rect 8260 11296 8294 11336
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 9398 11336 9404 11348
rect 8803 11308 9404 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10965 11339 11023 11345
rect 10965 11305 10977 11339
rect 11011 11336 11023 11339
rect 11422 11336 11428 11348
rect 11011 11308 11428 11336
rect 11011 11305 11023 11308
rect 10965 11299 11023 11305
rect 2924 11240 4660 11268
rect 5552 11268 5580 11296
rect 5997 11271 6055 11277
rect 5997 11268 6009 11271
rect 5552 11240 6009 11268
rect 2924 11228 2930 11240
rect 5997 11237 6009 11240
rect 6043 11237 6055 11271
rect 8266 11268 8294 11296
rect 8266 11240 9168 11268
rect 5997 11231 6055 11237
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 3936 11172 4752 11200
rect 3936 11160 3942 11172
rect 1486 11092 1492 11144
rect 1544 11132 1550 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1544 11104 1685 11132
rect 1544 11092 1550 11104
rect 1673 11101 1685 11104
rect 1719 11132 1731 11135
rect 3510 11132 3516 11144
rect 1719 11104 3516 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 1940 11067 1998 11073
rect 1940 11033 1952 11067
rect 1986 11064 1998 11067
rect 2590 11064 2596 11076
rect 1986 11036 2596 11064
rect 1986 11033 1998 11036
rect 1940 11027 1998 11033
rect 2590 11024 2596 11036
rect 2648 11024 2654 11076
rect 4448 10996 4476 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4724 11132 4752 11172
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6604 11172 7297 11200
rect 6604 11160 6610 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 8570 11200 8576 11212
rect 8251 11172 8576 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9140 11209 9168 11240
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 4724 11104 8524 11132
rect 4617 11095 4675 11101
rect 4522 11024 4528 11076
rect 4580 11064 4586 11076
rect 4862 11067 4920 11073
rect 4862 11064 4874 11067
rect 4580 11036 4874 11064
rect 4580 11024 4586 11036
rect 4862 11033 4874 11036
rect 4908 11033 4920 11067
rect 4862 11027 4920 11033
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5316 11036 7420 11064
rect 5316 11024 5322 11036
rect 5994 10996 6000 11008
rect 4448 10968 6000 10996
rect 5994 10956 6000 10968
rect 6052 10996 6058 11008
rect 6089 10999 6147 11005
rect 6089 10996 6101 10999
rect 6052 10968 6101 10996
rect 6052 10956 6058 10968
rect 6089 10965 6101 10968
rect 6135 10965 6147 10999
rect 6089 10959 6147 10965
rect 6641 10999 6699 11005
rect 6641 10965 6653 10999
rect 6687 10996 6699 10999
rect 7006 10996 7012 11008
rect 6687 10968 7012 10996
rect 6687 10965 6699 10968
rect 6641 10959 6699 10965
rect 7006 10956 7012 10968
rect 7064 10996 7070 11008
rect 7101 10999 7159 11005
rect 7101 10996 7113 10999
rect 7064 10968 7113 10996
rect 7064 10956 7070 10968
rect 7101 10965 7113 10968
rect 7147 10965 7159 10999
rect 7101 10959 7159 10965
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7392 10996 7420 11036
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7524 11036 7849 11064
rect 7524 11024 7530 11036
rect 7837 11033 7849 11036
rect 7883 11064 7895 11067
rect 8018 11064 8024 11076
rect 7883 11036 8024 11064
rect 7883 11033 7895 11036
rect 7837 11027 7895 11033
rect 8018 11024 8024 11036
rect 8076 11064 8082 11076
rect 8389 11067 8447 11073
rect 8389 11064 8401 11067
rect 8076 11036 8401 11064
rect 8076 11024 8082 11036
rect 8389 11033 8401 11036
rect 8435 11033 8447 11067
rect 8496 11064 8524 11104
rect 8662 11092 8668 11144
rect 8720 11132 8726 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8720 11104 8953 11132
rect 8720 11092 8726 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9381 11135 9439 11141
rect 9381 11132 9393 11135
rect 9272 11104 9393 11132
rect 9272 11092 9278 11104
rect 9381 11101 9393 11104
rect 9427 11101 9439 11135
rect 10980 11132 11008 11299
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13872 11308 14381 11336
rect 13872 11296 13878 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 14369 11299 14427 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 17770 11336 17776 11348
rect 16356 11308 17356 11336
rect 17731 11308 17776 11336
rect 16356 11296 16362 11308
rect 17328 11280 17356 11308
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 18598 11336 18604 11348
rect 18559 11308 18604 11336
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 19886 11336 19892 11348
rect 19383 11308 19892 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 12250 11268 12256 11280
rect 12176 11240 12256 11268
rect 11330 11200 11336 11212
rect 11291 11172 11336 11200
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 12176 11209 12204 11240
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12805 11271 12863 11277
rect 12805 11237 12817 11271
rect 12851 11268 12863 11271
rect 15381 11271 15439 11277
rect 15381 11268 15393 11271
rect 12851 11240 13400 11268
rect 12851 11237 12863 11240
rect 12805 11231 12863 11237
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11940 11172 12173 11200
rect 11940 11160 11946 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12342 11200 12348 11212
rect 12303 11172 12348 11200
rect 12161 11163 12219 11169
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 13372 11209 13400 11240
rect 14844 11240 15393 11268
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 13814 11200 13820 11212
rect 13504 11172 13549 11200
rect 13775 11172 13820 11200
rect 13504 11160 13510 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 14844 11209 14872 11240
rect 15381 11237 15393 11240
rect 15427 11237 15439 11271
rect 15381 11231 15439 11237
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 15620 11240 17172 11268
rect 15620 11228 15626 11240
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11169 14887 11203
rect 15838 11200 15844 11212
rect 15799 11172 15844 11200
rect 14829 11163 14887 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16025 11203 16083 11209
rect 16025 11169 16037 11203
rect 16071 11200 16083 11203
rect 16850 11200 16856 11212
rect 16071 11172 16856 11200
rect 16071 11169 16083 11172
rect 16025 11163 16083 11169
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 9381 11095 9439 11101
rect 9508 11104 11008 11132
rect 9508 11064 9536 11104
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11112 11104 11529 11132
rect 11112 11092 11118 11104
rect 11517 11101 11529 11104
rect 11563 11132 11575 11135
rect 12437 11135 12495 11141
rect 11563 11104 12388 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 8496 11036 9536 11064
rect 8389 11027 8447 11033
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10778 11064 10784 11076
rect 10008 11036 10784 11064
rect 10008 11024 10014 11036
rect 10778 11024 10784 11036
rect 10836 11064 10842 11076
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 10836 11036 11161 11064
rect 10836 11024 10842 11036
rect 11149 11033 11161 11036
rect 11195 11064 11207 11067
rect 12250 11064 12256 11076
rect 11195 11036 12256 11064
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12360 11064 12388 11104
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12618 11132 12624 11144
rect 12483 11104 12624 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 13832 11064 13860 11160
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16172 11104 16681 11132
rect 16172 11092 16178 11104
rect 16669 11101 16681 11104
rect 16715 11132 16727 11135
rect 17034 11132 17040 11144
rect 16715 11104 17040 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 17144 11132 17172 11240
rect 17310 11228 17316 11280
rect 17368 11268 17374 11280
rect 19429 11271 19487 11277
rect 19429 11268 19441 11271
rect 17368 11240 19441 11268
rect 17368 11228 17374 11240
rect 19429 11237 19441 11240
rect 19475 11237 19487 11271
rect 19429 11231 19487 11237
rect 17221 11203 17279 11209
rect 17221 11169 17233 11203
rect 17267 11200 17279 11203
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17267 11172 18061 11200
rect 17267 11169 17279 11172
rect 17221 11163 17279 11169
rect 18049 11169 18061 11172
rect 18095 11200 18107 11203
rect 18138 11200 18144 11212
rect 18095 11172 18144 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 17954 11132 17960 11144
rect 17144 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11132 18291 11135
rect 19536 11132 19564 11308
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20530 11296 20536 11348
rect 20588 11336 20594 11348
rect 21085 11339 21143 11345
rect 21085 11336 21097 11339
rect 20588 11308 21097 11336
rect 20588 11296 20594 11308
rect 21085 11305 21097 11308
rect 21131 11305 21143 11339
rect 21085 11299 21143 11305
rect 20809 11203 20867 11209
rect 20809 11169 20821 11203
rect 20855 11200 20867 11203
rect 20855 11172 20889 11200
rect 20855 11169 20867 11172
rect 20809 11163 20867 11169
rect 20824 11132 20852 11163
rect 18279 11104 19564 11132
rect 19628 11104 20852 11132
rect 18279 11101 18291 11104
rect 18233 11095 18291 11101
rect 12360 11036 13860 11064
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 15102 11064 15108 11076
rect 14608 11036 15108 11064
rect 14608 11024 14614 11036
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15749 11067 15807 11073
rect 15749 11033 15761 11067
rect 15795 11064 15807 11067
rect 16942 11064 16948 11076
rect 15795 11036 16948 11064
rect 15795 11033 15807 11036
rect 15749 11027 15807 11033
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 18877 11067 18935 11073
rect 18877 11064 18889 11067
rect 17359 11036 18889 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 18877 11033 18889 11036
rect 18923 11064 18935 11067
rect 19058 11064 19064 11076
rect 18923 11036 19064 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 19628 11064 19656 11104
rect 19208 11036 19656 11064
rect 19208 11024 19214 11036
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 20438 11064 20444 11076
rect 19760 11036 20444 11064
rect 19760 11024 19766 11036
rect 20438 11024 20444 11036
rect 20496 11064 20502 11076
rect 20542 11067 20600 11073
rect 20542 11064 20554 11067
rect 20496 11036 20554 11064
rect 20496 11024 20502 11036
rect 20542 11033 20554 11036
rect 20588 11033 20600 11067
rect 20824 11064 20852 11104
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11132 20959 11135
rect 21082 11132 21088 11144
rect 20947 11104 21088 11132
rect 20947 11101 20959 11104
rect 20901 11095 20959 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21266 11064 21272 11076
rect 20824 11036 21272 11064
rect 20542 11027 20600 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21545 11067 21603 11073
rect 21545 11033 21557 11067
rect 21591 11064 21603 11067
rect 21634 11064 21640 11076
rect 21591 11036 21640 11064
rect 21591 11033 21603 11036
rect 21545 11027 21603 11033
rect 21634 11024 21640 11036
rect 21692 11064 21698 11076
rect 22186 11064 22192 11076
rect 21692 11036 22192 11064
rect 21692 11024 21698 11036
rect 22186 11024 22192 11036
rect 22244 11024 22250 11076
rect 7653 10999 7711 11005
rect 7653 10996 7665 10999
rect 7248 10968 7293 10996
rect 7392 10968 7665 10996
rect 7248 10956 7254 10968
rect 7653 10965 7665 10968
rect 7699 10996 7711 10999
rect 8294 10996 8300 11008
rect 7699 10968 8300 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 10134 10956 10140 11008
rect 10192 10996 10198 11008
rect 10502 10996 10508 11008
rect 10192 10968 10508 10996
rect 10192 10956 10198 10968
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 11609 10999 11667 11005
rect 10652 10968 10697 10996
rect 10652 10956 10658 10968
rect 11609 10965 11621 10999
rect 11655 10996 11667 10999
rect 11698 10996 11704 11008
rect 11655 10968 11704 10996
rect 11655 10965 11667 10968
rect 11609 10959 11667 10965
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 11974 10996 11980 11008
rect 11935 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13262 10996 13268 11008
rect 12952 10968 12997 10996
rect 13223 10968 13268 10996
rect 12952 10956 12958 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 14918 10996 14924 11008
rect 14879 10968 14924 10996
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15378 10956 15384 11008
rect 15436 10996 15442 11008
rect 15838 10996 15844 11008
rect 15436 10968 15844 10996
rect 15436 10956 15442 10968
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 16209 10999 16267 11005
rect 16209 10996 16221 10999
rect 15988 10968 16221 10996
rect 15988 10956 15994 10968
rect 16209 10965 16221 10968
rect 16255 10965 16267 10999
rect 16209 10959 16267 10965
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16577 10999 16635 11005
rect 16577 10996 16589 10999
rect 16448 10968 16589 10996
rect 16448 10956 16454 10968
rect 16577 10965 16589 10968
rect 16623 10965 16635 10999
rect 16577 10959 16635 10965
rect 17405 10999 17463 11005
rect 17405 10965 17417 10999
rect 17451 10996 17463 10999
rect 17678 10996 17684 11008
rect 17451 10968 17684 10996
rect 17451 10965 17463 10968
rect 17405 10959 17463 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 18012 10968 18153 10996
rect 18012 10956 18018 10968
rect 18141 10965 18153 10968
rect 18187 10996 18199 10999
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 18187 10968 18705 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 18693 10965 18705 10968
rect 18739 10996 18751 10999
rect 18966 10996 18972 11008
rect 18739 10968 18972 10996
rect 18739 10965 18751 10968
rect 18693 10959 18751 10965
rect 18966 10956 18972 10968
rect 19024 10956 19030 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10761 4307 10795
rect 4249 10755 4307 10761
rect 2958 10684 2964 10736
rect 3016 10724 3022 10736
rect 3114 10727 3172 10733
rect 3114 10724 3126 10727
rect 3016 10696 3126 10724
rect 3016 10684 3022 10696
rect 3114 10693 3126 10696
rect 3160 10693 3172 10727
rect 3114 10687 3172 10693
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10656 1455 10659
rect 1486 10656 1492 10668
rect 1443 10628 1492 10656
rect 1443 10625 1455 10628
rect 1397 10619 1455 10625
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1670 10665 1676 10668
rect 1664 10619 1676 10665
rect 1728 10656 1734 10668
rect 2869 10659 2927 10665
rect 1728 10628 1764 10656
rect 1670 10616 1676 10619
rect 1728 10616 1734 10628
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3510 10656 3516 10668
rect 2915 10628 3516 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 4264 10656 4292 10755
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 5813 10795 5871 10801
rect 5813 10792 5825 10795
rect 4580 10764 5825 10792
rect 4580 10752 4586 10764
rect 5813 10761 5825 10764
rect 5859 10792 5871 10795
rect 6546 10792 6552 10804
rect 5859 10764 6552 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7248 10764 7481 10792
rect 7248 10752 7254 10764
rect 7469 10761 7481 10764
rect 7515 10761 7527 10795
rect 7469 10755 7527 10761
rect 8389 10795 8447 10801
rect 8389 10761 8401 10795
rect 8435 10792 8447 10795
rect 9214 10792 9220 10804
rect 8435 10764 9220 10792
rect 8435 10761 8447 10764
rect 8389 10755 8447 10761
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 5350 10724 5356 10736
rect 5132 10696 5356 10724
rect 5132 10684 5138 10696
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 6052 10696 6377 10724
rect 6052 10684 6058 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 6365 10687 6423 10693
rect 6454 10684 6460 10736
rect 6512 10724 6518 10736
rect 7101 10727 7159 10733
rect 7101 10724 7113 10727
rect 6512 10696 7113 10724
rect 6512 10684 6518 10696
rect 7101 10693 7113 10696
rect 7147 10724 7159 10727
rect 8404 10724 8432 10755
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9324 10764 9720 10792
rect 9324 10724 9352 10764
rect 7147 10696 7696 10724
rect 7147 10693 7159 10696
rect 7101 10687 7159 10693
rect 4700 10659 4758 10665
rect 4700 10656 4712 10659
rect 4264 10628 4712 10656
rect 4700 10625 4712 10628
rect 4746 10656 4758 10659
rect 4746 10628 6960 10656
rect 4746 10625 4758 10628
rect 4700 10619 4758 10625
rect 6932 10600 6960 10628
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4430 10588 4436 10600
rect 4304 10560 4436 10588
rect 4304 10548 4310 10560
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5902 10588 5908 10600
rect 5863 10560 5908 10588
rect 5902 10548 5908 10560
rect 5960 10548 5966 10600
rect 6454 10588 6460 10600
rect 6196 10560 6460 10588
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 6196 10520 6224 10560
rect 6454 10548 6460 10560
rect 6512 10588 6518 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6512 10560 6561 10588
rect 6512 10548 6518 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6914 10588 6920 10600
rect 6875 10560 6920 10588
rect 6549 10551 6607 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7064 10560 7109 10588
rect 7064 10548 7070 10560
rect 7466 10520 7472 10532
rect 5776 10492 6224 10520
rect 6288 10492 7472 10520
rect 5776 10480 5782 10492
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 2777 10455 2835 10461
rect 2777 10452 2789 10455
rect 2648 10424 2789 10452
rect 2648 10412 2654 10424
rect 2777 10421 2789 10424
rect 2823 10421 2835 10455
rect 2777 10415 2835 10421
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 6288 10452 6316 10492
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 7668 10520 7696 10696
rect 7852 10696 8432 10724
rect 8496 10696 9352 10724
rect 7852 10656 7880 10696
rect 7760 10628 7880 10656
rect 7929 10659 7987 10665
rect 7760 10597 7788 10628
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8294 10656 8300 10668
rect 7975 10628 8300 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8018 10588 8024 10600
rect 7883 10560 8024 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8496 10588 8524 10696
rect 9398 10684 9404 10736
rect 9456 10724 9462 10736
rect 9582 10724 9588 10736
rect 9456 10696 9588 10724
rect 9456 10684 9462 10696
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 9502 10659 9560 10665
rect 9502 10656 9514 10659
rect 8628 10628 9514 10656
rect 8628 10616 8634 10628
rect 9502 10625 9514 10628
rect 9548 10625 9560 10659
rect 9692 10656 9720 10764
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9824 10764 9873 10792
rect 9824 10752 9830 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10594 10792 10600 10804
rect 10275 10764 10600 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12802 10792 12808 10804
rect 12115 10764 12808 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13814 10792 13820 10804
rect 13775 10764 13820 10792
rect 13814 10752 13820 10764
rect 13872 10792 13878 10804
rect 14366 10792 14372 10804
rect 13872 10764 14372 10792
rect 13872 10752 13878 10764
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 14918 10792 14924 10804
rect 14691 10764 14924 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 16206 10792 16212 10804
rect 15028 10764 16212 10792
rect 10318 10724 10324 10736
rect 10279 10696 10324 10724
rect 10318 10684 10324 10696
rect 10376 10724 10382 10736
rect 10873 10727 10931 10733
rect 10873 10724 10885 10727
rect 10376 10696 10885 10724
rect 10376 10684 10382 10696
rect 10873 10693 10885 10696
rect 10919 10724 10931 10727
rect 11790 10724 11796 10736
rect 10919 10696 11796 10724
rect 10919 10693 10931 10696
rect 10873 10687 10931 10693
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 12520 10727 12578 10733
rect 12520 10693 12532 10727
rect 12566 10724 12578 10727
rect 13446 10724 13452 10736
rect 12566 10696 13452 10724
rect 12566 10693 12578 10696
rect 12520 10687 12578 10693
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 15028 10724 15056 10764
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 16390 10752 16396 10804
rect 16448 10792 16454 10804
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 16448 10764 16497 10792
rect 16448 10752 16454 10764
rect 16485 10761 16497 10764
rect 16531 10761 16543 10795
rect 16485 10755 16543 10761
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16724 10764 17141 10792
rect 16724 10752 16730 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 19610 10792 19616 10804
rect 19383 10764 19616 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 20220 10764 20269 10792
rect 20220 10752 20226 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 21266 10792 21272 10804
rect 21227 10764 21272 10792
rect 20257 10755 20315 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 13556 10696 15056 10724
rect 10962 10656 10968 10668
rect 9692 10628 10968 10656
rect 9502 10619 9560 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 12250 10656 12256 10668
rect 12211 10628 12256 10656
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 13556 10656 13584 10696
rect 15654 10684 15660 10736
rect 15712 10724 15718 10736
rect 15872 10727 15930 10733
rect 15872 10724 15884 10727
rect 15712 10696 15884 10724
rect 15712 10684 15718 10696
rect 15872 10693 15884 10696
rect 15918 10724 15930 10727
rect 17589 10727 17647 10733
rect 15918 10696 17264 10724
rect 15918 10693 15930 10696
rect 15872 10687 15930 10693
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 12360 10628 13584 10656
rect 13648 10628 14289 10656
rect 8220 10560 8524 10588
rect 9769 10591 9827 10597
rect 8220 10520 8248 10560
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 10505 10591 10563 10597
rect 9815 10560 10364 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 7668 10492 8248 10520
rect 8297 10523 8355 10529
rect 8297 10489 8309 10523
rect 8343 10520 8355 10523
rect 8343 10492 8892 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 4120 10424 6316 10452
rect 4120 10412 4126 10424
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8386 10452 8392 10464
rect 7708 10424 8392 10452
rect 7708 10412 7714 10424
rect 8386 10412 8392 10424
rect 8444 10452 8450 10464
rect 8662 10452 8668 10464
rect 8444 10424 8668 10452
rect 8444 10412 8450 10424
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8864 10452 8892 10492
rect 10336 10464 10364 10560
rect 10505 10557 10517 10591
rect 10551 10588 10563 10591
rect 10594 10588 10600 10600
rect 10551 10560 10600 10588
rect 10551 10557 10563 10560
rect 10505 10551 10563 10557
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 11330 10548 11336 10600
rect 11388 10588 11394 10600
rect 12360 10588 12388 10628
rect 11388 10560 12388 10588
rect 11388 10548 11394 10560
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13648 10588 13676 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 17034 10656 17040 10668
rect 16995 10628 17040 10656
rect 14277 10619 14335 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17236 10656 17264 10696
rect 17589 10693 17601 10727
rect 17635 10724 17647 10727
rect 19150 10724 19156 10736
rect 17635 10696 19156 10724
rect 17635 10693 17647 10696
rect 17589 10687 17647 10693
rect 17310 10656 17316 10668
rect 17236 10628 17316 10656
rect 13412 10560 13676 10588
rect 14093 10591 14151 10597
rect 13412 10548 13418 10560
rect 14093 10557 14105 10591
rect 14139 10557 14151 10591
rect 14093 10551 14151 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 15010 10588 15016 10600
rect 14231 10560 15016 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14108 10520 14136 10551
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 17236 10597 17264 10628
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17972 10597 18000 10696
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 19628 10724 19656 10752
rect 19628 10696 20852 10724
rect 18224 10659 18282 10665
rect 18224 10625 18236 10659
rect 18270 10656 18282 10659
rect 18598 10656 18604 10668
rect 18270 10628 18604 10656
rect 18270 10625 18282 10628
rect 18224 10619 18282 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 20070 10656 20076 10668
rect 19935 10628 20076 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20824 10656 20852 10696
rect 20824 10628 20944 10656
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 17221 10591 17279 10597
rect 16163 10560 17080 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 14458 10520 14464 10532
rect 14108 10492 14464 10520
rect 14458 10480 14464 10492
rect 14516 10520 14522 10532
rect 14737 10523 14795 10529
rect 14737 10520 14749 10523
rect 14516 10492 14749 10520
rect 14516 10480 14522 10492
rect 14737 10489 14749 10492
rect 14783 10489 14795 10523
rect 14737 10483 14795 10489
rect 16206 10480 16212 10532
rect 16264 10520 16270 10532
rect 16669 10523 16727 10529
rect 16264 10492 16528 10520
rect 16264 10480 16270 10492
rect 9582 10452 9588 10464
rect 8864 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 9950 10452 9956 10464
rect 9824 10424 9956 10452
rect 9824 10412 9830 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10778 10452 10784 10464
rect 10376 10424 10784 10452
rect 10376 10412 10382 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11149 10455 11207 10461
rect 11149 10421 11161 10455
rect 11195 10452 11207 10455
rect 11698 10452 11704 10464
rect 11195 10424 11704 10452
rect 11195 10421 11207 10424
rect 11149 10415 11207 10421
rect 11698 10412 11704 10424
rect 11756 10452 11762 10464
rect 12066 10452 12072 10464
rect 11756 10424 12072 10452
rect 11756 10412 11762 10424
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 13630 10452 13636 10464
rect 13591 10424 13636 10452
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 16500 10452 16528 10492
rect 16669 10489 16681 10523
rect 16715 10520 16727 10523
rect 16942 10520 16948 10532
rect 16715 10492 16948 10520
rect 16715 10489 16727 10492
rect 16669 10483 16727 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 17052 10520 17080 10560
rect 17221 10557 17233 10591
rect 17267 10557 17279 10591
rect 17957 10591 18015 10597
rect 17957 10588 17969 10591
rect 17221 10551 17279 10557
rect 17328 10560 17969 10588
rect 17328 10532 17356 10560
rect 17957 10557 17969 10560
rect 18003 10557 18015 10591
rect 19702 10588 19708 10600
rect 19663 10560 19708 10588
rect 17957 10551 18015 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 19797 10591 19855 10597
rect 19797 10557 19809 10591
rect 19843 10588 19855 10591
rect 20806 10588 20812 10600
rect 19843 10560 20392 10588
rect 20767 10560 20812 10588
rect 19843 10557 19855 10560
rect 19797 10551 19855 10557
rect 17310 10520 17316 10532
rect 17052 10492 17316 10520
rect 17310 10480 17316 10492
rect 17368 10480 17374 10532
rect 17420 10492 17816 10520
rect 17420 10452 17448 10492
rect 17678 10452 17684 10464
rect 16500 10424 17448 10452
rect 17639 10424 17684 10452
rect 17678 10412 17684 10424
rect 17736 10412 17742 10464
rect 17788 10452 17816 10492
rect 18966 10480 18972 10532
rect 19024 10520 19030 10532
rect 19150 10520 19156 10532
rect 19024 10492 19156 10520
rect 19024 10480 19030 10492
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 20364 10529 20392 10560
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 20916 10597 20944 10628
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 20349 10523 20407 10529
rect 20349 10489 20361 10523
rect 20395 10489 20407 10523
rect 21634 10520 21640 10532
rect 20349 10483 20407 10489
rect 20456 10492 21640 10520
rect 20456 10452 20484 10492
rect 21634 10480 21640 10492
rect 21692 10480 21698 10532
rect 17788 10424 20484 10452
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2501 10251 2559 10257
rect 2501 10217 2513 10251
rect 2547 10248 2559 10251
rect 2682 10248 2688 10260
rect 2547 10220 2688 10248
rect 2547 10217 2559 10220
rect 2501 10211 2559 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 2832 10220 2881 10248
rect 2832 10208 2838 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 5905 10251 5963 10257
rect 3936 10220 5856 10248
rect 3936 10208 3942 10220
rect 5534 10180 5540 10192
rect 5368 10152 5540 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2590 10112 2596 10124
rect 1995 10084 2596 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2590 10072 2596 10084
rect 2648 10112 2654 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 2648 10084 3433 10112
rect 2648 10072 2654 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 3421 10075 3479 10081
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5368 10121 5396 10152
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5828 10180 5856 10220
rect 5905 10217 5917 10251
rect 5951 10248 5963 10251
rect 6638 10248 6644 10260
rect 5951 10220 6644 10248
rect 5951 10217 5963 10220
rect 5905 10211 5963 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 8018 10248 8024 10260
rect 7979 10220 8024 10248
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 9030 10208 9036 10260
rect 9088 10248 9094 10260
rect 9214 10248 9220 10260
rect 9088 10220 9220 10248
rect 9088 10208 9094 10220
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 11698 10248 11704 10260
rect 9364 10220 11704 10248
rect 9364 10208 9370 10220
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 13262 10248 13268 10260
rect 12575 10220 13268 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 13412 10220 13737 10248
rect 13412 10208 13418 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 13725 10211 13783 10217
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16724 10220 17049 10248
rect 16724 10208 16730 10220
rect 17037 10217 17049 10220
rect 17083 10248 17095 10251
rect 18138 10248 18144 10260
rect 17083 10220 18144 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 18966 10248 18972 10260
rect 18831 10220 18972 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 20070 10248 20076 10260
rect 20031 10220 20076 10248
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20864 10220 20913 10248
rect 20864 10208 20870 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 5828 10152 6960 10180
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 5353 10075 5411 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 4338 10044 4344 10056
rect 3375 10016 4344 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 5902 10044 5908 10056
rect 4755 10016 5908 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 6052 10016 6377 10044
rect 6052 10004 6058 10016
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 6932 10044 6960 10152
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7745 10183 7803 10189
rect 7745 10180 7757 10183
rect 7064 10152 7757 10180
rect 7064 10140 7070 10152
rect 7745 10149 7757 10152
rect 7791 10180 7803 10183
rect 8202 10180 8208 10192
rect 7791 10152 8208 10180
rect 7791 10149 7803 10152
rect 7745 10143 7803 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 10134 10180 10140 10192
rect 9508 10152 10140 10180
rect 7374 10112 7380 10124
rect 7335 10084 7380 10112
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 8570 10112 8576 10124
rect 8531 10084 8576 10112
rect 8570 10072 8576 10084
rect 8628 10072 8634 10124
rect 9508 10121 9536 10152
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 10778 10180 10784 10192
rect 10739 10152 10784 10180
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 10962 10140 10968 10192
rect 11020 10180 11026 10192
rect 13630 10180 13636 10192
rect 11020 10152 12296 10180
rect 11020 10140 11026 10152
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 9640 10084 9685 10112
rect 9640 10072 9646 10084
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10318 10112 10324 10124
rect 10275 10084 10324 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10560 10084 11253 10112
rect 10560 10072 10566 10084
rect 11241 10081 11253 10084
rect 11287 10112 11299 10115
rect 11330 10112 11336 10124
rect 11287 10084 11336 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10081 11483 10115
rect 11882 10112 11888 10124
rect 11843 10084 11888 10112
rect 11425 10075 11483 10081
rect 9677 10047 9735 10053
rect 6932 10016 9545 10044
rect 6365 10007 6423 10013
rect 3237 9979 3295 9985
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 4522 9976 4528 9988
rect 3283 9948 4528 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5537 9979 5595 9985
rect 5537 9976 5549 9979
rect 5092 9948 5549 9976
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 2130 9868 2136 9920
rect 2188 9908 2194 9920
rect 2188 9880 2233 9908
rect 2188 9868 2194 9880
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 5092 9917 5120 9948
rect 5537 9945 5549 9948
rect 5583 9945 5595 9979
rect 5537 9939 5595 9945
rect 6457 9979 6515 9985
rect 6457 9945 6469 9979
rect 6503 9976 6515 9979
rect 6914 9976 6920 9988
rect 6503 9948 6920 9976
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 6914 9936 6920 9948
rect 6972 9936 6978 9988
rect 7193 9979 7251 9985
rect 7193 9945 7205 9979
rect 7239 9976 7251 9979
rect 7558 9976 7564 9988
rect 7239 9948 7564 9976
rect 7239 9945 7251 9948
rect 7193 9939 7251 9945
rect 7558 9936 7564 9948
rect 7616 9976 7622 9988
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7616 9948 7941 9976
rect 7616 9936 7622 9948
rect 7929 9945 7941 9948
rect 7975 9976 7987 9979
rect 9030 9976 9036 9988
rect 7975 9948 9036 9976
rect 7975 9945 7987 9948
rect 7929 9939 7987 9945
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 4249 9911 4307 9917
rect 4249 9908 4261 9911
rect 3108 9880 4261 9908
rect 3108 9868 3114 9880
rect 4249 9877 4261 9880
rect 4295 9908 4307 9911
rect 4617 9911 4675 9917
rect 4617 9908 4629 9911
rect 4295 9880 4629 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 4617 9877 4629 9880
rect 4663 9877 4675 9911
rect 4617 9871 4675 9877
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9877 5135 9911
rect 5077 9871 5135 9877
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 5997 9911 6055 9917
rect 5997 9908 6009 9911
rect 5491 9880 6009 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5997 9877 6009 9880
rect 6043 9877 6055 9911
rect 6822 9908 6828 9920
rect 6783 9880 6828 9908
rect 5997 9871 6055 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 8386 9908 8392 9920
rect 7340 9880 7385 9908
rect 8347 9880 8392 9908
rect 7340 9868 7346 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9517 9908 9545 10016
rect 9677 10013 9689 10047
rect 9723 10044 9735 10047
rect 9784 10044 9812 10072
rect 9723 10016 9812 10044
rect 9723 10013 9735 10016
rect 9677 10007 9735 10013
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10597 10047 10655 10053
rect 10597 10044 10609 10047
rect 10100 10016 10609 10044
rect 10100 10004 10106 10016
rect 10597 10013 10609 10016
rect 10643 10044 10655 10047
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 10643 10016 11161 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 11440 10044 11468 10075
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 12032 10084 12081 10112
rect 12032 10072 12038 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 12158 10044 12164 10056
rect 11440 10016 12164 10044
rect 11149 10007 11207 10013
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 12268 10044 12296 10152
rect 12728 10152 13636 10180
rect 12728 10121 12756 10152
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 14829 10183 14887 10189
rect 14829 10149 14841 10183
rect 14875 10180 14887 10183
rect 16758 10180 16764 10192
rect 14875 10152 16764 10180
rect 14875 10149 14887 10152
rect 14829 10143 14887 10149
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 18616 10180 18644 10208
rect 20438 10180 20444 10192
rect 18616 10152 20444 10180
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 12894 10112 12900 10124
rect 12855 10084 12900 10112
rect 12713 10075 12771 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 14182 10112 14188 10124
rect 14143 10084 14188 10112
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15933 10115 15991 10121
rect 15933 10081 15945 10115
rect 15979 10112 15991 10115
rect 16206 10112 16212 10124
rect 15979 10084 16212 10112
rect 15979 10081 15991 10084
rect 15933 10075 15991 10081
rect 12989 10047 13047 10053
rect 12268 10016 12434 10044
rect 10060 9976 10088 10004
rect 9876 9948 10088 9976
rect 12406 9976 12434 10016
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13170 10044 13176 10056
rect 13035 10016 13176 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13633 10047 13691 10053
rect 13633 10044 13645 10047
rect 13596 10016 13645 10044
rect 13596 10004 13602 10016
rect 13633 10013 13645 10016
rect 13679 10044 13691 10047
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13679 10016 14473 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 15948 10044 15976 10075
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 19521 10115 19579 10121
rect 16439 10084 16712 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 16482 10044 16488 10056
rect 15519 10016 15976 10044
rect 16443 10016 16488 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16684 10044 16712 10084
rect 19521 10081 19533 10115
rect 19567 10112 19579 10115
rect 19610 10112 19616 10124
rect 19567 10084 19616 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 20272 10121 20300 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 20257 10115 20315 10121
rect 20257 10081 20269 10115
rect 20303 10081 20315 10115
rect 20257 10075 20315 10081
rect 16758 10044 16764 10056
rect 16684 10016 16764 10044
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17126 10044 17132 10056
rect 17052 10016 17132 10044
rect 14918 9976 14924 9988
rect 12406 9948 14924 9976
rect 9876 9908 9904 9948
rect 14918 9936 14924 9948
rect 14976 9976 14982 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14976 9948 15393 9976
rect 14976 9936 14982 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 16577 9979 16635 9985
rect 16577 9945 16589 9979
rect 16623 9976 16635 9979
rect 17052 9976 17080 10016
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 17310 10044 17316 10056
rect 17267 10016 17316 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 18230 10004 18236 10056
rect 18288 10044 18294 10056
rect 20441 10047 20499 10053
rect 20441 10044 20453 10047
rect 18288 10016 20453 10044
rect 18288 10004 18294 10016
rect 20441 10013 20453 10016
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 17494 9985 17500 9988
rect 16623 9948 17080 9976
rect 17466 9979 17500 9985
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 17466 9945 17478 9979
rect 17552 9976 17558 9988
rect 17770 9976 17776 9988
rect 17552 9948 17776 9976
rect 17466 9939 17500 9945
rect 17494 9936 17500 9939
rect 17552 9936 17558 9948
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 19613 9979 19671 9985
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 20806 9976 20812 9988
rect 19659 9948 20812 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 8536 9880 8581 9908
rect 9517 9880 9904 9908
rect 8536 9868 8542 9880
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 11701 9911 11759 9917
rect 10100 9880 10145 9908
rect 10100 9868 10106 9880
rect 11701 9877 11713 9911
rect 11747 9908 11759 9911
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 11747 9880 12173 9908
rect 11747 9877 11759 9880
rect 11701 9871 11759 9877
rect 12161 9877 12173 9880
rect 12207 9908 12219 9911
rect 13262 9908 13268 9920
rect 12207 9880 13268 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 13357 9911 13415 9917
rect 13357 9877 13369 9911
rect 13403 9908 13415 9911
rect 13814 9908 13820 9920
rect 13403 9880 13820 9908
rect 13403 9877 13415 9880
rect 13357 9871 13415 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 14366 9908 14372 9920
rect 14327 9880 14372 9908
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 16666 9908 16672 9920
rect 14792 9880 16672 9908
rect 14792 9868 14798 9880
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19760 9880 19805 9908
rect 19760 9868 19766 9880
rect 20530 9868 20536 9920
rect 20588 9908 20594 9920
rect 20588 9880 20633 9908
rect 20588 9868 20594 9880
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20956 9880 21005 9908
rect 20956 9868 20962 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 21266 9908 21272 9920
rect 21227 9880 21272 9908
rect 20993 9871 21051 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 21545 9911 21603 9917
rect 21545 9877 21557 9911
rect 21591 9908 21603 9911
rect 21634 9908 21640 9920
rect 21591 9880 21640 9908
rect 21591 9877 21603 9880
rect 21545 9871 21603 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1765 9707 1823 9713
rect 1765 9673 1777 9707
rect 1811 9704 1823 9707
rect 2038 9704 2044 9716
rect 1811 9676 2044 9704
rect 1811 9673 1823 9676
rect 1765 9667 1823 9673
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 4157 9707 4215 9713
rect 4157 9673 4169 9707
rect 4203 9704 4215 9707
rect 4430 9704 4436 9716
rect 4203 9676 4436 9704
rect 4203 9673 4215 9676
rect 4157 9667 4215 9673
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 2838 9639 2896 9645
rect 2838 9636 2850 9639
rect 2648 9608 2850 9636
rect 2648 9596 2654 9608
rect 2838 9605 2850 9608
rect 2884 9605 2896 9639
rect 2838 9599 2896 9605
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 2096 9540 2145 9568
rect 2096 9528 2102 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 4172 9568 4200 9667
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4580 9676 4629 9704
rect 4580 9664 4586 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4617 9667 4675 9673
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 5132 9676 5177 9704
rect 5132 9664 5138 9676
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5718 9704 5724 9716
rect 5592 9676 5724 9704
rect 5592 9664 5598 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 7929 9707 7987 9713
rect 7929 9704 7941 9707
rect 7668 9676 7941 9704
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 2133 9531 2191 9537
rect 2608 9540 4200 9568
rect 4632 9608 5825 9636
rect 2222 9500 2228 9512
rect 2183 9472 2228 9500
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2608 9509 2636 9540
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9469 2651 9503
rect 2593 9463 2651 9469
rect 1670 9392 1676 9444
rect 1728 9432 1734 9444
rect 2332 9432 2360 9463
rect 4632 9432 4660 9608
rect 5813 9605 5825 9608
rect 5859 9636 5871 9639
rect 5994 9636 6000 9648
rect 5859 9608 6000 9636
rect 5859 9605 5871 9608
rect 5813 9599 5871 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6604 9608 6837 9636
rect 6604 9596 6610 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 7668 9636 7696 9676
rect 7929 9673 7941 9676
rect 7975 9673 7987 9707
rect 8294 9704 8300 9716
rect 8255 9676 8300 9704
rect 7929 9667 7987 9673
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 8628 9676 9781 9704
rect 8628 9664 8634 9676
rect 9769 9673 9781 9676
rect 9815 9704 9827 9707
rect 10594 9704 10600 9716
rect 9815 9676 10600 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 10836 9676 11069 9704
rect 10836 9664 10842 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 13446 9704 13452 9716
rect 11756 9676 13452 9704
rect 11756 9664 11762 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14182 9704 14188 9716
rect 13556 9676 14188 9704
rect 8588 9636 8616 9664
rect 8662 9645 8668 9648
rect 6825 9599 6883 9605
rect 7484 9608 7696 9636
rect 7760 9608 8616 9636
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 6733 9571 6791 9577
rect 5031 9540 5488 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 1728 9404 2360 9432
rect 1728 9392 1734 9404
rect 2332 9364 2360 9404
rect 4448 9404 4660 9432
rect 4448 9376 4476 9404
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 5184 9432 5212 9463
rect 5460 9441 5488 9540
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 7006 9568 7012 9580
rect 6779 9540 7012 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7484 9512 7512 9608
rect 5902 9500 5908 9512
rect 5863 9472 5908 9500
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6917 9503 6975 9509
rect 6052 9472 6097 9500
rect 6052 9460 6058 9472
rect 6917 9469 6929 9503
rect 6963 9500 6975 9503
rect 7374 9500 7380 9512
rect 6963 9472 7380 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 5040 9404 5212 9432
rect 5445 9435 5503 9441
rect 5040 9392 5046 9404
rect 5445 9401 5457 9435
rect 5491 9401 5503 9435
rect 6012 9432 6040 9460
rect 6932 9432 6960 9463
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7760 9509 7788 9608
rect 8656 9599 8668 9645
rect 8720 9636 8726 9648
rect 10410 9636 10416 9648
rect 8720 9608 8756 9636
rect 10371 9608 10416 9636
rect 8662 9596 8668 9599
rect 8720 9596 8726 9608
rect 10410 9596 10416 9608
rect 10468 9636 10474 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 10468 9608 11989 9636
rect 10468 9596 10474 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 13556 9636 13584 9676
rect 14182 9664 14188 9676
rect 14240 9704 14246 9716
rect 16298 9704 16304 9716
rect 14240 9676 16304 9704
rect 14240 9664 14246 9676
rect 16298 9664 16304 9676
rect 16356 9704 16362 9716
rect 16356 9686 16528 9704
rect 16356 9676 16488 9686
rect 16356 9664 16362 9676
rect 11977 9599 12035 9605
rect 12636 9608 13584 9636
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 10965 9571 11023 9577
rect 8076 9540 10088 9568
rect 8076 9528 8082 9540
rect 7745 9503 7803 9509
rect 7524 9472 7569 9500
rect 7524 9460 7530 9472
rect 7745 9469 7757 9503
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 8294 9500 8300 9512
rect 7883 9472 8300 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 6012 9404 6960 9432
rect 5445 9395 5503 9401
rect 3970 9364 3976 9376
rect 2332 9336 3976 9364
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4430 9364 4436 9376
rect 4387 9336 4436 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4890 9364 4896 9376
rect 4571 9336 4896 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5074 9324 5080 9376
rect 5132 9364 5138 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5132 9336 6377 9364
rect 5132 9324 5138 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 6972 9336 7297 9364
rect 6972 9324 6978 9336
rect 7285 9333 7297 9336
rect 7331 9364 7343 9367
rect 7742 9364 7748 9376
rect 7331 9336 7748 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8404 9364 8432 9463
rect 10060 9432 10088 9540
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11882 9568 11888 9580
rect 11011 9540 11560 9568
rect 11843 9540 11888 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10560 9472 11161 9500
rect 10560 9460 10566 9472
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 11532 9441 11560 9540
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12158 9500 12164 9512
rect 12119 9472 12164 9500
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 12636 9509 12664 9608
rect 13630 9596 13636 9648
rect 13688 9645 13694 9648
rect 13688 9639 13752 9645
rect 13688 9605 13706 9639
rect 13740 9605 13752 9639
rect 14918 9636 14924 9648
rect 14879 9608 14924 9636
rect 13688 9599 13752 9605
rect 13688 9596 13694 9599
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 16482 9634 16488 9676
rect 16540 9634 16546 9686
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 17954 9704 17960 9716
rect 16908 9676 17960 9704
rect 16908 9664 16914 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 18966 9704 18972 9716
rect 18748 9676 18972 9704
rect 18748 9664 18754 9676
rect 18966 9664 18972 9676
rect 19024 9664 19030 9716
rect 19702 9664 19708 9716
rect 19760 9704 19766 9716
rect 19889 9707 19947 9713
rect 19889 9704 19901 9707
rect 19760 9676 19901 9704
rect 19760 9664 19766 9676
rect 19889 9673 19901 9676
rect 19935 9673 19947 9707
rect 19889 9667 19947 9673
rect 20717 9707 20775 9713
rect 20717 9673 20729 9707
rect 20763 9704 20775 9707
rect 20806 9704 20812 9716
rect 20763 9676 20812 9704
rect 20763 9673 20775 9676
rect 20717 9667 20775 9673
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17034 9636 17040 9648
rect 16632 9608 17040 9636
rect 16632 9596 16638 9608
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 17218 9596 17224 9648
rect 17276 9596 17282 9648
rect 17862 9636 17868 9648
rect 17604 9608 17868 9636
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 14608 9540 15485 9568
rect 14608 9528 14614 9540
rect 15473 9537 15485 9540
rect 15519 9537 15531 9571
rect 17236 9568 17264 9596
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 15473 9531 15531 9537
rect 16408 9540 17325 9568
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9469 12679 9503
rect 12621 9463 12679 9469
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 11517 9435 11575 9441
rect 10060 9404 11468 9432
rect 9398 9364 9404 9376
rect 8404 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9364 9462 9376
rect 9861 9367 9919 9373
rect 9861 9364 9873 9367
rect 9456 9336 9873 9364
rect 9456 9324 9462 9336
rect 9861 9333 9873 9336
rect 9907 9333 9919 9367
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 9861 9327 9919 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11440 9364 11468 9404
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12342 9432 12348 9444
rect 11756 9404 12348 9432
rect 11756 9392 11762 9404
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 12250 9364 12256 9376
rect 11440 9336 12256 9364
rect 12250 9324 12256 9336
rect 12308 9364 12314 9376
rect 12728 9364 12756 9463
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 13412 9472 13461 9500
rect 13412 9460 13418 9472
rect 13449 9469 13461 9472
rect 13495 9469 13507 9503
rect 15194 9500 15200 9512
rect 15155 9472 15200 9500
rect 13449 9463 13507 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9500 15439 9503
rect 15654 9500 15660 9512
rect 15427 9472 15660 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15286 9432 15292 9444
rect 14752 9404 15292 9432
rect 12308 9336 12756 9364
rect 13173 9367 13231 9373
rect 12308 9324 12314 9336
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 14752 9364 14780 9404
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 13219 9336 14780 9364
rect 14829 9367 14887 9373
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15010 9364 15016 9376
rect 14875 9336 15016 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 15470 9364 15476 9376
rect 15252 9336 15476 9364
rect 15252 9324 15258 9336
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16022 9364 16028 9376
rect 15887 9336 16028 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16408 9373 16436 9540
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 17604 9568 17632 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19518 9596 19524 9648
rect 19576 9645 19582 9648
rect 19576 9636 19588 9645
rect 20349 9639 20407 9645
rect 20349 9636 20361 9639
rect 19576 9608 19621 9636
rect 19720 9608 20361 9636
rect 19576 9599 19588 9608
rect 19576 9596 19582 9599
rect 19720 9568 19748 9608
rect 20349 9605 20361 9608
rect 20395 9605 20407 9639
rect 21174 9636 21180 9648
rect 20349 9599 20407 9605
rect 20548 9608 21180 9636
rect 20254 9568 20260 9580
rect 17552 9540 17632 9568
rect 17696 9540 19748 9568
rect 20215 9540 20260 9568
rect 17552 9528 17558 9540
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16540 9472 17049 9500
rect 16540 9460 16546 9472
rect 17037 9469 17049 9472
rect 17083 9469 17095 9503
rect 17037 9463 17095 9469
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17236 9432 17264 9463
rect 17696 9441 17724 9540
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 17957 9503 18015 9509
rect 17957 9500 17969 9503
rect 17920 9472 17969 9500
rect 17920 9460 17926 9472
rect 17957 9469 17969 9472
rect 18003 9469 18015 9503
rect 17957 9463 18015 9469
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9469 19855 9503
rect 20438 9500 20444 9512
rect 20399 9472 20444 9500
rect 19797 9463 19855 9469
rect 16684 9404 17264 9432
rect 17681 9435 17739 9441
rect 16684 9376 16712 9404
rect 17681 9401 17693 9435
rect 17727 9401 17739 9435
rect 18233 9435 18291 9441
rect 18233 9432 18245 9435
rect 17681 9395 17739 9401
rect 17880 9404 18245 9432
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 16393 9327 16451 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17880 9364 17908 9404
rect 18233 9401 18245 9404
rect 18279 9432 18291 9435
rect 18690 9432 18696 9444
rect 18279 9404 18696 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18690 9392 18696 9404
rect 18748 9392 18754 9444
rect 18046 9364 18052 9376
rect 16816 9336 17908 9364
rect 18007 9336 18052 9364
rect 16816 9324 16822 9336
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 18417 9367 18475 9373
rect 18417 9333 18429 9367
rect 18463 9364 18475 9367
rect 18506 9364 18512 9376
rect 18463 9336 18512 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 18708 9364 18736 9392
rect 19812 9364 19840 9463
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 20548 9500 20576 9608
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 21085 9571 21143 9577
rect 21085 9568 21097 9571
rect 20680 9540 21097 9568
rect 20680 9528 20686 9540
rect 21085 9537 21097 9540
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 20806 9500 20812 9512
rect 20548 9472 20812 9500
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 21174 9500 21180 9512
rect 21135 9472 21180 9500
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9469 21327 9503
rect 21269 9463 21327 9469
rect 20456 9432 20484 9460
rect 21284 9432 21312 9463
rect 20456 9404 21312 9432
rect 18708 9336 19840 9364
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2280 9132 2329 9160
rect 2280 9120 2286 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4396 9132 4445 9160
rect 4396 9120 4402 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6086 9160 6092 9172
rect 5868 9132 5948 9160
rect 6047 9132 6092 9160
rect 5868 9120 5874 9132
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 5920 9092 5948 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 7006 9160 7012 9172
rect 6411 9132 7012 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 7006 9120 7012 9132
rect 7064 9160 7070 9172
rect 7282 9160 7288 9172
rect 7064 9132 7144 9160
rect 7243 9132 7288 9160
rect 7064 9120 7070 9132
rect 6454 9092 6460 9104
rect 3476 9064 5856 9092
rect 5920 9064 6460 9092
rect 3476 9052 3482 9064
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2746 8996 2881 9024
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 2746 8956 2774 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 3326 9024 3332 9036
rect 3287 8996 3332 9024
rect 2869 8987 2927 8993
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4338 9024 4344 9036
rect 3927 8996 4344 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 3142 8956 3148 8968
rect 2648 8928 2774 8956
rect 3103 8928 3148 8956
rect 2648 8916 2654 8928
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 1636 8860 1869 8888
rect 1636 8848 1642 8860
rect 1857 8857 1869 8860
rect 1903 8857 1915 8891
rect 1857 8851 1915 8857
rect 2685 8891 2743 8897
rect 2685 8857 2697 8891
rect 2731 8888 2743 8891
rect 2866 8888 2872 8900
rect 2731 8860 2872 8888
rect 2731 8857 2743 8860
rect 2685 8851 2743 8857
rect 2866 8848 2872 8860
rect 2924 8888 2930 8900
rect 3234 8888 3240 8900
rect 2924 8860 3240 8888
rect 2924 8848 2930 8860
rect 3234 8848 3240 8860
rect 3292 8888 3298 8900
rect 3510 8888 3516 8900
rect 3292 8860 3516 8888
rect 3292 8848 3298 8860
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 2130 8780 2136 8832
rect 2188 8820 2194 8832
rect 2225 8823 2283 8829
rect 2225 8820 2237 8823
rect 2188 8792 2237 8820
rect 2188 8780 2194 8792
rect 2225 8789 2237 8792
rect 2271 8789 2283 8823
rect 2225 8783 2283 8789
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 3896 8820 3924 8987
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 4798 9024 4804 9036
rect 4396 8996 4804 9024
rect 4396 8984 4402 8996
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5718 9024 5724 9036
rect 5132 8996 5724 9024
rect 5132 8984 5138 8996
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5828 9033 5856 9064
rect 6454 9052 6460 9064
rect 6512 9052 6518 9104
rect 7116 9092 7144 9132
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 8018 9160 8024 9172
rect 7392 9132 8024 9160
rect 7392 9092 7420 9132
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8444 9132 9045 9160
rect 8444 9120 8450 9132
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9033 9123 9091 9129
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9180 9132 10241 9160
rect 9180 9120 9186 9132
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10502 9160 10508 9172
rect 10463 9132 10508 9160
rect 10229 9123 10287 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 11974 9160 11980 9172
rect 10980 9132 11980 9160
rect 7116 9064 7420 9092
rect 7300 9036 7328 9064
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 8757 9095 8815 9101
rect 8757 9092 8769 9095
rect 8720 9064 8769 9092
rect 8720 9052 8726 9064
rect 8757 9061 8769 9064
rect 8803 9092 8815 9095
rect 8803 9064 9628 9092
rect 8803 9061 8815 9064
rect 8757 9055 8815 9061
rect 9600 9036 9628 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 9732 9064 10057 9092
rect 9732 9052 9738 9064
rect 10045 9061 10057 9064
rect 10091 9092 10103 9095
rect 10980 9092 11008 9132
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12250 9160 12256 9172
rect 12211 9132 12256 9160
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12802 9160 12808 9172
rect 12575 9132 12808 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9160 13507 9163
rect 14366 9160 14372 9172
rect 13495 9132 14372 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 17954 9160 17960 9172
rect 14844 9132 17960 9160
rect 10091 9064 11008 9092
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 11882 9052 11888 9104
rect 11940 9092 11946 9104
rect 11940 9064 12020 9092
rect 11940 9052 11946 9064
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 5902 9024 5908 9036
rect 5859 8996 5908 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 6604 8996 6653 9024
rect 6604 8984 6610 8996
rect 6641 8993 6653 8996
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 9582 9024 9588 9036
rect 9495 8996 9588 9024
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4430 8956 4436 8968
rect 4028 8928 4436 8956
rect 4028 8916 4034 8928
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 6822 8956 6828 8968
rect 4939 8928 6828 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 9401 8959 9459 8965
rect 7484 8928 8524 8956
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8888 4399 8891
rect 4614 8888 4620 8900
rect 4387 8860 4620 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 4614 8848 4620 8860
rect 4672 8888 4678 8900
rect 5074 8888 5080 8900
rect 4672 8860 5080 8888
rect 4672 8848 4678 8860
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 7484 8888 7512 8928
rect 5408 8860 7512 8888
rect 7644 8891 7702 8897
rect 5408 8848 5414 8860
rect 7644 8857 7656 8891
rect 7690 8888 7702 8891
rect 8202 8888 8208 8900
rect 7690 8860 8208 8888
rect 7690 8857 7702 8860
rect 7644 8851 7702 8857
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 4798 8820 4804 8832
rect 2823 8792 3924 8820
rect 4759 8792 4804 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 5040 8792 5273 8820
rect 5040 8780 5046 8792
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 5718 8820 5724 8832
rect 5675 8792 5724 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6822 8820 6828 8832
rect 6512 8792 6828 8820
rect 6512 8780 6518 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 8386 8820 8392 8832
rect 6963 8792 8392 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8496 8820 8524 8928
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9692 8956 9720 9052
rect 11992 9033 12020 9064
rect 13170 9052 13176 9104
rect 13228 9092 13234 9104
rect 14844 9092 14872 9132
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 20714 9160 20720 9172
rect 18432 9132 20208 9160
rect 20675 9132 20720 9160
rect 13228 9064 14872 9092
rect 13228 9052 13234 9064
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 12805 9027 12863 9033
rect 12805 8993 12817 9027
rect 12851 8993 12863 9027
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12805 8987 12863 8993
rect 9447 8928 9720 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11204 8928 11897 8956
rect 11204 8916 11210 8928
rect 11885 8925 11897 8928
rect 11931 8925 11943 8959
rect 12820 8956 12848 8987
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 14550 9024 14556 9036
rect 13136 8996 14556 9024
rect 13136 8984 13142 8996
rect 14550 8984 14556 8996
rect 14608 9024 14614 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14608 8996 14749 9024
rect 14608 8984 14614 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 15102 9024 15108 9036
rect 15015 8996 15108 9024
rect 14737 8987 14795 8993
rect 14642 8956 14648 8968
rect 12820 8928 14648 8956
rect 11885 8919 11943 8925
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9766 8888 9772 8900
rect 8720 8860 9772 8888
rect 8720 8848 8726 8860
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 11640 8891 11698 8897
rect 11640 8857 11652 8891
rect 11686 8888 11698 8891
rect 12158 8888 12164 8900
rect 11686 8860 12164 8888
rect 11686 8857 11698 8860
rect 11640 8851 11698 8857
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 15028 8888 15056 8996
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 16592 8996 16896 9024
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 15556 8959 15614 8965
rect 15556 8925 15568 8959
rect 15602 8956 15614 8959
rect 16592 8956 16620 8996
rect 16758 8956 16764 8968
rect 15602 8928 16620 8956
rect 16719 8928 16764 8956
rect 15602 8925 15614 8928
rect 15556 8919 15614 8925
rect 12584 8860 15056 8888
rect 12584 8848 12590 8860
rect 9493 8823 9551 8829
rect 9493 8820 9505 8823
rect 8496 8792 9505 8820
rect 9493 8789 9505 8792
rect 9539 8820 9551 8823
rect 9953 8823 10011 8829
rect 9953 8820 9965 8823
rect 9539 8792 9965 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 9953 8789 9965 8792
rect 9999 8820 10011 8823
rect 11790 8820 11796 8832
rect 9999 8792 11796 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 13078 8820 13084 8832
rect 13039 8792 13084 8820
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 13630 8820 13636 8832
rect 13412 8792 13636 8820
rect 13412 8780 13418 8792
rect 13630 8780 13636 8792
rect 13688 8820 13694 8832
rect 14458 8820 14464 8832
rect 13688 8792 14464 8820
rect 13688 8780 13694 8792
rect 14458 8780 14464 8792
rect 14516 8820 14522 8832
rect 14921 8823 14979 8829
rect 14921 8820 14933 8823
rect 14516 8792 14933 8820
rect 14516 8780 14522 8792
rect 14921 8789 14933 8792
rect 14967 8820 14979 8823
rect 15304 8820 15332 8919
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 15571 8888 15599 8919
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16868 8956 16896 8996
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 18432 9033 18460 9132
rect 20180 9092 20208 9132
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 20625 9095 20683 9101
rect 20625 9092 20637 9095
rect 20180 9064 20637 9092
rect 20625 9061 20637 9064
rect 20671 9092 20683 9095
rect 20806 9092 20812 9104
rect 20671 9064 20812 9092
rect 20671 9061 20683 9064
rect 20625 9055 20683 9061
rect 20806 9052 20812 9064
rect 20864 9052 20870 9104
rect 18417 9027 18475 9033
rect 18417 9024 18429 9027
rect 17828 8996 18429 9024
rect 17828 8984 17834 8996
rect 18417 8993 18429 8996
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 18647 8996 19380 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 18506 8956 18512 8968
rect 16868 8928 18512 8956
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 18690 8916 18696 8968
rect 18748 8956 18754 8968
rect 19242 8956 19248 8968
rect 18748 8928 19248 8956
rect 18748 8916 18754 8928
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19352 8956 19380 8996
rect 20438 8984 20444 9036
rect 20496 9024 20502 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20496 8996 21281 9024
rect 20496 8984 20502 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 19886 8956 19892 8968
rect 19352 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21358 8956 21364 8968
rect 21131 8928 21364 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 17006 8891 17064 8897
rect 17006 8888 17018 8891
rect 15528 8860 15599 8888
rect 16684 8860 17018 8888
rect 15528 8848 15534 8860
rect 14967 8792 15332 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16574 8820 16580 8832
rect 15988 8792 16580 8820
rect 15988 8780 15994 8792
rect 16574 8780 16580 8792
rect 16632 8820 16638 8832
rect 16684 8829 16712 8860
rect 17006 8857 17018 8860
rect 17052 8857 17064 8891
rect 17006 8851 17064 8857
rect 18414 8848 18420 8900
rect 18472 8888 18478 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 18472 8860 19502 8888
rect 18472 8848 18478 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 21177 8891 21235 8897
rect 21177 8888 21189 8891
rect 19490 8851 19548 8857
rect 20180 8860 21189 8888
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16632 8792 16681 8820
rect 16632 8780 16638 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 18141 8823 18199 8829
rect 18141 8820 18153 8823
rect 17276 8792 18153 8820
rect 17276 8780 17282 8792
rect 18141 8789 18153 8792
rect 18187 8789 18199 8823
rect 18690 8820 18696 8832
rect 18651 8792 18696 8820
rect 18141 8783 18199 8789
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 19061 8823 19119 8829
rect 19061 8789 19073 8823
rect 19107 8820 19119 8823
rect 20180 8820 20208 8860
rect 21177 8857 21189 8860
rect 21223 8857 21235 8891
rect 21177 8851 21235 8857
rect 19107 8792 20208 8820
rect 19107 8789 19119 8792
rect 19061 8783 19119 8789
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 2041 8619 2099 8625
rect 2041 8616 2053 8619
rect 1820 8588 2053 8616
rect 1820 8576 1826 8588
rect 2041 8585 2053 8588
rect 2087 8585 2099 8619
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2041 8579 2099 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 4522 8616 4528 8628
rect 2556 8588 2601 8616
rect 4483 8588 4528 8616
rect 2556 8576 2562 8588
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4856 8588 5089 8616
rect 4856 8576 4862 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 5408 8588 5549 8616
rect 5408 8576 5414 8588
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 5537 8579 5595 8585
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5868 8588 5917 8616
rect 5868 8576 5874 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 1854 8548 1860 8560
rect 1627 8520 1860 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 1854 8508 1860 8520
rect 1912 8548 1918 8560
rect 2424 8548 2452 8576
rect 1912 8520 2452 8548
rect 1912 8508 1918 8520
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 5994 8548 6000 8560
rect 2648 8520 6000 8548
rect 2648 8508 2654 8520
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2866 8480 2872 8492
rect 1995 8452 2872 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3234 8489 3240 8492
rect 3228 8480 3240 8489
rect 3195 8452 3240 8480
rect 3228 8443 3240 8452
rect 3234 8440 3240 8443
rect 3292 8440 3298 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4614 8480 4620 8492
rect 4212 8452 4620 8480
rect 4212 8440 4218 8452
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5442 8480 5448 8492
rect 4847 8452 5448 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 1728 8384 1777 8412
rect 1728 8372 1734 8384
rect 1765 8381 1777 8384
rect 1811 8412 1823 8415
rect 2498 8412 2504 8424
rect 1811 8384 2504 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2590 8372 2596 8424
rect 2648 8412 2654 8424
rect 2961 8415 3019 8421
rect 2648 8384 2693 8412
rect 2648 8372 2654 8384
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 4522 8412 4528 8424
rect 2961 8375 3019 8381
rect 3988 8384 4528 8412
rect 1210 8304 1216 8356
rect 1268 8344 1274 8356
rect 2774 8344 2780 8356
rect 1268 8316 2780 8344
rect 1268 8304 1274 8316
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 2130 8236 2136 8288
rect 2188 8276 2194 8288
rect 2976 8276 3004 8375
rect 3988 8276 4016 8384
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5350 8412 5356 8424
rect 5031 8384 5356 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5644 8421 5672 8520
rect 5994 8508 6000 8520
rect 6052 8548 6058 8560
rect 6380 8548 6408 8579
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8536 8588 8953 8616
rect 8536 8576 8542 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 9180 8588 9321 8616
rect 9180 8576 9186 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 9309 8579 9367 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 12805 8619 12863 8625
rect 10428 8588 11284 8616
rect 7929 8551 7987 8557
rect 6052 8520 6408 8548
rect 6472 8520 7880 8548
rect 6052 8508 6058 8520
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 6270 8480 6276 8492
rect 5776 8452 6276 8480
rect 5776 8440 5782 8452
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 6086 8412 6092 8424
rect 6047 8384 6092 8412
rect 5629 8375 5687 8381
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4341 8347 4399 8353
rect 4120 8316 4200 8344
rect 4120 8304 4126 8316
rect 2188 8248 4016 8276
rect 4172 8276 4200 8316
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4798 8344 4804 8356
rect 4387 8316 4804 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5368 8344 5396 8372
rect 6472 8344 6500 8520
rect 7478 8483 7536 8489
rect 7478 8480 7490 8483
rect 6748 8452 7490 8480
rect 5368 8316 6500 8344
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 6748 8344 6776 8452
rect 7478 8449 7490 8452
rect 7524 8449 7536 8483
rect 7852 8480 7880 8520
rect 7929 8517 7941 8551
rect 7975 8548 7987 8551
rect 8386 8548 8392 8560
rect 7975 8520 8392 8548
rect 7975 8517 7987 8520
rect 7929 8511 7987 8517
rect 8386 8508 8392 8520
rect 8444 8548 8450 8560
rect 9490 8548 9496 8560
rect 8444 8520 9496 8548
rect 8444 8508 8450 8520
rect 9490 8508 9496 8520
rect 9548 8548 9554 8560
rect 10428 8548 10456 8588
rect 9548 8520 10456 8548
rect 9548 8508 9554 8520
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 10893 8551 10951 8557
rect 10893 8548 10905 8551
rect 10560 8520 10905 8548
rect 10560 8508 10566 8520
rect 10893 8517 10905 8520
rect 10939 8517 10951 8551
rect 10893 8511 10951 8517
rect 8202 8480 8208 8492
rect 7852 8452 8208 8480
rect 7478 8443 7536 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 8711 8452 9413 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 9401 8449 9413 8452
rect 9447 8480 9459 8483
rect 11054 8480 11060 8492
rect 9447 8452 11060 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 11256 8480 11284 8588
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 12986 8616 12992 8628
rect 12851 8588 12992 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13538 8616 13544 8628
rect 13499 8588 13544 8616
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 14332 8588 14749 8616
rect 14332 8576 14338 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 16022 8616 16028 8628
rect 15983 8588 16028 8616
rect 14737 8579 14795 8585
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 16485 8619 16543 8625
rect 16485 8585 16497 8619
rect 16531 8616 16543 8619
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16531 8588 16957 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 16945 8579 17003 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18414 8616 18420 8628
rect 18327 8588 18420 8616
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 20070 8616 20076 8628
rect 18748 8588 20076 8616
rect 18748 8576 18754 8588
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20257 8619 20315 8625
rect 20257 8585 20269 8619
rect 20303 8616 20315 8619
rect 20530 8616 20536 8628
rect 20303 8588 20536 8616
rect 20303 8585 20315 8588
rect 20257 8579 20315 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20625 8619 20683 8625
rect 20625 8585 20637 8619
rect 20671 8616 20683 8619
rect 21726 8616 21732 8628
rect 20671 8588 21732 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11756 8520 11805 8548
rect 11756 8508 11762 8520
rect 11793 8517 11805 8520
rect 11839 8548 11851 8551
rect 13354 8548 13360 8560
rect 11839 8520 13360 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 12250 8480 12256 8492
rect 11256 8452 11376 8480
rect 12211 8452 12256 8480
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7791 8384 8033 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8021 8381 8033 8384
rect 8067 8412 8079 8415
rect 9582 8412 9588 8424
rect 8067 8384 8294 8412
rect 9543 8384 9588 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 6604 8316 6776 8344
rect 6604 8304 6610 8316
rect 7006 8276 7012 8288
rect 4172 8248 7012 8276
rect 2188 8236 2194 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7760 8276 7788 8375
rect 8266 8344 8294 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 8266 8316 8892 8344
rect 7432 8248 7788 8276
rect 8297 8279 8355 8285
rect 7432 8236 7438 8248
rect 8297 8245 8309 8279
rect 8343 8276 8355 8279
rect 8478 8276 8484 8288
rect 8343 8248 8484 8276
rect 8343 8245 8355 8248
rect 8297 8239 8355 8245
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 8864 8285 8892 8316
rect 11164 8288 11192 8375
rect 11348 8344 11376 8452
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12894 8480 12900 8492
rect 12391 8452 12900 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13556 8480 13584 8576
rect 15470 8548 15476 8560
rect 14752 8520 15476 8548
rect 13219 8452 13584 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12216 8384 12449 8412
rect 12216 8372 12222 8384
rect 12437 8381 12449 8384
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 13188 8344 13216 8443
rect 13722 8440 13728 8492
rect 13780 8440 13786 8492
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 13740 8412 13768 8440
rect 13596 8384 13768 8412
rect 14645 8415 14703 8421
rect 13596 8372 13602 8384
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 14752 8412 14780 8520
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 18432 8548 18460 8576
rect 21358 8548 21364 8560
rect 15948 8520 18460 8548
rect 19306 8520 21364 8548
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 15948 8480 15976 8520
rect 16114 8480 16120 8492
rect 14829 8443 14887 8449
rect 14936 8452 15976 8480
rect 16075 8452 16120 8480
rect 14691 8384 14780 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 11348 8316 13216 8344
rect 13357 8347 13415 8353
rect 13357 8313 13369 8347
rect 13403 8344 13415 8347
rect 13722 8344 13728 8356
rect 13403 8316 13728 8344
rect 13403 8313 13415 8316
rect 13357 8307 13415 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 14185 8347 14243 8353
rect 14185 8313 14197 8347
rect 14231 8344 14243 8347
rect 14550 8344 14556 8356
rect 14231 8316 14556 8344
rect 14231 8313 14243 8316
rect 14185 8307 14243 8313
rect 14550 8304 14556 8316
rect 14608 8344 14614 8356
rect 14844 8344 14872 8443
rect 14608 8316 14872 8344
rect 14608 8304 14614 8316
rect 8849 8279 8907 8285
rect 8849 8245 8861 8279
rect 8895 8276 8907 8279
rect 9398 8276 9404 8288
rect 8895 8248 9404 8276
rect 8895 8245 8907 8248
rect 8849 8239 8907 8245
rect 9398 8236 9404 8248
rect 9456 8276 9462 8288
rect 11146 8276 11152 8288
rect 9456 8248 11152 8276
rect 9456 8236 9462 8248
rect 11146 8236 11152 8248
rect 11204 8276 11210 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 11204 8248 11253 8276
rect 11204 8236 11210 8248
rect 11241 8245 11253 8248
rect 11287 8245 11299 8279
rect 11241 8239 11299 8245
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 11885 8279 11943 8285
rect 11885 8276 11897 8279
rect 11848 8248 11897 8276
rect 11848 8236 11854 8248
rect 11885 8245 11897 8248
rect 11931 8245 11943 8279
rect 11885 8239 11943 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12802 8276 12808 8288
rect 12032 8248 12808 8276
rect 12032 8236 12038 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 12986 8276 12992 8288
rect 12947 8248 12992 8276
rect 12986 8236 12992 8248
rect 13044 8236 13050 8288
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 14274 8276 14280 8288
rect 13136 8248 14280 8276
rect 13136 8236 13142 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 14936 8276 14964 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 17000 8452 17049 8480
rect 17000 8440 17006 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 18506 8480 18512 8492
rect 17037 8443 17095 8449
rect 18156 8452 18512 8480
rect 15286 8412 15292 8424
rect 15247 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15930 8412 15936 8424
rect 15891 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17218 8412 17224 8424
rect 16899 8384 17224 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 18156 8421 18184 8452
rect 18506 8440 18512 8452
rect 18564 8480 18570 8492
rect 19306 8480 19334 8520
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 19518 8480 19524 8492
rect 19576 8489 19582 8492
rect 18564 8452 19334 8480
rect 19488 8452 19524 8480
rect 18564 8440 18570 8452
rect 19518 8440 19524 8452
rect 19576 8443 19588 8489
rect 19576 8440 19582 8443
rect 19702 8440 19708 8492
rect 19760 8480 19766 8492
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 19760 8452 19809 8480
rect 19760 8440 19766 8452
rect 19797 8449 19809 8452
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8480 20775 8483
rect 20763 8452 21588 8480
rect 20763 8449 20775 8452
rect 20717 8443 20775 8449
rect 17957 8415 18015 8421
rect 17957 8412 17969 8415
rect 17736 8384 17969 8412
rect 17736 8372 17742 8384
rect 17957 8381 17969 8384
rect 18003 8381 18015 8415
rect 17957 8375 18015 8381
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8381 18199 8415
rect 20806 8412 20812 8424
rect 20767 8384 20812 8412
rect 18141 8375 18199 8381
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 21560 8421 21588 8452
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8412 21603 8415
rect 22278 8412 22284 8424
rect 21591 8384 22284 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 15197 8347 15255 8353
rect 15197 8313 15209 8347
rect 15243 8344 15255 8347
rect 17126 8344 17132 8356
rect 15243 8316 17132 8344
rect 15243 8313 15255 8316
rect 15197 8307 15255 8313
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 17368 8316 17509 8344
rect 17368 8304 17374 8316
rect 17497 8313 17509 8316
rect 17543 8313 17555 8347
rect 19886 8344 19892 8356
rect 19847 8316 19892 8344
rect 17497 8307 17555 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 20070 8304 20076 8356
rect 20128 8344 20134 8356
rect 20165 8347 20223 8353
rect 20165 8344 20177 8347
rect 20128 8316 20177 8344
rect 20128 8304 20134 8316
rect 20165 8313 20177 8316
rect 20211 8344 20223 8347
rect 21634 8344 21640 8356
rect 20211 8316 21640 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 21634 8304 21640 8316
rect 21692 8304 21698 8356
rect 14700 8248 14964 8276
rect 14700 8236 14706 8248
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15565 8279 15623 8285
rect 15565 8276 15577 8279
rect 15160 8248 15577 8276
rect 15160 8236 15166 8248
rect 15565 8245 15577 8248
rect 15611 8276 15623 8279
rect 15654 8276 15660 8288
rect 15611 8248 15660 8276
rect 15611 8245 15623 8248
rect 15565 8239 15623 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 18782 8276 18788 8288
rect 16264 8248 18788 8276
rect 16264 8236 16270 8248
rect 18782 8236 18788 8248
rect 18840 8236 18846 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19610 8276 19616 8288
rect 19484 8248 19616 8276
rect 19484 8236 19490 8248
rect 19610 8236 19616 8248
rect 19668 8276 19674 8288
rect 21085 8279 21143 8285
rect 21085 8276 21097 8279
rect 19668 8248 21097 8276
rect 19668 8236 19674 8248
rect 21085 8245 21097 8248
rect 21131 8276 21143 8279
rect 21269 8279 21327 8285
rect 21269 8276 21281 8279
rect 21131 8248 21281 8276
rect 21131 8245 21143 8248
rect 21085 8239 21143 8245
rect 21269 8245 21281 8248
rect 21315 8245 21327 8279
rect 21269 8239 21327 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2866 8072 2872 8084
rect 2827 8044 2872 8072
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6546 8072 6552 8084
rect 6420 8044 6552 8072
rect 6420 8032 6426 8044
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 6822 8072 6828 8084
rect 6779 8044 6828 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 3234 8004 3240 8016
rect 2240 7976 3240 8004
rect 2240 7948 2268 7976
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 6748 8004 6776 8035
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 6972 8044 7573 8072
rect 6972 8032 6978 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 7374 8004 7380 8016
rect 6328 7976 6776 8004
rect 6840 7976 7380 8004
rect 6328 7964 6334 7976
rect 2222 7936 2228 7948
rect 2135 7908 2228 7936
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 4154 7936 4160 7948
rect 3559 7908 4160 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4890 7936 4896 7948
rect 4851 7908 4896 7936
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 6840 7945 6868 7976
rect 7374 7964 7380 7976
rect 7432 7964 7438 8016
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3016 7840 3801 7868
rect 3016 7828 3022 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4430 7868 4436 7880
rect 4295 7840 4436 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4430 7828 4436 7840
rect 4488 7868 4494 7880
rect 4801 7871 4859 7877
rect 4488 7840 4568 7868
rect 4488 7828 4494 7840
rect 2317 7803 2375 7809
rect 2317 7769 2329 7803
rect 2363 7800 2375 7803
rect 3050 7800 3056 7812
rect 2363 7772 3056 7800
rect 2363 7769 2375 7772
rect 2317 7763 2375 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 3329 7803 3387 7809
rect 3329 7769 3341 7803
rect 3375 7800 3387 7803
rect 4540 7800 4568 7840
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 4982 7868 4988 7880
rect 4847 7840 4988 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5184 7800 5212 7831
rect 3375 7772 4384 7800
rect 4540 7772 5212 7800
rect 3375 7769 3387 7772
rect 3329 7763 3387 7769
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 1762 7732 1768 7744
rect 1719 7704 1768 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 2498 7732 2504 7744
rect 2455 7704 2504 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 3237 7735 3295 7741
rect 2832 7704 2877 7732
rect 2832 7692 2838 7704
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3602 7732 3608 7744
rect 3283 7704 3608 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 4356 7741 4384 7772
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7701 4399 7735
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4341 7695 4399 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5184 7732 5212 7772
rect 5350 7760 5356 7812
rect 5408 7809 5414 7812
rect 5408 7803 5472 7809
rect 5408 7769 5426 7803
rect 5460 7769 5472 7803
rect 5408 7763 5472 7769
rect 5408 7760 5414 7763
rect 5718 7760 5724 7812
rect 5776 7800 5782 7812
rect 6730 7800 6736 7812
rect 5776 7772 6736 7800
rect 5776 7760 5782 7772
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 6840 7732 6868 7899
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7282 7936 7288 7948
rect 6972 7908 7288 7936
rect 6972 7896 6978 7908
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7576 7800 7604 8035
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8352 8044 8953 8072
rect 8352 8032 8358 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 11425 8075 11483 8081
rect 8941 8035 8999 8041
rect 9048 8044 10824 8072
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 9048 8004 9076 8044
rect 10686 8004 10692 8016
rect 7800 7976 9076 8004
rect 9416 7976 10692 8004
rect 7800 7964 7806 7976
rect 9416 7948 9444 7976
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 10796 8004 10824 8044
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 12158 8072 12164 8084
rect 11471 8044 12164 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13817 8075 13875 8081
rect 13817 8072 13829 8075
rect 13504 8044 13829 8072
rect 13504 8032 13510 8044
rect 13817 8041 13829 8044
rect 13863 8072 13875 8075
rect 14734 8072 14740 8084
rect 13863 8044 14740 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 11698 8004 11704 8016
rect 10796 7976 11704 8004
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 8570 7936 8576 7948
rect 8531 7908 8576 7936
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9398 7936 9404 7948
rect 9359 7908 9404 7936
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9582 7936 9588 7948
rect 9543 7908 9588 7936
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9824 7908 9873 7936
rect 9824 7896 9830 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 9968 7908 10824 7936
rect 8386 7868 8392 7880
rect 8347 7840 8392 7868
rect 8386 7828 8392 7840
rect 8444 7828 8450 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 8536 7840 9321 7868
rect 8536 7828 8542 7840
rect 9309 7837 9321 7840
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9968 7800 9996 7908
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10594 7868 10600 7880
rect 10183 7840 10600 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 7576 7772 9996 7800
rect 10045 7803 10103 7809
rect 7006 7732 7012 7744
rect 5132 7704 6868 7732
rect 6967 7704 7012 7732
rect 5132 7692 5138 7704
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7190 7732 7196 7744
rect 7151 7704 7196 7732
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8202 7732 8208 7744
rect 8067 7704 8208 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8496 7741 8524 7772
rect 10045 7769 10057 7803
rect 10091 7800 10103 7803
rect 10796 7800 10824 7908
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 11020 7908 11161 7936
rect 11020 7896 11026 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 12894 7936 12900 7948
rect 11149 7899 11207 7905
rect 12728 7908 12900 7936
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11790 7868 11796 7880
rect 11103 7840 11796 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12549 7871 12607 7877
rect 12549 7837 12561 7871
rect 12595 7868 12607 7871
rect 12728 7868 12756 7908
rect 12894 7896 12900 7908
rect 12952 7936 12958 7948
rect 13449 7939 13507 7945
rect 13449 7936 13461 7939
rect 12952 7908 13461 7936
rect 12952 7896 12958 7908
rect 13449 7905 13461 7908
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 12595 7840 12756 7868
rect 12805 7871 12863 7877
rect 12595 7837 12607 7840
rect 12549 7831 12607 7837
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13832 7868 13860 8035
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 14884 8044 15240 8072
rect 14884 8032 14890 8044
rect 15212 8004 15240 8044
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 19061 8075 19119 8081
rect 16172 8044 18644 8072
rect 16172 8032 16178 8044
rect 17313 8007 17371 8013
rect 17313 8004 17325 8007
rect 15212 7976 17325 8004
rect 17313 7973 17325 7976
rect 17359 8004 17371 8007
rect 17678 8004 17684 8016
rect 17359 7976 17684 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17678 7964 17684 7976
rect 17736 7964 17742 8016
rect 18616 8004 18644 8044
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19518 8072 19524 8084
rect 19107 8044 19524 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19981 8075 20039 8081
rect 19981 8041 19993 8075
rect 20027 8072 20039 8075
rect 20254 8072 20260 8084
rect 20027 8044 20260 8072
rect 20027 8041 20039 8044
rect 19981 8035 20039 8041
rect 20254 8032 20260 8044
rect 20312 8032 20318 8084
rect 20809 8007 20867 8013
rect 20809 8004 20821 8007
rect 18616 7976 20821 8004
rect 20809 7973 20821 7976
rect 20855 7973 20867 8007
rect 20809 7967 20867 7973
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 16022 7936 16028 7948
rect 15712 7908 16028 7936
rect 15712 7896 15718 7908
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 13311 7840 13860 7868
rect 14093 7871 14151 7877
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 16132 7868 16160 7899
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 20438 7936 20444 7948
rect 16448 7908 17816 7936
rect 20399 7908 20444 7936
rect 16448 7896 16454 7908
rect 14093 7831 14151 7837
rect 15028 7840 16160 7868
rect 16669 7871 16727 7877
rect 12820 7800 12848 7831
rect 13722 7800 13728 7812
rect 10091 7772 10640 7800
rect 10796 7772 12434 7800
rect 12820 7772 13728 7800
rect 10091 7769 10103 7772
rect 10045 7763 10103 7769
rect 8481 7735 8539 7741
rect 8481 7701 8493 7735
rect 8527 7701 8539 7735
rect 8481 7695 8539 7701
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10318 7732 10324 7744
rect 9916 7704 10324 7732
rect 9916 7692 9922 7704
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10502 7732 10508 7744
rect 10463 7704 10508 7732
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10612 7741 10640 7772
rect 10597 7735 10655 7741
rect 10597 7701 10609 7735
rect 10643 7701 10655 7735
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10597 7695 10655 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12406 7732 12434 7772
rect 13722 7760 13728 7772
rect 13780 7800 13786 7812
rect 14108 7800 14136 7831
rect 15028 7812 15056 7840
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 16715 7840 17172 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 13780 7772 14136 7800
rect 14360 7803 14418 7809
rect 13780 7760 13786 7772
rect 14360 7769 14372 7803
rect 14406 7800 14418 7803
rect 15010 7800 15016 7812
rect 14406 7772 15016 7800
rect 14406 7769 14418 7772
rect 14360 7763 14418 7769
rect 15010 7760 15016 7772
rect 15068 7760 15074 7812
rect 16684 7800 16712 7831
rect 16408 7772 16712 7800
rect 17144 7800 17172 7840
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17368 7840 17693 7868
rect 17368 7828 17374 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17788 7868 17816 7908
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 20625 7939 20683 7945
rect 20625 7905 20637 7939
rect 20671 7936 20683 7939
rect 20714 7936 20720 7948
rect 20671 7908 20720 7936
rect 20671 7905 20683 7908
rect 20625 7899 20683 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 21358 7936 21364 7948
rect 21319 7908 21364 7936
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 18506 7868 18512 7880
rect 17788 7840 18512 7868
rect 17681 7831 17739 7837
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20898 7868 20904 7880
rect 20395 7840 20904 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21266 7868 21272 7880
rect 21192 7840 21272 7868
rect 17948 7803 18006 7809
rect 17144 7772 17356 7800
rect 12986 7732 12992 7744
rect 12406 7704 12992 7732
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 15470 7732 15476 7744
rect 13412 7704 13457 7732
rect 15431 7704 15476 7732
rect 13412 7692 13418 7704
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15562 7692 15568 7744
rect 15620 7732 15626 7744
rect 15620 7704 15665 7732
rect 15620 7692 15626 7704
rect 15838 7692 15844 7744
rect 15896 7732 15902 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15896 7704 15945 7732
rect 15896 7692 15902 7704
rect 15933 7701 15945 7704
rect 15979 7732 15991 7735
rect 16408 7732 16436 7772
rect 15979 7704 16436 7732
rect 16485 7735 16543 7741
rect 15979 7701 15991 7704
rect 15933 7695 15991 7701
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 16761 7735 16819 7741
rect 16761 7732 16773 7735
rect 16531 7704 16773 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 16761 7701 16773 7704
rect 16807 7732 16819 7735
rect 17218 7732 17224 7744
rect 16807 7704 17224 7732
rect 16807 7701 16819 7704
rect 16761 7695 16819 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17328 7732 17356 7772
rect 17948 7769 17960 7803
rect 17994 7800 18006 7803
rect 18874 7800 18880 7812
rect 17994 7772 18880 7800
rect 17994 7769 18006 7772
rect 17948 7763 18006 7769
rect 18874 7760 18880 7772
rect 18932 7760 18938 7812
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 21082 7800 21088 7812
rect 19751 7772 21088 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 18138 7732 18144 7744
rect 17328 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 19334 7732 19340 7744
rect 19295 7704 19340 7732
rect 19334 7692 19340 7704
rect 19392 7732 19398 7744
rect 19610 7732 19616 7744
rect 19392 7704 19616 7732
rect 19392 7692 19398 7704
rect 19610 7692 19616 7704
rect 19668 7692 19674 7744
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 21192 7741 21220 7840
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 21726 7800 21732 7812
rect 21416 7772 21732 7800
rect 21416 7760 21422 7772
rect 21726 7760 21732 7772
rect 21784 7760 21790 7812
rect 21177 7735 21235 7741
rect 21177 7732 21189 7735
rect 20956 7704 21189 7732
rect 20956 7692 20962 7704
rect 21177 7701 21189 7704
rect 21223 7701 21235 7735
rect 21177 7695 21235 7701
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 21634 7732 21640 7744
rect 21324 7704 21640 7732
rect 21324 7692 21330 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2832 7500 3157 7528
rect 2832 7488 2838 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3602 7528 3608 7540
rect 3563 7500 3608 7528
rect 3145 7491 3203 7497
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 4764 7500 5365 7528
rect 4764 7488 4770 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7497 7987 7531
rect 7929 7491 7987 7497
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 10226 7528 10232 7540
rect 9447 7500 9536 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 1949 7463 2007 7469
rect 1949 7460 1961 7463
rect 1544 7432 1961 7460
rect 1544 7420 1550 7432
rect 1949 7429 1961 7432
rect 1995 7460 2007 7463
rect 2130 7460 2136 7472
rect 1995 7432 2136 7460
rect 1995 7429 2007 7432
rect 1949 7423 2007 7429
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 2498 7460 2504 7472
rect 2459 7432 2504 7460
rect 2498 7420 2504 7432
rect 2556 7420 2562 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4430 7460 4436 7472
rect 4304 7432 4436 7460
rect 4304 7420 4310 7432
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4890 7420 4896 7472
rect 4948 7420 4954 7472
rect 4982 7420 4988 7472
rect 5040 7460 5046 7472
rect 5169 7463 5227 7469
rect 5169 7460 5181 7463
rect 5040 7432 5181 7460
rect 5040 7420 5046 7432
rect 5169 7429 5181 7432
rect 5215 7460 5227 7463
rect 5810 7460 5816 7472
rect 5215 7432 5816 7460
rect 5215 7429 5227 7432
rect 5169 7423 5227 7429
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 7374 7460 7380 7472
rect 6564 7432 7380 7460
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 1627 7364 2421 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2409 7361 2421 7364
rect 2455 7392 2467 7395
rect 2866 7392 2872 7404
rect 2455 7364 2872 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2866 7352 2872 7364
rect 2924 7352 2930 7404
rect 3234 7392 3240 7404
rect 3195 7364 3240 7392
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 4810 7395 4868 7401
rect 4810 7392 4822 7395
rect 4080 7364 4822 7392
rect 2590 7324 2596 7336
rect 2503 7296 2596 7324
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 2406 7216 2412 7268
rect 2464 7256 2470 7268
rect 2608 7256 2636 7284
rect 2464 7228 2636 7256
rect 2884 7256 2912 7352
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 4080 7324 4108 7364
rect 4810 7361 4822 7364
rect 4856 7392 4868 7395
rect 4908 7392 4936 7420
rect 5074 7392 5080 7404
rect 4856 7364 4936 7392
rect 5035 7364 5080 7392
rect 4856 7361 4868 7364
rect 4810 7355 4868 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 6564 7401 6592 7432
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 7944 7460 7972 7491
rect 8288 7463 8346 7469
rect 8288 7460 8300 7463
rect 7432 7432 7687 7460
rect 7944 7432 8300 7460
rect 7432 7420 7438 7432
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 6549 7395 6607 7401
rect 5767 7364 6500 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 3099 7296 4108 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 5960 7296 6005 7324
rect 5960 7284 5966 7296
rect 3418 7256 3424 7268
rect 2884 7228 3424 7256
rect 2464 7216 2470 7228
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 1762 7188 1768 7200
rect 1675 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7188 1826 7200
rect 2590 7188 2596 7200
rect 1820 7160 2596 7188
rect 1820 7148 1826 7160
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 3697 7191 3755 7197
rect 3697 7157 3709 7191
rect 3743 7188 3755 7191
rect 4154 7188 4160 7200
rect 3743 7160 4160 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 4154 7148 4160 7160
rect 4212 7188 4218 7200
rect 4798 7188 4804 7200
rect 4212 7160 4804 7188
rect 4212 7148 4218 7160
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6472 7197 6500 7364
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6816 7395 6874 7401
rect 6816 7361 6828 7395
rect 6862 7392 6874 7395
rect 7558 7392 7564 7404
rect 6862 7364 7564 7392
rect 6862 7361 6874 7364
rect 6816 7355 6874 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 7659 7392 7687 7432
rect 8288 7429 8300 7432
rect 8334 7460 8346 7463
rect 8570 7460 8576 7472
rect 8334 7432 8576 7460
rect 8334 7429 8346 7432
rect 8288 7423 8346 7429
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7659 7364 8033 7392
rect 8021 7361 8033 7364
rect 8067 7392 8079 7395
rect 8662 7392 8668 7404
rect 8067 7364 8668 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9398 7352 9404 7404
rect 9456 7392 9462 7404
rect 9508 7392 9536 7500
rect 10152 7500 10232 7528
rect 9858 7460 9864 7472
rect 9819 7432 9864 7460
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 9953 7463 10011 7469
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 10152 7460 10180 7500
rect 10226 7488 10232 7500
rect 10284 7528 10290 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 10284 7500 10517 7528
rect 10284 7488 10290 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10505 7491 10563 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11020 7500 11529 7528
rect 11020 7488 11026 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12308 7500 12357 7528
rect 12308 7488 12314 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 14737 7531 14795 7537
rect 12860 7500 14412 7528
rect 12860 7488 12866 7500
rect 10318 7460 10324 7472
rect 9999 7432 10180 7460
rect 10279 7432 10324 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 11146 7460 11152 7472
rect 10980 7432 11152 7460
rect 10980 7404 11008 7432
rect 11146 7420 11152 7432
rect 11204 7420 11210 7472
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 12713 7463 12771 7469
rect 12713 7460 12725 7463
rect 11296 7432 12725 7460
rect 11296 7420 11302 7432
rect 12713 7429 12725 7432
rect 12759 7460 12771 7463
rect 14384 7460 14412 7500
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15286 7528 15292 7540
rect 14783 7500 15292 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15473 7531 15531 7537
rect 15473 7497 15485 7531
rect 15519 7528 15531 7531
rect 15562 7528 15568 7540
rect 15519 7500 15568 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15654 7488 15660 7540
rect 15712 7528 15718 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15712 7500 16129 7528
rect 15712 7488 15718 7500
rect 16117 7497 16129 7500
rect 16163 7528 16175 7531
rect 16206 7528 16212 7540
rect 16163 7500 16212 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 17218 7488 17224 7540
rect 17276 7528 17282 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17276 7500 17693 7528
rect 17276 7488 17282 7500
rect 17681 7497 17693 7500
rect 17727 7528 17739 7531
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 17727 7500 18245 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 18233 7497 18245 7500
rect 18279 7528 18291 7531
rect 18598 7528 18604 7540
rect 18279 7500 18604 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 21174 7528 21180 7540
rect 20588 7500 20852 7528
rect 21135 7500 21180 7528
rect 20588 7488 20594 7500
rect 17954 7460 17960 7472
rect 12759 7432 14320 7460
rect 14384 7432 17960 7460
rect 12759 7429 12771 7432
rect 12713 7423 12771 7429
rect 9456 7364 10088 7392
rect 9456 7352 9462 7364
rect 10060 7333 10088 7364
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11882 7392 11888 7404
rect 11843 7364 11888 7392
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 14292 7401 14320 7432
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 19518 7460 19524 7472
rect 18892 7432 19524 7460
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 13044 7364 13277 7392
rect 13044 7352 13050 7364
rect 13265 7361 13277 7364
rect 13311 7392 13323 7395
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13311 7364 13829 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7392 14335 7395
rect 15102 7392 15108 7404
rect 14323 7364 15108 7392
rect 14323 7361 14335 7364
rect 14277 7355 14335 7361
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17494 7392 17500 7404
rect 17083 7364 17500 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 10045 7287 10103 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12802 7324 12808 7336
rect 12763 7296 12808 7324
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 12952 7296 13045 7324
rect 13096 7296 14105 7324
rect 12952 7284 12958 7296
rect 9122 7216 9128 7268
rect 9180 7256 9186 7268
rect 12526 7256 12532 7268
rect 9180 7228 12532 7256
rect 9180 7216 9186 7228
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12912 7256 12940 7284
rect 12676 7228 12940 7256
rect 12676 7216 12682 7228
rect 12986 7216 12992 7268
rect 13044 7256 13050 7268
rect 13096 7256 13124 7296
rect 14093 7293 14105 7296
rect 14139 7324 14151 7327
rect 14458 7324 14464 7336
rect 14139 7296 14464 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14826 7324 14832 7336
rect 14787 7296 14832 7324
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15010 7324 15016 7336
rect 14971 7296 15016 7324
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7324 15439 7327
rect 15470 7324 15476 7336
rect 15427 7296 15476 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7293 16819 7327
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16761 7287 16819 7293
rect 13044 7228 13124 7256
rect 13449 7259 13507 7265
rect 13044 7216 13050 7228
rect 13449 7225 13461 7259
rect 13495 7256 13507 7259
rect 14734 7256 14740 7268
rect 13495 7228 14740 7256
rect 13495 7225 13507 7228
rect 13449 7219 13507 7225
rect 14734 7216 14740 7228
rect 14792 7216 14798 7268
rect 16776 7256 16804 7287
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 17770 7324 17776 7336
rect 17328 7296 17776 7324
rect 17328 7256 17356 7296
rect 17770 7284 17776 7296
rect 17828 7324 17834 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17828 7296 17969 7324
rect 17828 7284 17834 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 18138 7324 18144 7336
rect 18099 7296 18144 7324
rect 17957 7287 18015 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18892 7333 18920 7432
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 20717 7463 20775 7469
rect 20717 7460 20729 7463
rect 19720 7432 20729 7460
rect 19058 7392 19064 7404
rect 19019 7364 19064 7392
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19720 7392 19748 7432
rect 20717 7429 20729 7432
rect 20763 7429 20775 7463
rect 20824 7460 20852 7500
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 21269 7463 21327 7469
rect 21269 7460 21281 7463
rect 20824 7432 21281 7460
rect 20717 7423 20775 7429
rect 21269 7429 21281 7432
rect 21315 7429 21327 7463
rect 21269 7423 21327 7429
rect 19886 7392 19892 7404
rect 19208 7364 19748 7392
rect 19847 7364 19892 7392
rect 19208 7352 19214 7364
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7392 20867 7395
rect 20898 7392 20904 7404
rect 20855 7364 20904 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 20898 7352 20904 7364
rect 20956 7392 20962 7404
rect 21082 7392 21088 7404
rect 20956 7364 21088 7392
rect 20956 7352 20962 7364
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 18877 7327 18935 7333
rect 18877 7293 18889 7327
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 18969 7327 19027 7333
rect 18969 7293 18981 7327
rect 19015 7324 19027 7327
rect 19981 7327 20039 7333
rect 19015 7296 19564 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19536 7265 19564 7296
rect 19981 7293 19993 7327
rect 20027 7293 20039 7327
rect 19981 7287 20039 7293
rect 16776 7228 17356 7256
rect 17405 7259 17463 7265
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 19521 7259 19579 7265
rect 17451 7228 18736 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 6457 7191 6515 7197
rect 6457 7157 6469 7191
rect 6503 7188 6515 7191
rect 6730 7188 6736 7200
rect 6503 7160 6736 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 10962 7188 10968 7200
rect 9548 7160 9593 7188
rect 10923 7160 10968 7188
rect 9548 7148 9554 7160
rect 10962 7148 10968 7160
rect 11020 7188 11026 7200
rect 11057 7191 11115 7197
rect 11057 7188 11069 7191
rect 11020 7160 11069 7188
rect 11020 7148 11026 7160
rect 11057 7157 11069 7160
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11882 7188 11888 7200
rect 11379 7160 11888 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 13170 7188 13176 7200
rect 12216 7160 13176 7188
rect 12216 7148 12222 7160
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13722 7188 13728 7200
rect 13683 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14366 7188 14372 7200
rect 14327 7160 14372 7188
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 17497 7191 17555 7197
rect 17497 7188 17509 7191
rect 17368 7160 17509 7188
rect 17368 7148 17374 7160
rect 17497 7157 17509 7160
rect 17543 7157 17555 7191
rect 18598 7188 18604 7200
rect 18559 7160 18604 7188
rect 17497 7151 17555 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18708 7188 18736 7228
rect 19521 7225 19533 7259
rect 19567 7225 19579 7259
rect 19521 7219 19579 7225
rect 19996 7188 20024 7287
rect 20070 7284 20076 7336
rect 20128 7324 20134 7336
rect 20625 7327 20683 7333
rect 20128 7296 20173 7324
rect 20128 7284 20134 7296
rect 20625 7293 20637 7327
rect 20671 7324 20683 7327
rect 20714 7324 20720 7336
rect 20671 7296 20720 7324
rect 20671 7293 20683 7296
rect 20625 7287 20683 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 21358 7216 21364 7268
rect 21416 7256 21422 7268
rect 21453 7259 21511 7265
rect 21453 7256 21465 7259
rect 21416 7228 21465 7256
rect 21416 7216 21422 7228
rect 21453 7225 21465 7228
rect 21499 7225 21511 7259
rect 21453 7219 21511 7225
rect 18708 7160 20024 7188
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2866 6984 2872 6996
rect 2280 6956 2872 6984
rect 2280 6944 2286 6956
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3786 6984 3792 6996
rect 3108 6956 3792 6984
rect 3108 6944 3114 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 9122 6984 9128 6996
rect 4120 6956 9128 6984
rect 4120 6944 4126 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 12032 6956 12081 6984
rect 12032 6944 12038 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 13909 6987 13967 6993
rect 13909 6984 13921 6987
rect 12584 6956 13921 6984
rect 12584 6944 12590 6956
rect 13909 6953 13921 6956
rect 13955 6984 13967 6987
rect 14826 6984 14832 6996
rect 13955 6956 14832 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15620 6956 15669 6984
rect 15620 6944 15626 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 18874 6984 18880 6996
rect 18835 6956 18880 6984
rect 15657 6947 15715 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 19058 6944 19064 6996
rect 19116 6984 19122 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 19116 6956 19257 6984
rect 19116 6944 19122 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 5902 6916 5908 6928
rect 4816 6888 5908 6916
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 3510 6808 3516 6860
rect 3568 6848 3574 6860
rect 3605 6851 3663 6857
rect 3605 6848 3617 6851
rect 3568 6820 3617 6848
rect 3568 6808 3574 6820
rect 3605 6817 3617 6820
rect 3651 6848 3663 6851
rect 3786 6848 3792 6860
rect 3651 6820 3792 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 4430 6780 4436 6792
rect 3283 6752 4436 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 4430 6740 4436 6752
rect 4488 6780 4494 6792
rect 4816 6780 4844 6888
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5258 6848 5264 6860
rect 5040 6820 5264 6848
rect 5040 6808 5046 6820
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5718 6848 5724 6860
rect 5679 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5828 6857 5856 6888
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 7190 6916 7196 6928
rect 6748 6888 7196 6916
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 6748 6848 6776 6888
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 9582 6916 9588 6928
rect 7616 6888 9588 6916
rect 7616 6876 7622 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 13630 6916 13636 6928
rect 11112 6888 13636 6916
rect 11112 6876 11118 6888
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 15286 6916 15292 6928
rect 13872 6888 15292 6916
rect 13872 6876 13878 6888
rect 15286 6876 15292 6888
rect 15344 6876 15350 6928
rect 18892 6916 18920 6944
rect 20070 6916 20076 6928
rect 18892 6888 20076 6916
rect 5813 6811 5871 6817
rect 5920 6820 6776 6848
rect 5350 6780 5356 6792
rect 4488 6752 4844 6780
rect 5000 6752 5356 6780
rect 4488 6740 4494 6752
rect 1756 6715 1814 6721
rect 1756 6681 1768 6715
rect 1802 6712 1814 6715
rect 2130 6712 2136 6724
rect 1802 6684 2136 6712
rect 1802 6681 1814 6684
rect 1756 6675 1814 6681
rect 2130 6672 2136 6684
rect 2188 6672 2194 6724
rect 3694 6712 3700 6724
rect 2884 6684 3700 6712
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2884 6653 2912 6684
rect 3694 6672 3700 6684
rect 3752 6712 3758 6724
rect 4045 6715 4103 6721
rect 4045 6712 4057 6715
rect 3752 6684 4057 6712
rect 3752 6672 3758 6684
rect 4045 6681 4057 6684
rect 4091 6681 4103 6715
rect 4045 6675 4103 6681
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2280 6616 2881 6644
rect 2280 6604 2286 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3329 6647 3387 6653
rect 3329 6644 3341 6647
rect 3108 6616 3341 6644
rect 3108 6604 3114 6616
rect 3329 6613 3341 6616
rect 3375 6613 3387 6647
rect 3329 6607 3387 6613
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5000 6644 5028 6752
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5920 6780 5948 6820
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6880 6820 6929 6848
rect 6880 6808 6886 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 7374 6848 7380 6860
rect 7287 6820 7380 6848
rect 6917 6811 6975 6817
rect 7374 6808 7380 6820
rect 7432 6848 7438 6860
rect 8113 6851 8171 6857
rect 8113 6848 8125 6851
rect 7432 6820 8125 6848
rect 7432 6808 7438 6820
rect 8113 6817 8125 6820
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 5644 6752 5948 6780
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5644 6721 5672 6752
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 7064 6752 7481 6780
rect 7064 6740 7070 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 7469 6743 7527 6749
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7742 6780 7748 6792
rect 7607 6752 7748 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8128 6780 8156 6811
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 8260 6820 8309 6848
rect 8260 6808 8266 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8938 6848 8944 6860
rect 8444 6820 8944 6848
rect 8444 6808 8450 6820
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9674 6848 9680 6860
rect 9180 6820 9680 6848
rect 9180 6808 9186 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 10962 6848 10968 6860
rect 10923 6820 10968 6848
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11698 6848 11704 6860
rect 11659 6820 11704 6848
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 12618 6848 12624 6860
rect 12579 6820 12624 6848
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 12986 6848 12992 6860
rect 12947 6820 12992 6848
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 14274 6848 14280 6860
rect 14187 6820 14280 6848
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 15010 6848 15016 6860
rect 14332 6820 14780 6848
rect 14971 6820 15016 6848
rect 14332 6808 14338 6820
rect 9398 6780 9404 6792
rect 8128 6752 9404 6780
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 12158 6780 12164 6792
rect 9646 6752 12164 6780
rect 5629 6715 5687 6721
rect 5629 6712 5641 6715
rect 5132 6684 5641 6712
rect 5132 6672 5138 6684
rect 5629 6681 5641 6684
rect 5675 6681 5687 6715
rect 5629 6675 5687 6681
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 5868 6684 6408 6712
rect 5868 6672 5874 6684
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 4764 6616 5181 6644
rect 4764 6604 4770 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 6270 6644 6276 6656
rect 5316 6616 5361 6644
rect 6231 6616 6276 6644
rect 5316 6604 5322 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6380 6653 6408 6684
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 6825 6715 6883 6721
rect 6825 6712 6837 6715
rect 6696 6684 6837 6712
rect 6696 6672 6702 6684
rect 6825 6681 6837 6684
rect 6871 6681 6883 6715
rect 6825 6675 6883 6681
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 9646 6712 9674 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13004 6780 13032 6808
rect 12575 6752 13032 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 14366 6740 14372 6792
rect 14424 6780 14430 6792
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14424 6752 14473 6780
rect 14424 6740 14430 6752
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14752 6780 14780 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15160 6820 15884 6848
rect 15160 6808 15166 6820
rect 15470 6780 15476 6792
rect 14752 6752 15476 6780
rect 14461 6743 14519 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 7248 6684 9674 6712
rect 7248 6672 7254 6684
rect 10410 6672 10416 6724
rect 10468 6712 10474 6724
rect 10698 6715 10756 6721
rect 10698 6712 10710 6715
rect 10468 6684 10710 6712
rect 10468 6672 10474 6684
rect 10698 6681 10710 6684
rect 10744 6681 10756 6715
rect 15289 6715 15347 6721
rect 15289 6712 15301 6715
rect 10698 6675 10756 6681
rect 10796 6684 15301 6712
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6613 6423 6647
rect 6365 6607 6423 6613
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6512 6616 6745 6644
rect 6512 6604 6518 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7616 6616 7941 6644
rect 7616 6604 7622 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 8352 6616 8401 6644
rect 8352 6604 8358 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8389 6607 8447 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9122 6644 9128 6656
rect 8904 6616 9128 6644
rect 8904 6604 8910 6616
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 10796 6644 10824 6684
rect 15289 6681 15301 6684
rect 15335 6712 15347 6715
rect 15749 6715 15807 6721
rect 15749 6712 15761 6715
rect 15335 6684 15761 6712
rect 15335 6681 15347 6684
rect 15289 6675 15347 6681
rect 15749 6681 15761 6684
rect 15795 6681 15807 6715
rect 15856 6712 15884 6820
rect 18598 6808 18604 6860
rect 18656 6848 18662 6860
rect 19812 6857 19840 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 18656 6820 19717 6848
rect 18656 6808 18662 6820
rect 19705 6817 19717 6820
rect 19751 6817 19763 6851
rect 19705 6811 19763 6817
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6817 19855 6851
rect 19797 6811 19855 6817
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 20404 6820 20637 6848
rect 20404 6808 20410 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 17126 6740 17132 6792
rect 17184 6789 17190 6792
rect 17184 6780 17196 6789
rect 17184 6752 17229 6780
rect 17184 6743 17196 6752
rect 17184 6740 17190 6743
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17770 6789 17776 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 17368 6752 17417 6780
rect 17368 6740 17374 6752
rect 17405 6749 17417 6752
rect 17451 6780 17463 6783
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17451 6752 17509 6780
rect 17451 6749 17463 6752
rect 17405 6743 17463 6749
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17764 6780 17776 6789
rect 17731 6752 17776 6780
rect 17497 6743 17555 6749
rect 17764 6743 17776 6752
rect 17770 6740 17776 6743
rect 17828 6740 17834 6792
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 20530 6780 20536 6792
rect 19484 6752 20536 6780
rect 19484 6740 19490 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20898 6780 20904 6792
rect 20859 6752 20904 6780
rect 20898 6740 20904 6752
rect 20956 6740 20962 6792
rect 17954 6712 17960 6724
rect 15856 6684 17960 6712
rect 15749 6675 15807 6681
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 20441 6715 20499 6721
rect 19659 6684 20116 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 11054 6644 11060 6656
rect 9456 6616 10824 6644
rect 11015 6616 11060 6644
rect 9456 6604 9462 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11296 6616 11437 6644
rect 11296 6604 11302 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 11517 6647 11575 6653
rect 11517 6613 11529 6647
rect 11563 6644 11575 6647
rect 11790 6644 11796 6656
rect 11563 6616 11796 6644
rect 11563 6613 11575 6616
rect 11517 6607 11575 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 11977 6647 12035 6653
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12437 6647 12495 6653
rect 12437 6644 12449 6647
rect 12023 6616 12449 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12437 6613 12449 6616
rect 12483 6644 12495 6647
rect 12710 6644 12716 6656
rect 12483 6616 12716 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 14366 6644 14372 6656
rect 14327 6616 14372 6644
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15197 6647 15255 6653
rect 15197 6613 15209 6647
rect 15243 6644 15255 6647
rect 15654 6644 15660 6656
rect 15243 6616 15660 6644
rect 15243 6613 15255 6616
rect 15197 6607 15255 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 16022 6644 16028 6656
rect 15983 6616 16028 6644
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 17034 6644 17040 6656
rect 16264 6616 17040 6644
rect 16264 6604 16270 6616
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 18874 6604 18880 6656
rect 18932 6644 18938 6656
rect 18969 6647 19027 6653
rect 18969 6644 18981 6647
rect 18932 6616 18981 6644
rect 18932 6604 18938 6616
rect 18969 6613 18981 6616
rect 19015 6644 19027 6647
rect 19518 6644 19524 6656
rect 19015 6616 19524 6644
rect 19015 6613 19027 6616
rect 18969 6607 19027 6613
rect 19518 6604 19524 6616
rect 19576 6644 19582 6656
rect 19702 6644 19708 6656
rect 19576 6616 19708 6644
rect 19576 6604 19582 6616
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 20088 6653 20116 6684
rect 20441 6681 20453 6715
rect 20487 6712 20499 6715
rect 21269 6715 21327 6721
rect 21269 6712 21281 6715
rect 20487 6684 21281 6712
rect 20487 6681 20499 6684
rect 20441 6675 20499 6681
rect 21269 6681 21281 6684
rect 21315 6681 21327 6715
rect 21269 6675 21327 6681
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 21085 6647 21143 6653
rect 21085 6613 21097 6647
rect 21131 6644 21143 6647
rect 21542 6644 21548 6656
rect 21131 6616 21548 6644
rect 21131 6613 21143 6616
rect 21085 6607 21143 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2958 6440 2964 6452
rect 2823 6412 2964 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3234 6440 3240 6452
rect 3191 6412 3240 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 3844 6412 6009 6440
rect 3844 6400 3850 6412
rect 5997 6409 6009 6412
rect 6043 6440 6055 6443
rect 7561 6443 7619 6449
rect 7561 6440 7573 6443
rect 6043 6412 7573 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 7561 6409 7573 6412
rect 7607 6440 7619 6443
rect 8110 6440 8116 6452
rect 7607 6412 8116 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8754 6440 8760 6452
rect 8343 6412 8760 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 8938 6440 8944 6452
rect 8899 6412 8944 6440
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9861 6443 9919 6449
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 9907 6412 10333 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 10735 6412 11529 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11974 6440 11980 6452
rect 11517 6403 11575 6409
rect 11624 6412 11980 6440
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3881 6375 3939 6381
rect 3881 6372 3893 6375
rect 3660 6344 3893 6372
rect 3660 6332 3666 6344
rect 3881 6341 3893 6344
rect 3927 6341 3939 6375
rect 3881 6335 3939 6341
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4430 6372 4436 6384
rect 4019 6344 4436 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 4522 6332 4528 6384
rect 4580 6381 4586 6384
rect 4580 6375 4644 6381
rect 4580 6341 4598 6375
rect 4632 6341 4644 6375
rect 4580 6335 4644 6341
rect 4580 6332 4586 6335
rect 6638 6332 6644 6384
rect 6696 6372 6702 6384
rect 6825 6375 6883 6381
rect 6825 6372 6837 6375
rect 6696 6344 6837 6372
rect 6696 6332 6702 6344
rect 6825 6341 6837 6344
rect 6871 6341 6883 6375
rect 6825 6335 6883 6341
rect 7469 6375 7527 6381
rect 7469 6341 7481 6375
rect 7515 6372 7527 6375
rect 7742 6372 7748 6384
rect 7515 6344 7748 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8389 6375 8447 6381
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 9490 6372 9496 6384
rect 8435 6344 9496 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 9490 6332 9496 6344
rect 9548 6332 9554 6384
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 11624 6372 11652 6412
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 13541 6443 13599 6449
rect 13541 6409 13553 6443
rect 13587 6440 13599 6443
rect 14366 6440 14372 6452
rect 13587 6412 14372 6440
rect 13587 6409 13599 6412
rect 13541 6403 13599 6409
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 15657 6443 15715 6449
rect 15657 6409 15669 6443
rect 15703 6440 15715 6443
rect 15930 6440 15936 6452
rect 15703 6412 15936 6440
rect 15703 6409 15715 6412
rect 15657 6403 15715 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17000 6412 17417 6440
rect 17000 6400 17006 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17405 6403 17463 6409
rect 17494 6400 17500 6452
rect 17552 6440 17558 6452
rect 17552 6412 17597 6440
rect 17552 6400 17558 6412
rect 17770 6400 17776 6452
rect 17828 6440 17834 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 17828 6412 18337 6440
rect 17828 6400 17834 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6440 19855 6443
rect 19886 6440 19892 6452
rect 19843 6412 19892 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 11885 6375 11943 6381
rect 11885 6372 11897 6375
rect 10100 6344 11652 6372
rect 11808 6344 11897 6372
rect 10100 6332 10106 6344
rect 2866 6304 2872 6316
rect 2608 6276 2872 6304
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6205 2099 6239
rect 2041 6199 2099 6205
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2406 6236 2412 6248
rect 2271 6208 2412 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2056 6168 2084 6199
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2608 6245 2636 6276
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2700 6168 2728 6199
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2832 6208 3249 6236
rect 2832 6196 2838 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3510 6196 3516 6248
rect 3568 6196 3574 6248
rect 3694 6196 3700 6248
rect 3752 6236 3758 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3752 6208 4077 6236
rect 3752 6196 3758 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 2056 6140 2728 6168
rect 3528 6168 3556 6196
rect 4246 6168 4252 6180
rect 3528 6140 4252 6168
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6100 1550 6112
rect 2056 6100 2084 6140
rect 4246 6128 4252 6140
rect 4304 6168 4310 6180
rect 4356 6168 4384 6267
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6604 6276 6745 6304
rect 6604 6264 6610 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 7650 6304 7656 6316
rect 6733 6267 6791 6273
rect 6840 6276 7656 6304
rect 6840 6236 6868 6276
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7760 6304 7788 6332
rect 11333 6307 11391 6313
rect 7760 6276 11284 6304
rect 4304 6140 4384 6168
rect 5552 6208 6868 6236
rect 4304 6128 4310 6140
rect 1544 6072 2084 6100
rect 1544 6060 1550 6072
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 3384 6072 3525 6100
rect 3384 6060 3390 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 3513 6063 3571 6069
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5552 6100 5580 6208
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7374 6236 7380 6248
rect 6972 6208 7017 6236
rect 7335 6208 7380 6236
rect 6972 6196 6978 6208
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 6178 6168 6184 6180
rect 6091 6140 6184 6168
rect 6178 6128 6184 6140
rect 6236 6168 6242 6180
rect 7760 6168 7788 6276
rect 8110 6236 8116 6248
rect 8071 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9766 6236 9772 6248
rect 9727 6208 9772 6236
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 10778 6236 10784 6248
rect 10739 6208 10784 6236
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10873 6239 10931 6245
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 11256 6236 11284 6276
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11808 6304 11836 6344
rect 11885 6341 11897 6344
rect 11931 6341 11943 6375
rect 11885 6335 11943 6341
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 13078 6372 13084 6384
rect 12216 6344 12434 6372
rect 13039 6344 13084 6372
rect 12216 6332 12222 6344
rect 12406 6304 12434 6344
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 14176 6375 14234 6381
rect 14176 6341 14188 6375
rect 14222 6372 14234 6375
rect 14274 6372 14280 6384
rect 14222 6344 14280 6372
rect 14222 6341 14234 6344
rect 14176 6335 14234 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 14826 6332 14832 6384
rect 14884 6372 14890 6384
rect 15749 6375 15807 6381
rect 15749 6372 15761 6375
rect 14884 6344 15761 6372
rect 14884 6332 14890 6344
rect 15749 6341 15761 6344
rect 15795 6341 15807 6375
rect 18340 6372 18368 6403
rect 19886 6400 19892 6412
rect 19944 6400 19950 6452
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20211 6412 20637 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 20346 6372 20352 6384
rect 18340 6344 20352 6372
rect 15749 6335 15807 6341
rect 20346 6332 20352 6344
rect 20404 6332 20410 6384
rect 20530 6332 20536 6384
rect 20588 6372 20594 6384
rect 21453 6375 21511 6381
rect 21453 6372 21465 6375
rect 20588 6344 21465 6372
rect 20588 6332 20594 6344
rect 21453 6341 21465 6344
rect 21499 6372 21511 6375
rect 22462 6372 22468 6384
rect 21499 6344 22468 6372
rect 21499 6341 21511 6344
rect 21453 6335 21511 6341
rect 22462 6332 22468 6344
rect 22520 6332 22526 6384
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 11379 6276 11836 6304
rect 11900 6276 12296 6304
rect 12406 6276 12541 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11900 6236 11928 6276
rect 11256 6208 11928 6236
rect 12069 6239 12127 6245
rect 10873 6199 10931 6205
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12268 6236 12296 6276
rect 12529 6273 12541 6276
rect 12575 6304 12587 6307
rect 13173 6307 13231 6313
rect 13173 6304 13185 6307
rect 12575 6276 13185 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 13173 6273 13185 6276
rect 13219 6273 13231 6307
rect 15010 6304 15016 6316
rect 13173 6267 13231 6273
rect 13832 6276 15016 6304
rect 12894 6236 12900 6248
rect 12268 6208 12900 6236
rect 12069 6199 12127 6205
rect 6236 6140 6776 6168
rect 6236 6128 6242 6140
rect 5718 6100 5724 6112
rect 4120 6072 5580 6100
rect 5679 6072 5724 6100
rect 4120 6060 4126 6072
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6362 6100 6368 6112
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6748 6100 6776 6140
rect 7300 6140 7788 6168
rect 9600 6140 10364 6168
rect 7300 6100 7328 6140
rect 9600 6112 9628 6140
rect 6748 6072 7328 6100
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7708 6072 7941 6100
rect 7708 6060 7714 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8570 6060 8576 6112
rect 8628 6100 8634 6112
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8628 6072 8769 6100
rect 8628 6060 8634 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 10100 6072 10241 6100
rect 10100 6060 10106 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10336 6100 10364 6140
rect 10410 6128 10416 6180
rect 10468 6168 10474 6180
rect 10888 6168 10916 6199
rect 10468 6140 10916 6168
rect 10468 6128 10474 6140
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 11606 6168 11612 6180
rect 11204 6140 11612 6168
rect 11204 6128 11210 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 11698 6100 11704 6112
rect 10336 6072 11704 6100
rect 10229 6063 10287 6069
rect 11698 6060 11704 6072
rect 11756 6100 11762 6112
rect 12084 6100 12112 6199
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6236 13047 6239
rect 13832 6236 13860 6276
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 16393 6307 16451 6313
rect 16393 6304 16405 6307
rect 15160 6276 16405 6304
rect 15160 6264 15166 6276
rect 16393 6273 16405 6276
rect 16439 6304 16451 6307
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16439 6276 17049 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17552 6276 17877 6304
rect 17552 6264 17558 6276
rect 17865 6273 17877 6276
rect 17911 6273 17923 6307
rect 19438 6307 19496 6313
rect 19438 6304 19450 6307
rect 17865 6267 17923 6273
rect 18064 6276 19450 6304
rect 13035 6208 13860 6236
rect 13909 6239 13967 6245
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 12621 6171 12679 6177
rect 12621 6168 12633 6171
rect 12216 6140 12633 6168
rect 12216 6128 12222 6140
rect 12621 6137 12633 6140
rect 12667 6168 12679 6171
rect 13078 6168 13084 6180
rect 12667 6140 13084 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13814 6128 13820 6180
rect 13872 6168 13878 6180
rect 13924 6168 13952 6199
rect 13872 6140 13952 6168
rect 15289 6171 15347 6177
rect 13872 6128 13878 6140
rect 15289 6137 15301 6171
rect 15335 6168 15347 6171
rect 15378 6168 15384 6180
rect 15335 6140 15384 6168
rect 15335 6137 15347 6140
rect 15289 6131 15347 6137
rect 15378 6128 15384 6140
rect 15436 6168 15442 6180
rect 15488 6168 15516 6199
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 15988 6208 16773 6236
rect 15988 6196 15994 6208
rect 16761 6205 16773 6208
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6236 17003 6239
rect 17402 6236 17408 6248
rect 16991 6208 17408 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 15436 6140 15516 6168
rect 15436 6128 15442 6140
rect 15746 6128 15752 6180
rect 15804 6168 15810 6180
rect 16209 6171 16267 6177
rect 16209 6168 16221 6171
rect 15804 6140 16221 6168
rect 15804 6128 15810 6140
rect 16209 6137 16221 6140
rect 16255 6137 16267 6171
rect 16776 6168 16804 6199
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18064 6245 18092 6276
rect 19438 6273 19450 6276
rect 19484 6304 19496 6307
rect 19886 6304 19892 6316
rect 19484 6276 19892 6304
rect 19484 6273 19496 6276
rect 19438 6267 19496 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17828 6208 17969 6236
rect 17828 6196 17834 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 19702 6236 19708 6248
rect 19663 6208 19708 6236
rect 18049 6199 18107 6205
rect 18064 6168 18092 6199
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 20254 6236 20260 6248
rect 20215 6208 20260 6236
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 20364 6245 20392 6332
rect 20806 6264 20812 6316
rect 20864 6304 20870 6316
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20864 6276 21005 6304
rect 20864 6264 20870 6276
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 21542 6304 21548 6316
rect 21140 6276 21548 6304
rect 21140 6264 21146 6276
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20349 6199 20407 6205
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 16776 6140 18092 6168
rect 16209 6131 16267 6137
rect 11756 6072 12112 6100
rect 11756 6060 11762 6072
rect 15838 6060 15844 6112
rect 15896 6100 15902 6112
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 15896 6072 16129 6100
rect 15896 6060 15902 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16224 6100 16252 6131
rect 19886 6128 19892 6180
rect 19944 6168 19950 6180
rect 21192 6168 21220 6199
rect 19944 6140 21220 6168
rect 19944 6128 19950 6140
rect 17310 6100 17316 6112
rect 16224 6072 17316 6100
rect 16117 6063 16175 6069
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17494 6060 17500 6112
rect 17552 6100 17558 6112
rect 21358 6100 21364 6112
rect 17552 6072 21364 6100
rect 17552 6060 17558 6072
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1857 5899 1915 5905
rect 1857 5896 1869 5899
rect 1452 5868 1869 5896
rect 1452 5856 1458 5868
rect 1857 5865 1869 5868
rect 1903 5865 1915 5899
rect 1857 5859 1915 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3142 5896 3148 5908
rect 2915 5868 3148 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 4709 5899 4767 5905
rect 4709 5896 4721 5899
rect 4488 5868 4721 5896
rect 4488 5856 4494 5868
rect 4709 5865 4721 5868
rect 4755 5865 4767 5899
rect 4709 5859 4767 5865
rect 5276 5868 6132 5896
rect 5276 5828 5304 5868
rect 5534 5828 5540 5840
rect 4448 5800 5304 5828
rect 5495 5800 5540 5828
rect 4448 5772 4476 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 2188 5732 2605 5760
rect 2188 5720 2194 5732
rect 2593 5729 2605 5732
rect 2639 5729 2651 5763
rect 3326 5760 3332 5772
rect 3287 5732 3332 5760
rect 2593 5723 2651 5729
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 2608 5692 2636 5723
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 4062 5760 4068 5772
rect 3559 5732 4068 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4430 5760 4436 5772
rect 4391 5732 4436 5760
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5261 5763 5319 5769
rect 5261 5760 5273 5763
rect 4908 5732 5273 5760
rect 4908 5692 4936 5732
rect 5261 5729 5273 5732
rect 5307 5760 5319 5763
rect 5718 5760 5724 5772
rect 5307 5732 5724 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 5994 5760 6000 5772
rect 5955 5732 6000 5760
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6104 5769 6132 5868
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 9122 5896 9128 5908
rect 6788 5868 9128 5896
rect 6788 5856 6794 5868
rect 9122 5856 9128 5868
rect 9180 5896 9186 5908
rect 10318 5896 10324 5908
rect 9180 5868 10324 5896
rect 9180 5856 9186 5868
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 11698 5896 11704 5908
rect 11480 5868 11704 5896
rect 11480 5856 11486 5868
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 12032 5868 12173 5896
rect 12032 5856 12038 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 13538 5896 13544 5908
rect 13499 5868 13544 5896
rect 12161 5859 12219 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 17034 5896 17040 5908
rect 13740 5868 17040 5896
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 13556 5828 13584 5856
rect 8720 5800 8984 5828
rect 8720 5788 8726 5800
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5760 6147 5763
rect 6914 5760 6920 5772
rect 6135 5732 6920 5760
rect 6135 5729 6147 5732
rect 6089 5723 6147 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7650 5760 7656 5772
rect 7611 5732 7656 5760
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 8110 5760 8116 5772
rect 7883 5732 8116 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8846 5760 8852 5772
rect 8251 5732 8852 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8956 5769 8984 5800
rect 10704 5800 12112 5828
rect 10704 5769 10732 5800
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 11977 5763 12035 5769
rect 11977 5729 11989 5763
rect 12023 5760 12035 5763
rect 12084 5760 12112 5800
rect 13188 5800 13584 5828
rect 13188 5769 13216 5800
rect 12023 5732 12112 5760
rect 13173 5763 13231 5769
rect 12023 5729 12035 5732
rect 11977 5723 12035 5729
rect 13173 5729 13185 5763
rect 13219 5729 13231 5763
rect 13173 5723 13231 5729
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13630 5760 13636 5772
rect 13403 5732 13636 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 2608 5664 4936 5692
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 6362 5692 6368 5704
rect 5123 5664 6368 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7282 5692 7288 5704
rect 6779 5664 7288 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7282 5652 7288 5664
rect 7340 5652 7346 5704
rect 7558 5692 7564 5704
rect 7519 5664 7564 5692
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 8352 5664 8401 5692
rect 8352 5652 8358 5664
rect 8389 5661 8401 5664
rect 8435 5692 8447 5695
rect 8478 5692 8484 5704
rect 8435 5664 8484 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9197 5695 9255 5701
rect 9197 5692 9209 5695
rect 8812 5664 9209 5692
rect 8812 5652 8818 5664
rect 9197 5661 9209 5664
rect 9243 5692 9255 5695
rect 9243 5664 9444 5692
rect 9243 5661 9255 5664
rect 9197 5655 9255 5661
rect 1578 5584 1584 5636
rect 1636 5624 1642 5636
rect 2409 5627 2467 5633
rect 2409 5624 2421 5627
rect 1636 5596 2421 5624
rect 1636 5584 1642 5596
rect 2409 5593 2421 5596
rect 2455 5593 2467 5627
rect 2409 5587 2467 5593
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 2547 5596 3832 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 3234 5556 3240 5568
rect 3195 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3804 5565 3832 5596
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 4706 5624 4712 5636
rect 4120 5596 4712 5624
rect 4120 5584 4126 5596
rect 4706 5584 4712 5596
rect 4764 5584 4770 5636
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 5215 5596 6408 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5525 3847 5559
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 3789 5519 3847 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4338 5556 4344 5568
rect 4295 5528 4344 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 6380 5565 6408 5596
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 9416 5624 9444 5664
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 10704 5692 10732 5723
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 10870 5692 10876 5704
rect 9548 5664 10732 5692
rect 10831 5664 10876 5692
rect 9548 5652 9554 5664
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11664 5664 11713 5692
rect 11664 5652 11670 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5661 11851 5695
rect 12158 5692 12164 5704
rect 11793 5655 11851 5661
rect 11992 5664 12164 5692
rect 9582 5624 9588 5636
rect 6604 5596 8892 5624
rect 9416 5596 9588 5624
rect 6604 5584 6610 5596
rect 5905 5559 5963 5565
rect 5905 5556 5917 5559
rect 5040 5528 5917 5556
rect 5040 5516 5046 5528
rect 5905 5525 5917 5528
rect 5951 5525 5963 5559
rect 5905 5519 5963 5525
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5525 6423 5559
rect 6822 5556 6828 5568
rect 6783 5528 6828 5556
rect 6365 5519 6423 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7190 5556 7196 5568
rect 7151 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8386 5556 8392 5568
rect 8343 5528 8392 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8536 5528 8769 5556
rect 8536 5516 8542 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8864 5556 8892 5596
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 10134 5584 10140 5636
rect 10192 5624 10198 5636
rect 10888 5624 10916 5652
rect 11146 5624 11152 5636
rect 10192 5596 10824 5624
rect 10888 5596 11152 5624
rect 10192 5584 10198 5596
rect 10152 5556 10180 5584
rect 8864 5528 10180 5556
rect 10321 5559 10379 5565
rect 8757 5519 8815 5525
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10410 5556 10416 5568
rect 10367 5528 10416 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 10796 5565 10824 5596
rect 11146 5584 11152 5596
rect 11204 5584 11210 5636
rect 11808 5624 11836 5655
rect 11992 5624 12020 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 12308 5664 12357 5692
rect 12308 5652 12314 5664
rect 12345 5661 12357 5664
rect 12391 5692 12403 5695
rect 13740 5692 13768 5868
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 19886 5856 19892 5908
rect 19944 5896 19950 5908
rect 19944 5868 20208 5896
rect 19944 5856 19950 5868
rect 16485 5831 16543 5837
rect 16485 5797 16497 5831
rect 16531 5828 16543 5831
rect 18138 5828 18144 5840
rect 16531 5800 18144 5828
rect 16531 5797 16543 5800
rect 16485 5791 16543 5797
rect 18138 5788 18144 5800
rect 18196 5788 18202 5840
rect 20180 5828 20208 5868
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20717 5899 20775 5905
rect 20717 5896 20729 5899
rect 20312 5868 20729 5896
rect 20312 5856 20318 5868
rect 20717 5865 20729 5868
rect 20763 5865 20775 5899
rect 20717 5859 20775 5865
rect 21082 5856 21088 5908
rect 21140 5896 21146 5908
rect 22094 5896 22100 5908
rect 21140 5868 22100 5896
rect 21140 5856 21146 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 20625 5831 20683 5837
rect 20625 5828 20637 5831
rect 20180 5800 20637 5828
rect 20625 5797 20637 5800
rect 20671 5828 20683 5831
rect 20671 5800 21312 5828
rect 20671 5797 20683 5800
rect 20625 5791 20683 5797
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16758 5760 16764 5772
rect 16719 5732 16764 5760
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 16960 5732 17877 5760
rect 12391 5664 13768 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 15378 5652 15384 5704
rect 15436 5701 15442 5704
rect 15436 5692 15448 5701
rect 15657 5695 15715 5701
rect 15436 5664 15481 5692
rect 15436 5655 15448 5664
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 15746 5692 15752 5704
rect 15703 5664 15752 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 15436 5652 15442 5655
rect 11808 5596 12020 5624
rect 12621 5627 12679 5633
rect 12621 5593 12633 5627
rect 12667 5624 12679 5627
rect 12802 5624 12808 5636
rect 12667 5596 12808 5624
rect 12667 5593 12679 5596
rect 12621 5587 12679 5593
rect 12802 5584 12808 5596
rect 12860 5624 12866 5636
rect 13081 5627 13139 5633
rect 13081 5624 13093 5627
rect 12860 5596 13093 5624
rect 12860 5584 12866 5596
rect 13081 5593 13093 5596
rect 13127 5593 13139 5627
rect 15672 5624 15700 5655
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 16114 5692 16120 5704
rect 16075 5664 16120 5692
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16960 5701 16988 5732
rect 17865 5729 17877 5732
rect 17911 5760 17923 5763
rect 18046 5760 18052 5772
rect 17911 5732 18052 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 18046 5720 18052 5732
rect 18104 5760 18110 5772
rect 21284 5769 21312 5800
rect 21269 5763 21327 5769
rect 18104 5732 19380 5760
rect 18104 5720 18110 5732
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 17402 5692 17408 5704
rect 17363 5664 17408 5692
rect 16945 5655 17003 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 17770 5692 17776 5704
rect 17727 5664 17776 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19352 5692 19380 5732
rect 21269 5729 21281 5763
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 22278 5692 22284 5704
rect 19352 5664 22284 5692
rect 19245 5655 19303 5661
rect 13081 5587 13139 5593
rect 15396 5596 15700 5624
rect 15396 5568 15424 5596
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 16853 5627 16911 5633
rect 16853 5624 16865 5627
rect 16632 5596 16865 5624
rect 16632 5584 16638 5596
rect 16853 5593 16865 5596
rect 16899 5593 16911 5627
rect 16853 5587 16911 5593
rect 17494 5584 17500 5636
rect 17552 5624 17558 5636
rect 18325 5627 18383 5633
rect 18325 5624 18337 5627
rect 17552 5596 18337 5624
rect 17552 5584 17558 5596
rect 18325 5593 18337 5596
rect 18371 5593 18383 5627
rect 18325 5587 18383 5593
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5525 10839 5559
rect 11238 5556 11244 5568
rect 11199 5528 11244 5556
rect 10781 5519 10839 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11333 5559 11391 5565
rect 11333 5525 11345 5559
rect 11379 5556 11391 5559
rect 11422 5556 11428 5568
rect 11379 5528 11428 5556
rect 11379 5525 11391 5528
rect 11333 5519 11391 5525
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 14274 5556 14280 5568
rect 12768 5528 12813 5556
rect 14235 5528 14280 5556
rect 12768 5516 12774 5528
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15378 5516 15384 5568
rect 15436 5516 15442 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 16025 5559 16083 5565
rect 16025 5556 16037 5559
rect 15620 5528 16037 5556
rect 15620 5516 15626 5528
rect 16025 5525 16037 5528
rect 16071 5525 16083 5559
rect 17310 5556 17316 5568
rect 17271 5528 17316 5556
rect 16025 5519 16083 5525
rect 17310 5516 17316 5528
rect 17368 5516 17374 5568
rect 18874 5516 18880 5568
rect 18932 5556 18938 5568
rect 18969 5559 19027 5565
rect 18969 5556 18981 5559
rect 18932 5528 18981 5556
rect 18932 5516 18938 5528
rect 18969 5525 18981 5528
rect 19015 5556 19027 5559
rect 19260 5556 19288 5655
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 19518 5633 19524 5636
rect 19512 5587 19524 5633
rect 19576 5624 19582 5636
rect 19576 5596 19612 5624
rect 19518 5584 19524 5587
rect 19576 5584 19582 5596
rect 21358 5584 21364 5636
rect 21416 5624 21422 5636
rect 22186 5624 22192 5636
rect 21416 5596 22192 5624
rect 21416 5584 21422 5596
rect 22186 5584 22192 5596
rect 22244 5584 22250 5636
rect 20070 5556 20076 5568
rect 19015 5528 20076 5556
rect 19015 5525 19027 5528
rect 18969 5519 19027 5525
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 21082 5556 21088 5568
rect 21043 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21266 5556 21272 5568
rect 21223 5528 21272 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21266 5516 21272 5528
rect 21324 5556 21330 5568
rect 21634 5556 21640 5568
rect 21324 5528 21640 5556
rect 21324 5516 21330 5528
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2317 5355 2375 5361
rect 2317 5352 2329 5355
rect 2096 5324 2329 5352
rect 2096 5312 2102 5324
rect 2317 5321 2329 5324
rect 2363 5321 2375 5355
rect 2317 5315 2375 5321
rect 2777 5355 2835 5361
rect 2777 5321 2789 5355
rect 2823 5352 2835 5355
rect 3234 5352 3240 5364
rect 2823 5324 3240 5352
rect 2823 5321 2835 5324
rect 2777 5315 2835 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4304 5324 4445 5352
rect 4304 5312 4310 5324
rect 4433 5321 4445 5324
rect 4479 5352 4491 5355
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4479 5324 5273 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 5261 5321 5273 5324
rect 5307 5321 5319 5355
rect 5261 5315 5319 5321
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5408 5324 5457 5352
rect 5408 5312 5414 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5905 5355 5963 5361
rect 5905 5352 5917 5355
rect 5592 5324 5917 5352
rect 5592 5312 5598 5324
rect 5905 5321 5917 5324
rect 5951 5321 5963 5355
rect 5905 5315 5963 5321
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7193 5355 7251 5361
rect 7193 5352 7205 5355
rect 6604 5324 7205 5352
rect 6604 5312 6610 5324
rect 7193 5321 7205 5324
rect 7239 5321 7251 5355
rect 7193 5315 7251 5321
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7340 5324 7389 5352
rect 7340 5312 7346 5324
rect 7377 5321 7389 5324
rect 7423 5352 7435 5355
rect 7834 5352 7840 5364
rect 7423 5324 7840 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8478 5352 8484 5364
rect 8343 5324 8484 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8588 5324 9536 5352
rect 1670 5284 1676 5296
rect 1631 5256 1676 5284
rect 1670 5244 1676 5256
rect 1728 5244 1734 5296
rect 1762 5244 1768 5296
rect 1820 5284 1826 5296
rect 2590 5284 2596 5296
rect 1820 5256 2596 5284
rect 1820 5244 1826 5256
rect 2590 5244 2596 5256
rect 2648 5284 2654 5296
rect 3114 5287 3172 5293
rect 3114 5284 3126 5287
rect 2648 5256 3126 5284
rect 2648 5244 2654 5256
rect 3114 5253 3126 5256
rect 3160 5253 3172 5287
rect 5074 5284 5080 5296
rect 5035 5256 5080 5284
rect 3114 5247 3172 5253
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 5810 5284 5816 5296
rect 5771 5256 5816 5284
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 7653 5287 7711 5293
rect 7653 5284 7665 5287
rect 7616 5256 7665 5284
rect 7616 5244 7622 5256
rect 7653 5253 7665 5256
rect 7699 5284 7711 5287
rect 8588 5284 8616 5324
rect 7699 5256 8616 5284
rect 7699 5253 7711 5256
rect 7653 5247 7711 5253
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 9094 5287 9152 5293
rect 9094 5284 9106 5287
rect 8904 5256 9106 5284
rect 8904 5244 8910 5256
rect 9094 5253 9106 5256
rect 9140 5284 9152 5287
rect 9508 5284 9536 5324
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 9640 5324 10241 5352
rect 9640 5312 9646 5324
rect 10229 5321 10241 5324
rect 10275 5352 10287 5355
rect 10318 5352 10324 5364
rect 10275 5324 10324 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 10778 5352 10784 5364
rect 10643 5324 10784 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 10870 5312 10876 5364
rect 10928 5352 10934 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10928 5324 10977 5352
rect 10928 5312 10934 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 10965 5315 11023 5321
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12710 5352 12716 5364
rect 12483 5324 12716 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 15562 5352 15568 5364
rect 15523 5324 15568 5352
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 16390 5352 16396 5364
rect 16351 5324 16396 5352
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17310 5352 17316 5364
rect 17083 5324 17316 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 19518 5352 19524 5364
rect 19479 5324 19524 5352
rect 19518 5312 19524 5324
rect 19576 5312 19582 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20864 5324 21005 5352
rect 20864 5312 20870 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 9140 5256 9444 5284
rect 9508 5256 9628 5284
rect 9140 5253 9152 5256
rect 9094 5247 9152 5253
rect 1946 5216 1952 5228
rect 1907 5188 1952 5216
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2406 5216 2412 5228
rect 2367 5188 2412 5216
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 4246 5216 4252 5228
rect 2915 5188 4252 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4982 5216 4988 5228
rect 4943 5188 4988 5216
rect 4982 5176 4988 5188
rect 5040 5216 5046 5228
rect 5166 5216 5172 5228
rect 5040 5188 5172 5216
rect 5040 5176 5046 5188
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 5592 5188 6745 5216
rect 5592 5176 5598 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 8386 5216 8392 5228
rect 8347 5188 8392 5216
rect 6733 5179 6791 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 8938 5216 8944 5228
rect 8720 5188 8944 5216
rect 8720 5176 8726 5188
rect 2222 5148 2228 5160
rect 2183 5120 2228 5148
rect 2222 5108 2228 5120
rect 2280 5108 2286 5160
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4801 5151 4859 5157
rect 4120 5120 4752 5148
rect 4120 5108 4126 5120
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 4430 5080 4436 5092
rect 4295 5052 4436 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 4430 5040 4436 5052
rect 4488 5040 4494 5092
rect 4724 5080 4752 5120
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 4890 5148 4896 5160
rect 4847 5120 4896 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5776 5120 6009 5148
rect 5776 5108 5782 5120
rect 5997 5117 6009 5120
rect 6043 5117 6055 5151
rect 5997 5111 6055 5117
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6604 5120 6837 5148
rect 6604 5108 6610 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 6972 5120 7021 5148
rect 6972 5108 6978 5120
rect 7009 5117 7021 5120
rect 7055 5148 7067 5151
rect 7282 5148 7288 5160
rect 7055 5120 7288 5148
rect 7055 5117 7067 5120
rect 7009 5111 7067 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8754 5148 8760 5160
rect 8251 5120 8760 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8864 5157 8892 5188
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9416 5216 9444 5256
rect 9490 5216 9496 5228
rect 9416 5188 9496 5216
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 9600 5216 9628 5256
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 10505 5287 10563 5293
rect 10505 5284 10517 5287
rect 9916 5256 10517 5284
rect 9916 5244 9922 5256
rect 10505 5253 10517 5256
rect 10551 5284 10563 5287
rect 10686 5284 10692 5296
rect 10551 5256 10692 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 13630 5244 13636 5296
rect 13688 5284 13694 5296
rect 14124 5287 14182 5293
rect 14124 5284 14136 5287
rect 13688 5256 14136 5284
rect 13688 5244 13694 5256
rect 14124 5253 14136 5256
rect 14170 5284 14182 5287
rect 16022 5284 16028 5296
rect 14170 5256 16028 5284
rect 14170 5253 14182 5256
rect 14124 5247 14182 5253
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 16114 5244 16120 5296
rect 16172 5244 16178 5296
rect 18874 5284 18880 5296
rect 18156 5256 18880 5284
rect 11057 5219 11115 5225
rect 9600 5188 10272 5216
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8662 5080 8668 5092
rect 4724 5052 8668 5080
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4396 4984 4537 5012
rect 4396 4972 4402 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 4525 4975 4583 4981
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 6052 4984 6377 5012
rect 6052 4972 6058 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6365 4975 6423 4981
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7708 4984 7849 5012
rect 7708 4972 7714 4984
rect 7837 4981 7849 4984
rect 7883 5012 7895 5015
rect 8294 5012 8300 5024
rect 7883 4984 8300 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8757 5015 8815 5021
rect 8757 4981 8769 5015
rect 8803 5012 8815 5015
rect 10134 5012 10140 5024
rect 8803 4984 10140 5012
rect 8803 4981 8815 4984
rect 8757 4975 8815 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10244 5012 10272 5188
rect 11057 5185 11069 5219
rect 11103 5216 11115 5219
rect 11698 5216 11704 5228
rect 11103 5188 11704 5216
rect 11103 5185 11115 5188
rect 11057 5179 11115 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12526 5216 12532 5228
rect 12487 5188 12532 5216
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 14826 5216 14832 5228
rect 14787 5188 14832 5216
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 15470 5216 15476 5228
rect 15383 5188 15476 5216
rect 15470 5176 15476 5188
rect 15528 5216 15534 5228
rect 16132 5216 16160 5244
rect 15528 5188 16160 5216
rect 15528 5176 15534 5188
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 18156 5225 18184 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 18966 5244 18972 5296
rect 19024 5284 19030 5296
rect 20717 5287 20775 5293
rect 19024 5256 20576 5284
rect 19024 5244 19030 5256
rect 18141 5219 18199 5225
rect 18141 5216 18153 5219
rect 17092 5188 18153 5216
rect 17092 5176 17098 5188
rect 18141 5185 18153 5188
rect 18187 5185 18199 5219
rect 18141 5179 18199 5185
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 18397 5219 18455 5225
rect 18397 5216 18409 5219
rect 18288 5188 18409 5216
rect 18288 5176 18294 5188
rect 18397 5185 18409 5188
rect 18443 5185 18455 5219
rect 18397 5179 18455 5185
rect 19610 5176 19616 5228
rect 19668 5216 19674 5228
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 19668 5188 19993 5216
rect 19668 5176 19674 5188
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 20441 5219 20499 5225
rect 20441 5216 20453 5219
rect 19981 5179 20039 5185
rect 20364 5188 20453 5216
rect 10318 5108 10324 5160
rect 10376 5148 10382 5160
rect 11195 5151 11253 5157
rect 11195 5148 11207 5151
rect 10376 5120 11207 5148
rect 10376 5108 10382 5120
rect 11195 5117 11207 5120
rect 11241 5117 11253 5151
rect 11195 5111 11253 5117
rect 11330 5108 11336 5160
rect 11388 5148 11394 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11388 5120 11529 5148
rect 11388 5108 11394 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 14369 5151 14427 5157
rect 12391 5120 12848 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12158 5080 12164 5092
rect 11716 5052 12164 5080
rect 10686 5012 10692 5024
rect 10244 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 11146 4972 11152 5024
rect 11204 5012 11210 5024
rect 11716 5021 11744 5052
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11204 4984 11713 5012
rect 11204 4972 11210 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11882 5012 11888 5024
rect 11843 4984 11888 5012
rect 11701 4975 11759 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12820 5012 12848 5120
rect 14369 5117 14381 5151
rect 14415 5148 14427 5151
rect 15378 5148 15384 5160
rect 14415 5120 15384 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 12943 5052 13492 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 12986 5012 12992 5024
rect 12820 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13464 5012 13492 5052
rect 14476 5024 14504 5120
rect 15378 5108 15384 5120
rect 15436 5148 15442 5160
rect 15749 5151 15807 5157
rect 15749 5148 15761 5151
rect 15436 5120 15761 5148
rect 15436 5108 15442 5120
rect 15749 5117 15761 5120
rect 15795 5148 15807 5151
rect 15930 5148 15936 5160
rect 15795 5120 15936 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 16114 5148 16120 5160
rect 16075 5120 16120 5148
rect 16114 5108 16120 5120
rect 16172 5148 16178 5160
rect 16390 5148 16396 5160
rect 16172 5120 16396 5148
rect 16172 5108 16178 5120
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16758 5148 16764 5160
rect 16719 5120 16764 5148
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16908 5120 16957 5148
rect 16908 5108 16914 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 16945 5111 17003 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 19705 5151 19763 5157
rect 19705 5148 19717 5151
rect 19576 5120 19717 5148
rect 19576 5108 19582 5120
rect 19705 5117 19717 5120
rect 19751 5117 19763 5151
rect 19886 5148 19892 5160
rect 19847 5120 19892 5148
rect 19705 5111 19763 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 16025 5083 16083 5089
rect 16025 5049 16037 5083
rect 16071 5080 16083 5083
rect 16206 5080 16212 5092
rect 16071 5052 16212 5080
rect 16071 5049 16083 5052
rect 16025 5043 16083 5049
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 20364 5089 20392 5188
rect 20441 5185 20453 5188
rect 20487 5185 20499 5219
rect 20548 5216 20576 5256
rect 20717 5253 20729 5287
rect 20763 5284 20775 5287
rect 20898 5284 20904 5296
rect 20763 5256 20904 5284
rect 20763 5253 20775 5256
rect 20717 5247 20775 5253
rect 20898 5244 20904 5256
rect 20956 5244 20962 5296
rect 21269 5219 21327 5225
rect 21269 5216 21281 5219
rect 20548 5188 21281 5216
rect 20441 5179 20499 5185
rect 21269 5185 21281 5188
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 17681 5083 17739 5089
rect 17681 5080 17693 5083
rect 16316 5052 17693 5080
rect 14366 5012 14372 5024
rect 13464 4984 14372 5012
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 14642 5012 14648 5024
rect 14516 4984 14561 5012
rect 14603 4984 14648 5012
rect 14516 4972 14522 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 14918 4972 14924 5024
rect 14976 5012 14982 5024
rect 16316 5012 16344 5052
rect 17681 5049 17693 5052
rect 17727 5049 17739 5083
rect 17681 5043 17739 5049
rect 20349 5083 20407 5089
rect 20349 5049 20361 5083
rect 20395 5049 20407 5083
rect 20349 5043 20407 5049
rect 17402 5012 17408 5024
rect 14976 4984 16344 5012
rect 17363 4984 17408 5012
rect 14976 4972 14982 4984
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 17696 5012 17724 5043
rect 18874 5012 18880 5024
rect 17696 4984 18880 5012
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 21542 5012 21548 5024
rect 21503 4984 21548 5012
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1762 4808 1768 4820
rect 1723 4780 1768 4808
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 2556 4780 3893 4808
rect 2556 4768 2562 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 4430 4808 4436 4820
rect 3881 4771 3939 4777
rect 4264 4780 4436 4808
rect 4264 4752 4292 4780
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4672 4780 5764 4808
rect 4672 4768 4678 4780
rect 3329 4743 3387 4749
rect 3329 4740 3341 4743
rect 3160 4712 3341 4740
rect 3160 4681 3188 4712
rect 3329 4709 3341 4712
rect 3375 4740 3387 4743
rect 4246 4740 4252 4752
rect 3375 4712 4252 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 5445 4743 5503 4749
rect 5445 4709 5457 4743
rect 5491 4740 5503 4743
rect 5626 4740 5632 4752
rect 5491 4712 5632 4740
rect 5491 4709 5503 4712
rect 5445 4703 5503 4709
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 5736 4740 5764 4780
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 6144 4780 6377 4808
rect 6144 4768 6150 4780
rect 6365 4777 6377 4780
rect 6411 4777 6423 4811
rect 6365 4771 6423 4777
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 8202 4808 8208 4820
rect 7156 4780 8208 4808
rect 7156 4768 7162 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8444 4780 8953 4808
rect 8444 4768 8450 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9824 4780 9873 4808
rect 9824 4768 9830 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 9861 4771 9919 4777
rect 10781 4811 10839 4817
rect 10781 4777 10793 4811
rect 10827 4808 10839 4811
rect 10962 4808 10968 4820
rect 10827 4780 10968 4808
rect 10827 4777 10839 4780
rect 10781 4771 10839 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11606 4808 11612 4820
rect 11296 4780 11612 4808
rect 11296 4768 11302 4780
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12526 4808 12532 4820
rect 12299 4780 12532 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 15654 4808 15660 4820
rect 13780 4780 15660 4808
rect 13780 4768 13786 4780
rect 15654 4768 15660 4780
rect 15712 4768 15718 4820
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16761 4811 16819 4817
rect 15988 4780 16712 4808
rect 15988 4768 15994 4780
rect 5736 4712 7420 4740
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4641 3203 4675
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 3145 4635 3203 4641
rect 3988 4644 4445 4672
rect 2958 4545 2964 4548
rect 2900 4539 2964 4545
rect 2900 4536 2912 4539
rect 2871 4508 2912 4536
rect 2900 4505 2912 4508
rect 2946 4505 2964 4539
rect 2900 4499 2964 4505
rect 2958 4496 2964 4499
rect 3016 4536 3022 4548
rect 3988 4536 4016 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 4433 4635 4491 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5994 4672 6000 4684
rect 5040 4644 5085 4672
rect 5955 4644 6000 4672
rect 5040 4632 5046 4644
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6144 4644 6189 4672
rect 6144 4632 6150 4644
rect 6932 4545 6960 4712
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7098 4672 7104 4684
rect 7055 4644 7104 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7282 4672 7288 4684
rect 7239 4644 7288 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7392 4672 7420 4712
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 8754 4740 8760 4752
rect 7524 4712 8432 4740
rect 8667 4712 8760 4740
rect 7524 4700 7530 4712
rect 8404 4684 8432 4712
rect 8754 4700 8760 4712
rect 8812 4740 8818 4752
rect 9398 4740 9404 4752
rect 8812 4712 9404 4740
rect 8812 4700 8818 4712
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 10686 4740 10692 4752
rect 9508 4712 10692 4740
rect 9508 4684 9536 4712
rect 10686 4700 10692 4712
rect 10744 4740 10750 4752
rect 10744 4712 11284 4740
rect 10744 4700 10750 4712
rect 7558 4672 7564 4684
rect 7392 4644 7564 4672
rect 7558 4632 7564 4644
rect 7616 4632 7622 4684
rect 7926 4632 7932 4684
rect 7984 4672 7990 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7984 4644 8033 4672
rect 7984 4632 7990 4644
rect 8021 4641 8033 4644
rect 8067 4672 8079 4675
rect 8110 4672 8116 4684
rect 8067 4644 8116 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 8444 4644 8493 4672
rect 8444 4632 8450 4644
rect 8481 4641 8493 4644
rect 8527 4672 8539 4675
rect 9490 4672 9496 4684
rect 8527 4644 9352 4672
rect 9451 4644 9496 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 9324 4613 9352 4644
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 10410 4672 10416 4684
rect 10371 4644 10416 4672
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 11256 4681 11284 4712
rect 12158 4700 12164 4752
rect 12216 4740 12222 4752
rect 14274 4740 14280 4752
rect 12216 4712 14280 4740
rect 12216 4700 12222 4712
rect 14274 4700 14280 4712
rect 14332 4700 14338 4752
rect 16684 4740 16712 4780
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 16850 4808 16856 4820
rect 16807 4780 16856 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17126 4768 17132 4820
rect 17184 4808 17190 4820
rect 17862 4808 17868 4820
rect 17184 4780 17868 4808
rect 17184 4768 17190 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 19760 4780 20361 4808
rect 19760 4768 19766 4780
rect 20349 4777 20361 4780
rect 20395 4808 20407 4811
rect 22554 4808 22560 4820
rect 20395 4780 22560 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 20070 4740 20076 4752
rect 14568 4712 16160 4740
rect 16684 4712 16896 4740
rect 20031 4712 20076 4740
rect 11241 4675 11299 4681
rect 10652 4644 11192 4672
rect 10652 4632 10658 4644
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9456 4576 9501 4604
rect 9456 4564 9462 4576
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10192 4576 10241 4604
rect 10192 4564 10198 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 11054 4604 11060 4616
rect 10367 4576 11060 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 11164 4604 11192 4644
rect 11241 4641 11253 4675
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11882 4672 11888 4684
rect 11664 4644 11888 4672
rect 11664 4632 11670 4644
rect 11882 4632 11888 4644
rect 11940 4672 11946 4684
rect 12897 4675 12955 4681
rect 11940 4644 12664 4672
rect 11940 4632 11946 4644
rect 11425 4607 11483 4613
rect 11425 4604 11437 4607
rect 11164 4576 11437 4604
rect 11425 4573 11437 4576
rect 11471 4604 11483 4607
rect 11698 4604 11704 4616
rect 11471 4576 11704 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 12636 4613 12664 4644
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 13630 4672 13636 4684
rect 12943 4644 13636 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 14568 4681 14596 4712
rect 16132 4684 16160 4712
rect 16868 4684 16896 4712
rect 20070 4700 20076 4712
rect 20128 4740 20134 4752
rect 20441 4743 20499 4749
rect 20441 4740 20453 4743
rect 20128 4712 20453 4740
rect 20128 4700 20134 4712
rect 20441 4709 20453 4712
rect 20487 4740 20499 4743
rect 20717 4743 20775 4749
rect 20717 4740 20729 4743
rect 20487 4712 20729 4740
rect 20487 4709 20499 4712
rect 20441 4703 20499 4709
rect 20717 4709 20729 4712
rect 20763 4709 20775 4743
rect 20717 4703 20775 4709
rect 14553 4675 14611 4681
rect 14553 4641 14565 4675
rect 14599 4641 14611 4675
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 14553 4635 14611 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4672 15899 4675
rect 16022 4672 16028 4684
rect 15887 4644 16028 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 16172 4644 16221 4672
rect 16172 4632 16178 4644
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 16666 4672 16672 4684
rect 16255 4644 16672 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 16908 4644 17001 4672
rect 16908 4632 16914 4644
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 18969 4675 19027 4681
rect 18969 4672 18981 4675
rect 17920 4644 18981 4672
rect 17920 4632 17926 4644
rect 18969 4641 18981 4644
rect 19015 4672 19027 4675
rect 19797 4675 19855 4681
rect 19797 4672 19809 4675
rect 19015 4644 19809 4672
rect 19015 4641 19027 4644
rect 18969 4635 19027 4641
rect 19797 4641 19809 4644
rect 19843 4641 19855 4675
rect 19797 4635 19855 4641
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 13262 4564 13268 4616
rect 13320 4604 13326 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13320 4576 13553 4604
rect 13320 4564 13326 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 3016 4508 4016 4536
rect 4341 4539 4399 4545
rect 3016 4496 3022 4508
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 5905 4539 5963 4545
rect 4387 4508 5580 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2740 4440 3433 4468
rect 2740 4428 2746 4440
rect 3421 4437 3433 4440
rect 3467 4468 3479 4471
rect 4062 4468 4068 4480
rect 3467 4440 4068 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5074 4468 5080 4480
rect 5035 4440 5080 4468
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5552 4477 5580 4508
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 6917 4539 6975 4545
rect 5951 4508 6592 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 6564 4477 6592 4508
rect 6917 4505 6929 4539
rect 6963 4505 6975 4539
rect 7852 4536 7880 4564
rect 7852 4508 8064 4536
rect 6917 4499 6975 4505
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4437 5595 4471
rect 5537 4431 5595 4437
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4437 6607 4471
rect 7374 4468 7380 4480
rect 7335 4440 7380 4468
rect 6549 4431 6607 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 7745 4471 7803 4477
rect 7745 4468 7757 4471
rect 7616 4440 7757 4468
rect 7616 4428 7622 4440
rect 7745 4437 7757 4440
rect 7791 4437 7803 4471
rect 7745 4431 7803 4437
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8036 4468 8064 4508
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 8754 4536 8760 4548
rect 8536 4508 8760 4536
rect 8536 4496 8542 4508
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 8904 4508 12081 4536
rect 8904 4496 8910 4508
rect 12069 4505 12081 4508
rect 12115 4536 12127 4539
rect 12434 4536 12440 4548
rect 12115 4508 12440 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 12434 4496 12440 4508
rect 12492 4536 12498 4548
rect 13449 4539 13507 4545
rect 13449 4536 13461 4539
rect 12492 4508 13461 4536
rect 12492 4496 12498 4508
rect 13449 4505 13461 4508
rect 13495 4505 13507 4539
rect 13556 4536 13584 4567
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14642 4604 14648 4616
rect 13780 4576 14648 4604
rect 13780 4564 13786 4576
rect 14642 4564 14648 4576
rect 14700 4604 14706 4616
rect 14737 4607 14795 4613
rect 14737 4604 14749 4607
rect 14700 4576 14749 4604
rect 14700 4564 14706 4576
rect 14737 4573 14749 4576
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 15565 4607 15623 4613
rect 15565 4573 15577 4607
rect 15611 4604 15623 4607
rect 15746 4604 15752 4616
rect 15611 4576 15752 4604
rect 15611 4573 15623 4576
rect 15565 4567 15623 4573
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 16390 4604 16396 4616
rect 16351 4576 16396 4604
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16960 4576 17264 4604
rect 14093 4539 14151 4545
rect 14093 4536 14105 4539
rect 13556 4508 14105 4536
rect 13449 4499 13507 4505
rect 14093 4505 14105 4508
rect 14139 4505 14151 4539
rect 16960 4536 16988 4576
rect 14093 4499 14151 4505
rect 15120 4508 16988 4536
rect 17120 4539 17178 4545
rect 10410 4468 10416 4480
rect 7892 4440 7937 4468
rect 8036 4440 10416 4468
rect 7892 4428 7898 4440
rect 10410 4428 10416 4440
rect 10468 4468 10474 4480
rect 10594 4468 10600 4480
rect 10468 4440 10600 4468
rect 10468 4428 10474 4440
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 10870 4468 10876 4480
rect 10831 4440 10876 4468
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11333 4471 11391 4477
rect 11333 4468 11345 4471
rect 11112 4440 11345 4468
rect 11112 4428 11118 4440
rect 11333 4437 11345 4440
rect 11379 4437 11391 4471
rect 11974 4468 11980 4480
rect 11887 4440 11980 4468
rect 11333 4431 11391 4437
rect 11974 4428 11980 4440
rect 12032 4468 12038 4480
rect 12526 4468 12532 4480
rect 12032 4440 12532 4468
rect 12032 4428 12038 4440
rect 12526 4428 12532 4440
rect 12584 4468 12590 4480
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 12584 4440 12725 4468
rect 12584 4428 12590 4440
rect 12713 4437 12725 4440
rect 12759 4437 12771 4471
rect 13078 4468 13084 4480
rect 13039 4440 13084 4468
rect 12713 4431 12771 4437
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 14642 4468 14648 4480
rect 14555 4440 14648 4468
rect 14642 4428 14648 4440
rect 14700 4468 14706 4480
rect 14826 4468 14832 4480
rect 14700 4440 14832 4468
rect 14700 4428 14706 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15120 4477 15148 4508
rect 17120 4505 17132 4539
rect 17166 4505 17178 4539
rect 17236 4536 17264 4576
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 18104 4576 19625 4604
rect 18104 4564 18110 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 22370 4604 22376 4616
rect 19613 4567 19671 4573
rect 19720 4576 22376 4604
rect 18785 4539 18843 4545
rect 18785 4536 18797 4539
rect 17236 4508 18797 4536
rect 17120 4499 17178 4505
rect 18785 4505 18797 4508
rect 18831 4505 18843 4539
rect 19720 4536 19748 4576
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 18785 4499 18843 4505
rect 18892 4508 19748 4536
rect 21361 4539 21419 4545
rect 15105 4471 15163 4477
rect 15105 4437 15117 4471
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15252 4440 15297 4468
rect 15252 4428 15258 4440
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 16264 4440 16313 4468
rect 16264 4428 16270 4440
rect 16301 4437 16313 4440
rect 16347 4437 16359 4471
rect 16301 4431 16359 4437
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 16942 4468 16948 4480
rect 16816 4440 16948 4468
rect 16816 4428 16822 4440
rect 16942 4428 16948 4440
rect 17000 4468 17006 4480
rect 17144 4468 17172 4499
rect 18892 4480 18920 4508
rect 21361 4505 21373 4539
rect 21407 4536 21419 4539
rect 21634 4536 21640 4548
rect 21407 4508 21640 4536
rect 21407 4505 21419 4508
rect 21361 4499 21419 4505
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 17862 4468 17868 4480
rect 17000 4440 17868 4468
rect 17000 4428 17006 4440
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 18693 4471 18751 4477
rect 18380 4440 18425 4468
rect 18380 4428 18386 4440
rect 18693 4437 18705 4471
rect 18739 4468 18751 4471
rect 18874 4468 18880 4480
rect 18739 4440 18880 4468
rect 18739 4437 18751 4440
rect 18693 4431 18751 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19242 4468 19248 4480
rect 19203 4440 19248 4468
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 19702 4468 19708 4480
rect 19663 4440 19708 4468
rect 19702 4428 19708 4440
rect 19760 4428 19766 4480
rect 21174 4468 21180 4480
rect 21135 4440 21180 4468
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 21542 4468 21548 4480
rect 21503 4440 21548 4468
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2464 4236 2697 4264
rect 2464 4224 2470 4236
rect 2685 4233 2697 4236
rect 2731 4233 2743 4267
rect 2958 4264 2964 4276
rect 2919 4236 2964 4264
rect 2685 4227 2743 4233
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5997 4267 6055 4273
rect 5997 4264 6009 4267
rect 5592 4236 6009 4264
rect 5592 4224 5598 4236
rect 5997 4233 6009 4236
rect 6043 4264 6055 4267
rect 6546 4264 6552 4276
rect 6043 4236 6552 4264
rect 6043 4233 6055 4236
rect 5997 4227 6055 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 6914 4224 6920 4276
rect 6972 4224 6978 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 8570 4264 8576 4276
rect 7340 4236 8064 4264
rect 8531 4236 8576 4264
rect 7340 4224 7346 4236
rect 2317 4199 2375 4205
rect 2317 4165 2329 4199
rect 2363 4196 2375 4199
rect 2774 4196 2780 4208
rect 2363 4168 2780 4196
rect 2363 4165 2375 4168
rect 2317 4159 2375 4165
rect 2774 4156 2780 4168
rect 2832 4156 2838 4208
rect 4890 4156 4896 4208
rect 4948 4196 4954 4208
rect 5660 4199 5718 4205
rect 5660 4196 5672 4199
rect 4948 4168 5672 4196
rect 4948 4156 4954 4168
rect 5660 4165 5672 4168
rect 5706 4196 5718 4199
rect 6932 4196 6960 4224
rect 5706 4168 6960 4196
rect 7092 4199 7150 4205
rect 5706 4165 5718 4168
rect 5660 4159 5718 4165
rect 7092 4165 7104 4199
rect 7138 4196 7150 4199
rect 7926 4196 7932 4208
rect 7138 4168 7932 4196
rect 7138 4165 7150 4168
rect 7092 4159 7150 4165
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8036 4196 8064 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 9122 4264 9128 4276
rect 8720 4236 8892 4264
rect 9083 4236 9128 4264
rect 8720 4224 8726 4236
rect 8864 4196 8892 4236
rect 9122 4224 9128 4236
rect 9180 4264 9186 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9180 4236 9781 4264
rect 9180 4224 9186 4236
rect 9769 4233 9781 4236
rect 9815 4264 9827 4267
rect 11606 4264 11612 4276
rect 9815 4236 11612 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12250 4264 12256 4276
rect 12032 4236 12256 4264
rect 12032 4224 12038 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 13078 4264 13084 4276
rect 13039 4236 13084 4264
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 14645 4267 14703 4273
rect 13740 4236 14596 4264
rect 9674 4196 9680 4208
rect 8036 4168 8800 4196
rect 8864 4168 9680 4196
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3326 4128 3332 4140
rect 2915 4100 3332 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4085 4131 4143 4137
rect 4085 4097 4097 4131
rect 4131 4128 4143 4131
rect 4131 4100 4568 4128
rect 4131 4097 4143 4100
rect 4085 4091 4143 4097
rect 2130 4060 2136 4072
rect 2091 4032 2136 4060
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 4430 4060 4436 4072
rect 4387 4032 4436 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 1762 3924 1768 3936
rect 1544 3896 1768 3924
rect 1544 3884 1550 3896
rect 1762 3884 1768 3896
rect 1820 3924 1826 3936
rect 2240 3924 2268 4023
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4540 3936 4568 4100
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 5905 4131 5963 4137
rect 5132 4100 5856 4128
rect 5132 4088 5138 4100
rect 5828 4060 5856 4100
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6178 4128 6184 4140
rect 5951 4100 6184 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6178 4088 6184 4100
rect 6236 4128 6242 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6236 4100 6837 4128
rect 6236 4088 6242 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8662 4128 8668 4140
rect 6972 4100 8524 4128
rect 8623 4100 8668 4128
rect 6972 4088 6978 4100
rect 6086 4060 6092 4072
rect 5828 4032 6092 4060
rect 6086 4020 6092 4032
rect 6144 4060 6150 4072
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 6144 4032 6561 4060
rect 6144 4020 6150 4032
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 6549 4023 6607 4029
rect 8220 4032 8401 4060
rect 6457 3995 6515 4001
rect 6457 3961 6469 3995
rect 6503 3992 6515 3995
rect 6638 3992 6644 4004
rect 6503 3964 6644 3992
rect 6503 3961 6515 3964
rect 6457 3955 6515 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 4522 3924 4528 3936
rect 1820 3896 2268 3924
rect 4435 3896 4528 3924
rect 1820 3884 1826 3896
rect 4522 3884 4528 3896
rect 4580 3924 4586 3936
rect 5994 3924 6000 3936
rect 4580 3896 6000 3924
rect 4580 3884 4586 3896
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 8220 3933 8248 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7156 3896 8217 3924
rect 7156 3884 7162 3896
rect 8205 3893 8217 3896
rect 8251 3924 8263 3927
rect 8294 3924 8300 3936
rect 8251 3896 8300 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8496 3924 8524 4100
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 8772 4060 8800 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 9953 4199 10011 4205
rect 9953 4165 9965 4199
rect 9999 4196 10011 4199
rect 10965 4199 11023 4205
rect 10965 4196 10977 4199
rect 9999 4168 10977 4196
rect 9999 4165 10011 4168
rect 9953 4159 10011 4165
rect 10965 4165 10977 4168
rect 11011 4196 11023 4199
rect 11011 4168 11100 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9088 4100 9321 4128
rect 9088 4088 9094 4100
rect 9309 4097 9321 4100
rect 9355 4128 9367 4131
rect 9582 4128 9588 4140
rect 9355 4100 9588 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10042 4128 10048 4140
rect 10003 4100 10048 4128
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 10870 4128 10876 4140
rect 10244 4100 10876 4128
rect 9600 4060 9628 4088
rect 10244 4060 10272 4100
rect 10870 4088 10876 4100
rect 10928 4128 10934 4140
rect 11072 4128 11100 4168
rect 11330 4128 11336 4140
rect 10928 4100 11008 4128
rect 11072 4100 11336 4128
rect 10928 4088 10934 4100
rect 8772 4032 9352 4060
rect 9600 4032 10272 4060
rect 10321 4063 10379 4069
rect 9033 3995 9091 4001
rect 9033 3961 9045 3995
rect 9079 3992 9091 3995
rect 9214 3992 9220 4004
rect 9079 3964 9220 3992
rect 9079 3961 9091 3964
rect 9033 3955 9091 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9324 3992 9352 4032
rect 10321 4029 10333 4063
rect 10367 4060 10379 4063
rect 10980 4060 11008 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 12158 4128 12164 4140
rect 11440 4100 12164 4128
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 10367 4032 10916 4060
rect 10980 4032 11069 4060
rect 10367 4029 10379 4032
rect 10321 4023 10379 4029
rect 10888 3992 10916 4032
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11440 4060 11468 4100
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12342 4128 12348 4140
rect 12303 4100 12348 4128
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12492 4100 13185 4128
rect 12492 4088 12498 4100
rect 13173 4097 13185 4100
rect 13219 4128 13231 4131
rect 13740 4128 13768 4236
rect 14458 4156 14464 4208
rect 14516 4156 14522 4208
rect 14568 4196 14596 4236
rect 14645 4233 14657 4267
rect 14691 4264 14703 4267
rect 15194 4264 15200 4276
rect 14691 4236 15200 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 15194 4224 15200 4236
rect 15252 4224 15258 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 17126 4264 17132 4276
rect 15804 4236 17132 4264
rect 15804 4224 15810 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17402 4224 17408 4276
rect 17460 4264 17466 4276
rect 17589 4267 17647 4273
rect 17589 4264 17601 4267
rect 17460 4236 17601 4264
rect 17460 4224 17466 4236
rect 17589 4233 17601 4236
rect 17635 4233 17647 4267
rect 17589 4227 17647 4233
rect 18322 4224 18328 4276
rect 18380 4264 18386 4276
rect 18417 4267 18475 4273
rect 18417 4264 18429 4267
rect 18380 4236 18429 4264
rect 18380 4224 18386 4236
rect 18417 4233 18429 4236
rect 18463 4233 18475 4267
rect 18417 4227 18475 4233
rect 18509 4267 18567 4273
rect 18509 4233 18521 4267
rect 18555 4264 18567 4267
rect 19242 4264 19248 4276
rect 18555 4236 19248 4264
rect 18555 4233 18567 4236
rect 18509 4227 18567 4233
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 20070 4264 20076 4276
rect 19383 4236 20076 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 20070 4224 20076 4236
rect 20128 4264 20134 4276
rect 22094 4264 22100 4276
rect 20128 4236 22100 4264
rect 20128 4224 20134 4236
rect 22094 4224 22100 4236
rect 22152 4224 22158 4276
rect 14918 4196 14924 4208
rect 14568 4168 14924 4196
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 15654 4156 15660 4208
rect 15712 4196 15718 4208
rect 16853 4199 16911 4205
rect 16853 4196 16865 4199
rect 15712 4168 16865 4196
rect 15712 4156 15718 4168
rect 16853 4165 16865 4168
rect 16899 4196 16911 4199
rect 17218 4196 17224 4208
rect 16899 4168 17224 4196
rect 16899 4165 16911 4168
rect 16853 4159 16911 4165
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 19886 4196 19892 4208
rect 19260 4168 19892 4196
rect 13219 4100 13768 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14476 4128 14504 4156
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 13872 4100 15117 4128
rect 13872 4088 13878 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15372 4131 15430 4137
rect 15372 4097 15384 4131
rect 15418 4128 15430 4131
rect 16114 4128 16120 4140
rect 15418 4100 16120 4128
rect 15418 4097 15430 4100
rect 15372 4091 15430 4097
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 17034 4088 17040 4140
rect 17092 4128 17098 4140
rect 17678 4128 17684 4140
rect 17092 4100 17137 4128
rect 17639 4100 17684 4128
rect 17092 4088 17098 4100
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 11606 4060 11612 4072
rect 11287 4032 11468 4060
rect 11567 4032 11612 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 10962 3992 10968 4004
rect 9324 3964 10824 3992
rect 10888 3964 10968 3992
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 8496 3896 9505 3924
rect 9493 3893 9505 3896
rect 9539 3924 9551 3927
rect 10318 3924 10324 3936
rect 9539 3896 10324 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 10594 3924 10600 3936
rect 10555 3896 10600 3924
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 10796 3924 10824 3964
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 11256 3924 11284 4023
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12250 4060 12256 4072
rect 12211 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12986 4060 12992 4072
rect 12899 4032 12992 4060
rect 12986 4020 12992 4032
rect 13044 4060 13050 4072
rect 13722 4060 13728 4072
rect 13044 4032 13728 4060
rect 13044 4020 13050 4032
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14458 4060 14464 4072
rect 14231 4032 14464 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 14550 4020 14556 4072
rect 14608 4020 14614 4072
rect 14734 4060 14740 4072
rect 14695 4032 14740 4060
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 14918 4060 14924 4072
rect 14879 4032 14924 4060
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 16761 4063 16819 4069
rect 16761 4029 16773 4063
rect 16807 4060 16819 4063
rect 17126 4060 17132 4072
rect 16807 4032 17132 4060
rect 16807 4029 16819 4032
rect 16761 4023 16819 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17497 4063 17555 4069
rect 17497 4029 17509 4063
rect 17543 4060 17555 4063
rect 18230 4060 18236 4072
rect 17543 4032 18236 4060
rect 17543 4029 17555 4032
rect 17497 4023 17555 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 19260 4060 19288 4168
rect 19886 4156 19892 4168
rect 19944 4156 19950 4208
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 19794 4128 19800 4140
rect 19475 4100 19800 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 19794 4088 19800 4100
rect 19852 4128 19858 4140
rect 19852 4100 19932 4128
rect 19852 4088 19858 4100
rect 19518 4060 19524 4072
rect 18800 4032 19288 4060
rect 19479 4032 19524 4060
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 12158 3992 12164 4004
rect 11480 3964 12164 3992
rect 11480 3952 11486 3964
rect 12158 3952 12164 3964
rect 12216 3992 12222 4004
rect 14568 3992 14596 4020
rect 12216 3964 14596 3992
rect 16485 3995 16543 4001
rect 12216 3952 12222 3964
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 16850 3992 16856 4004
rect 16531 3964 16856 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 17954 3992 17960 4004
rect 16960 3964 17960 3992
rect 10796 3896 11284 3924
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11572 3896 11805 3924
rect 11572 3884 11578 3896
rect 11793 3893 11805 3896
rect 11839 3924 11851 3927
rect 12434 3924 12440 3936
rect 11839 3896 12440 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 12894 3924 12900 3936
rect 12759 3896 12900 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13538 3924 13544 3936
rect 13499 3896 13544 3924
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 13814 3924 13820 3936
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14277 3927 14335 3933
rect 14277 3893 14289 3927
rect 14323 3924 14335 3927
rect 14550 3924 14556 3936
rect 14323 3896 14556 3924
rect 14323 3893 14335 3896
rect 14277 3887 14335 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 16960 3924 16988 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 18049 3995 18107 4001
rect 18049 3961 18061 3995
rect 18095 3992 18107 3995
rect 18800 3992 18828 4032
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 18095 3964 18828 3992
rect 18877 3995 18935 4001
rect 18095 3961 18107 3964
rect 18049 3955 18107 3961
rect 18877 3961 18889 3995
rect 18923 3992 18935 3995
rect 19610 3992 19616 4004
rect 18923 3964 19616 3992
rect 18923 3961 18935 3964
rect 18877 3955 18935 3961
rect 19610 3952 19616 3964
rect 19668 3952 19674 4004
rect 19904 4001 19932 4100
rect 19889 3995 19947 4001
rect 19889 3961 19901 3995
rect 19935 3992 19947 3995
rect 20346 3992 20352 4004
rect 19935 3964 20352 3992
rect 19935 3961 19947 3964
rect 19889 3955 19947 3961
rect 20346 3952 20352 3964
rect 20404 3952 20410 4004
rect 15068 3896 16988 3924
rect 15068 3884 15074 3896
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 20070 3924 20076 3936
rect 19024 3896 19069 3924
rect 20031 3896 20076 3924
rect 19024 3884 19030 3896
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2041 3723 2099 3729
rect 2041 3720 2053 3723
rect 2004 3692 2053 3720
rect 2004 3680 2010 3692
rect 2041 3689 2053 3692
rect 2087 3689 2099 3723
rect 2041 3683 2099 3689
rect 4065 3723 4123 3729
rect 4065 3689 4077 3723
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4080 3652 4108 3683
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 4304 3692 5181 3720
rect 4304 3680 4310 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 5997 3723 6055 3729
rect 5997 3689 6009 3723
rect 6043 3689 6055 3723
rect 8662 3720 8668 3732
rect 5997 3683 6055 3689
rect 6104 3692 7696 3720
rect 3436 3624 4108 3652
rect 2498 3584 2504 3596
rect 2459 3556 2504 3584
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 2590 3544 2596 3596
rect 2648 3584 2654 3596
rect 3326 3584 3332 3596
rect 2648 3556 2693 3584
rect 3252 3556 3332 3584
rect 2648 3544 2654 3556
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3252 3525 3280 3556
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2832 3488 3249 3516
rect 2832 3476 2838 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3329 3451 3387 3457
rect 3329 3417 3341 3451
rect 3375 3448 3387 3451
rect 3436 3448 3464 3624
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 4430 3652 4436 3664
rect 4212 3624 4436 3652
rect 4212 3612 4218 3624
rect 4430 3612 4436 3624
rect 4488 3652 4494 3664
rect 4985 3655 5043 3661
rect 4985 3652 4997 3655
rect 4488 3624 4997 3652
rect 4488 3612 4494 3624
rect 4985 3621 4997 3624
rect 5031 3652 5043 3655
rect 5902 3652 5908 3664
rect 5031 3624 5908 3652
rect 5031 3621 5043 3624
rect 4985 3615 5043 3621
rect 5902 3612 5908 3624
rect 5960 3652 5966 3664
rect 6012 3652 6040 3683
rect 5960 3624 6040 3652
rect 5960 3612 5966 3624
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 4522 3584 4528 3596
rect 3559 3556 4528 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4709 3587 4767 3593
rect 4709 3553 4721 3587
rect 4755 3584 4767 3587
rect 4890 3584 4896 3596
rect 4755 3556 4896 3584
rect 4755 3553 4767 3556
rect 4709 3547 4767 3553
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 5626 3584 5632 3596
rect 5587 3556 5632 3584
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 5994 3584 6000 3596
rect 5859 3556 6000 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 5994 3544 6000 3556
rect 6052 3544 6058 3596
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 4154 3516 4160 3528
rect 4019 3488 4160 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 6104 3516 6132 3692
rect 7668 3652 7696 3692
rect 8036 3692 8340 3720
rect 8623 3692 8668 3720
rect 8036 3652 8064 3692
rect 7668 3624 8064 3652
rect 8312 3652 8340 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 10594 3720 10600 3732
rect 8772 3692 10600 3720
rect 8772 3652 8800 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 11664 3692 12020 3720
rect 11664 3680 11670 3692
rect 10410 3652 10416 3664
rect 8312 3624 8800 3652
rect 10371 3624 10416 3652
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8202 3584 8208 3596
rect 8159 3556 8208 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 5583 3488 6132 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 6178 3476 6184 3528
rect 6236 3516 6242 3528
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 6236 3488 7665 3516
rect 6236 3476 6242 3488
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 3375 3420 3464 3448
rect 3375 3417 3387 3420
rect 3329 3411 3387 3417
rect 3878 3408 3884 3460
rect 3936 3448 3942 3460
rect 4525 3451 4583 3457
rect 4525 3448 4537 3451
rect 3936 3420 4537 3448
rect 3936 3408 3942 3420
rect 4525 3417 4537 3420
rect 4571 3417 4583 3451
rect 4525 3411 4583 3417
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6196 3448 6224 3476
rect 5960 3420 6224 3448
rect 6448 3451 6506 3457
rect 5960 3408 5966 3420
rect 6448 3417 6460 3451
rect 6494 3448 6506 3451
rect 6494 3420 7052 3448
rect 6494 3417 6506 3420
rect 6448 3411 6506 3417
rect 2406 3380 2412 3392
rect 2367 3352 2412 3380
rect 2406 3340 2412 3352
rect 2464 3340 2470 3392
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 3142 3380 3148 3392
rect 2915 3352 3148 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 3292 3352 4445 3380
rect 3292 3340 3298 3352
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 7024 3380 7052 3420
rect 7466 3380 7472 3392
rect 7024 3352 7472 3380
rect 4433 3343 4491 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3380 7619 3383
rect 8128 3380 8156 3547
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 11992 3593 12020 3692
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 12308 3692 14105 3720
rect 12308 3680 12314 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15749 3723 15807 3729
rect 15749 3720 15761 3723
rect 14792 3692 15761 3720
rect 14792 3680 14798 3692
rect 15749 3689 15761 3692
rect 15795 3689 15807 3723
rect 15749 3683 15807 3689
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 17313 3723 17371 3729
rect 16172 3692 16804 3720
rect 16172 3680 16178 3692
rect 12345 3655 12403 3661
rect 12345 3621 12357 3655
rect 12391 3652 12403 3655
rect 16482 3652 16488 3664
rect 12391 3624 12940 3652
rect 12391 3621 12403 3624
rect 12345 3615 12403 3621
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8941 3519 8999 3525
rect 8352 3488 8708 3516
rect 8352 3476 8358 3488
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 8570 3448 8576 3460
rect 8251 3420 8576 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 8680 3448 8708 3488
rect 8941 3485 8953 3519
rect 8987 3516 8999 3519
rect 9030 3516 9036 3528
rect 8987 3488 9036 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9030 3476 9036 3488
rect 9088 3516 9094 3528
rect 9490 3516 9496 3528
rect 9088 3488 9496 3516
rect 9088 3476 9094 3488
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 12158 3516 12164 3528
rect 12119 3488 12164 3516
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12802 3516 12808 3528
rect 12400 3488 12808 3516
rect 12400 3476 12406 3488
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 12912 3516 12940 3624
rect 14108 3624 14964 3652
rect 13814 3516 13820 3528
rect 12912 3488 13820 3516
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 13964 3488 14009 3516
rect 13964 3476 13970 3488
rect 9186 3451 9244 3457
rect 9186 3448 9198 3451
rect 8680 3420 9198 3448
rect 9186 3417 9198 3420
rect 9232 3417 9244 3451
rect 9186 3411 9244 3417
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 11732 3451 11790 3457
rect 9824 3420 11652 3448
rect 9824 3408 9830 3420
rect 7607 3352 8156 3380
rect 8297 3383 8355 3389
rect 7607 3349 7619 3352
rect 7561 3343 7619 3349
rect 8297 3349 8309 3383
rect 8343 3380 8355 3383
rect 9030 3380 9036 3392
rect 8343 3352 9036 3380
rect 8343 3349 8355 3352
rect 8297 3343 8355 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 10318 3380 10324 3392
rect 10279 3352 10324 3380
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10597 3383 10655 3389
rect 10597 3349 10609 3383
rect 10643 3380 10655 3383
rect 10686 3380 10692 3392
rect 10643 3352 10692 3380
rect 10643 3349 10655 3352
rect 10597 3343 10655 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11624 3380 11652 3420
rect 11732 3417 11744 3451
rect 11778 3448 11790 3451
rect 12066 3448 12072 3460
rect 11778 3420 12072 3448
rect 11778 3417 11790 3420
rect 11732 3411 11790 3417
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 13446 3448 13452 3460
rect 12406 3420 13452 3448
rect 12406 3380 12434 3420
rect 13446 3408 13452 3420
rect 13504 3408 13510 3460
rect 13722 3457 13728 3460
rect 13664 3451 13728 3457
rect 13664 3448 13676 3451
rect 13635 3420 13676 3448
rect 13664 3417 13676 3420
rect 13710 3417 13728 3451
rect 13664 3411 13728 3417
rect 13722 3408 13728 3411
rect 13780 3448 13786 3460
rect 14108 3448 14136 3624
rect 14936 3596 14964 3624
rect 15948 3624 16488 3652
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 14700 3556 14745 3584
rect 14700 3544 14706 3556
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 14516 3488 15301 3516
rect 14516 3476 14522 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 15948 3516 15976 3624
rect 16482 3612 16488 3624
rect 16540 3612 16546 3664
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16301 3587 16359 3593
rect 16301 3584 16313 3587
rect 16080 3556 16313 3584
rect 16080 3544 16086 3556
rect 16301 3553 16313 3556
rect 16347 3553 16359 3587
rect 16776 3584 16804 3692
rect 17313 3689 17325 3723
rect 17359 3720 17371 3723
rect 17678 3720 17684 3732
rect 17359 3692 17684 3720
rect 17359 3689 17371 3692
rect 17313 3683 17371 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18012 3692 18153 3720
rect 18012 3680 18018 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 19116 3692 19257 3720
rect 19116 3680 19122 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17586 3652 17592 3664
rect 17267 3624 17592 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 18966 3652 18972 3664
rect 17788 3624 18972 3652
rect 17788 3593 17816 3624
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 17773 3587 17831 3593
rect 16776 3556 17724 3584
rect 16301 3547 16359 3553
rect 15436 3488 15976 3516
rect 16117 3519 16175 3525
rect 15436 3476 15442 3488
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16390 3516 16396 3528
rect 16163 3488 16396 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16390 3476 16396 3488
rect 16448 3516 16454 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16448 3488 16957 3516
rect 16448 3476 16454 3488
rect 16945 3485 16957 3488
rect 16991 3516 17003 3519
rect 17402 3516 17408 3528
rect 16991 3488 17408 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 17696 3516 17724 3556
rect 17773 3553 17785 3587
rect 17819 3553 17831 3587
rect 17773 3547 17831 3553
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 18693 3587 18751 3593
rect 18693 3584 18705 3587
rect 17920 3556 17965 3584
rect 18064 3556 18705 3584
rect 17920 3544 17926 3556
rect 18064 3516 18092 3556
rect 18693 3553 18705 3556
rect 18739 3584 18751 3587
rect 19518 3584 19524 3596
rect 18739 3556 19524 3584
rect 18739 3553 18751 3556
rect 18693 3547 18751 3553
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 17696 3488 18092 3516
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 19058 3516 19064 3528
rect 18647 3488 19064 3516
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 16761 3451 16819 3457
rect 16761 3448 16773 3451
rect 13780 3420 14136 3448
rect 16224 3420 16773 3448
rect 13780 3408 13786 3420
rect 16224 3392 16252 3420
rect 16761 3417 16773 3420
rect 16807 3417 16819 3451
rect 16761 3411 16819 3417
rect 17681 3451 17739 3457
rect 17681 3417 17693 3451
rect 17727 3448 17739 3451
rect 17954 3448 17960 3460
rect 17727 3420 17960 3448
rect 17727 3417 17739 3420
rect 17681 3411 17739 3417
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 18509 3451 18567 3457
rect 18509 3448 18521 3451
rect 18472 3420 18521 3448
rect 18472 3408 18478 3420
rect 18509 3417 18521 3420
rect 18555 3448 18567 3451
rect 18969 3451 19027 3457
rect 18969 3448 18981 3451
rect 18555 3420 18981 3448
rect 18555 3417 18567 3420
rect 18509 3411 18567 3417
rect 18969 3417 18981 3420
rect 19015 3417 19027 3451
rect 18969 3411 19027 3417
rect 12526 3380 12532 3392
rect 11624 3352 12434 3380
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 14424 3352 14473 3380
rect 14424 3340 14430 3352
rect 14461 3349 14473 3352
rect 14507 3349 14519 3383
rect 14918 3380 14924 3392
rect 14879 3352 14924 3380
rect 14461 3343 14519 3349
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 16264 3352 16309 3380
rect 16264 3340 16270 3352
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 16540 3352 16681 3380
rect 16540 3340 16546 3352
rect 16669 3349 16681 3352
rect 16715 3380 16727 3383
rect 19702 3380 19708 3392
rect 16715 3352 19708 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2464 3148 2697 3176
rect 2464 3136 2470 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 2685 3139 2743 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3510 3176 3516 3188
rect 3292 3148 3516 3176
rect 3292 3136 3298 3148
rect 3510 3136 3516 3148
rect 3568 3176 3574 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3568 3148 3709 3176
rect 3568 3136 3574 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7374 3176 7380 3188
rect 7331 3148 7380 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 9214 3176 9220 3188
rect 8987 3148 9220 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 12618 3176 12624 3188
rect 11379 3148 12624 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 13633 3179 13691 3185
rect 13633 3176 13645 3179
rect 12860 3148 13645 3176
rect 12860 3136 12866 3148
rect 13633 3145 13645 3148
rect 13679 3145 13691 3179
rect 13633 3139 13691 3145
rect 14001 3179 14059 3185
rect 14001 3145 14013 3179
rect 14047 3176 14059 3179
rect 14918 3176 14924 3188
rect 14047 3148 14924 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 15160 3148 16405 3176
rect 15160 3136 15166 3148
rect 16393 3145 16405 3148
rect 16439 3145 16451 3179
rect 16393 3139 16451 3145
rect 2958 3068 2964 3120
rect 3016 3108 3022 3120
rect 6638 3108 6644 3120
rect 3016 3080 6644 3108
rect 3016 3068 3022 3080
rect 6638 3068 6644 3080
rect 6696 3068 6702 3120
rect 7650 3108 7656 3120
rect 7116 3080 7656 3108
rect 3050 3040 3056 3052
rect 3011 3012 3056 3040
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3160 3012 4384 3040
rect 1854 2932 1860 2984
rect 1912 2972 1918 2984
rect 3160 2972 3188 3012
rect 1912 2944 3188 2972
rect 3237 2975 3295 2981
rect 1912 2932 1918 2944
rect 3237 2941 3249 2975
rect 3283 2941 3295 2975
rect 4356 2972 4384 3012
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 4488 3012 5733 3040
rect 4488 3000 4494 3012
rect 5721 3009 5733 3012
rect 5767 3040 5779 3043
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5767 3012 6377 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 7116 3040 7144 3080
rect 7650 3068 7656 3080
rect 7708 3108 7714 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 7708 3080 8217 3108
rect 7708 3068 7714 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 10198 3111 10256 3117
rect 10198 3108 10210 3111
rect 8205 3071 8263 3077
rect 8864 3080 10210 3108
rect 6365 3003 6423 3009
rect 6656 3012 7144 3040
rect 6656 2981 6684 3012
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7248 3012 7389 3040
rect 7248 3000 7254 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 4356 2944 6653 2972
rect 3237 2935 3295 2941
rect 6641 2941 6653 2944
rect 6687 2941 6699 2975
rect 6914 2972 6920 2984
rect 6875 2944 6920 2972
rect 6641 2935 6699 2941
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 3252 2904 3280 2935
rect 6914 2932 6920 2944
rect 6972 2932 6978 2984
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 7466 2972 7472 2984
rect 7340 2944 7472 2972
rect 7340 2932 7346 2944
rect 7466 2932 7472 2944
rect 7524 2972 7530 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7524 2944 7941 2972
rect 7524 2932 7530 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 8864 2981 8892 3080
rect 10198 3077 10210 3080
rect 10244 3108 10256 3111
rect 10318 3108 10324 3120
rect 10244 3080 10324 3108
rect 10244 3077 10256 3080
rect 10198 3071 10256 3077
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 11793 3111 11851 3117
rect 10560 3080 11560 3108
rect 10560 3068 10566 3080
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 8113 2975 8171 2981
rect 8113 2972 8125 2975
rect 8076 2944 8125 2972
rect 8076 2932 8082 2944
rect 8113 2941 8125 2944
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 2924 2876 3280 2904
rect 2924 2864 2930 2876
rect 6546 2864 6552 2916
rect 6604 2864 6610 2916
rect 7745 2907 7803 2913
rect 7745 2873 7757 2907
rect 7791 2904 7803 2907
rect 9048 2904 9076 3003
rect 9490 3000 9496 3052
rect 9548 3040 9554 3052
rect 9861 3043 9919 3049
rect 9548 3012 9674 3040
rect 9548 3000 9554 3012
rect 9646 2972 9674 3012
rect 9861 3009 9873 3043
rect 9907 3040 9919 3043
rect 10778 3040 10784 3052
rect 9907 3012 10784 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11532 3049 11560 3080
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 12158 3108 12164 3120
rect 11839 3080 12164 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 13274 3111 13332 3117
rect 13274 3108 13286 3111
rect 12584 3080 13286 3108
rect 12584 3068 12590 3080
rect 13274 3077 13286 3080
rect 13320 3108 13332 3111
rect 13320 3080 13492 3108
rect 13320 3077 13332 3080
rect 13274 3071 13332 3077
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 13464 3040 13492 3080
rect 13538 3068 13544 3120
rect 13596 3108 13602 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13596 3080 14105 3108
rect 13596 3068 13602 3080
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 16206 3108 16212 3120
rect 14093 3071 14151 3077
rect 14752 3080 16212 3108
rect 14642 3040 14648 3052
rect 13464 3012 14648 3040
rect 11517 3003 11575 3009
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9646 2944 9965 2972
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 13538 2972 13544 2984
rect 13499 2944 13544 2972
rect 9953 2935 10011 2941
rect 13538 2932 13544 2944
rect 13596 2972 13602 2984
rect 13906 2972 13912 2984
rect 13596 2944 13912 2972
rect 13596 2932 13602 2944
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14200 2981 14228 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 14752 3049 14780 3080
rect 16206 3068 16212 3080
rect 16264 3068 16270 3120
rect 17586 3108 17592 3120
rect 17328 3080 17592 3108
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 14737 3003 14795 3009
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 14752 2972 14780 3003
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15286 3040 15292 3052
rect 15247 3012 15292 3040
rect 15286 3000 15292 3012
rect 15344 3000 15350 3052
rect 15838 3040 15844 3052
rect 15799 3012 15844 3040
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 16666 3040 16672 3052
rect 16356 3012 16672 3040
rect 16356 3000 16362 3012
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17328 3049 17356 3080
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 17770 3040 17776 3052
rect 17460 3012 17505 3040
rect 17731 3012 17776 3040
rect 17460 3000 17466 3012
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18782 3000 18788 3052
rect 18840 3040 18846 3052
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18840 3012 18889 3040
rect 18840 3000 18846 3012
rect 18877 3009 18889 3012
rect 18923 3040 18935 3043
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18923 3012 19257 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 15562 2972 15568 2984
rect 14332 2944 14780 2972
rect 15523 2944 15568 2972
rect 14332 2932 14338 2944
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 16114 2972 16120 2984
rect 16075 2944 16120 2972
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 9766 2904 9772 2916
rect 7791 2876 9076 2904
rect 9324 2876 9772 2904
rect 7791 2873 7803 2876
rect 7745 2867 7803 2873
rect 3878 2836 3884 2848
rect 3839 2808 3884 2836
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4985 2839 5043 2845
rect 4985 2805 4997 2839
rect 5031 2836 5043 2839
rect 5074 2836 5080 2848
rect 5031 2808 5080 2836
rect 5031 2805 5043 2808
rect 4985 2799 5043 2805
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 6564 2836 6592 2864
rect 9324 2836 9352 2876
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 11256 2876 12434 2904
rect 6564 2808 9352 2836
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9582 2836 9588 2848
rect 9447 2808 9588 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9677 2839 9735 2845
rect 9677 2805 9689 2839
rect 9723 2836 9735 2839
rect 11256 2836 11284 2876
rect 9723 2808 11284 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 12124 2808 12173 2836
rect 12124 2796 12130 2808
rect 12161 2805 12173 2808
rect 12207 2805 12219 2839
rect 12406 2836 12434 2876
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 14921 2907 14979 2913
rect 14921 2904 14933 2907
rect 14424 2876 14933 2904
rect 14424 2864 14430 2876
rect 14921 2873 14933 2876
rect 14967 2873 14979 2907
rect 14921 2867 14979 2873
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 17129 2907 17187 2913
rect 17129 2904 17141 2907
rect 16264 2876 17141 2904
rect 16264 2864 16270 2876
rect 17129 2873 17141 2876
rect 17175 2873 17187 2907
rect 17129 2867 17187 2873
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 18782 2904 18788 2916
rect 18371 2876 18788 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 19061 2907 19119 2913
rect 19061 2873 19073 2907
rect 19107 2904 19119 2907
rect 19518 2904 19524 2916
rect 19107 2876 19524 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 13262 2836 13268 2848
rect 12406 2808 13268 2836
rect 12161 2799 12219 2805
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 13780 2808 14565 2836
rect 13780 2796 13786 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 16942 2836 16948 2848
rect 16899 2808 16948 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17368 2808 17601 2836
rect 17368 2796 17374 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 17589 2799 17647 2805
rect 17678 2796 17684 2848
rect 17736 2836 17742 2848
rect 17957 2839 18015 2845
rect 17957 2836 17969 2839
rect 17736 2808 17969 2836
rect 17736 2796 17742 2808
rect 17957 2805 17969 2808
rect 18003 2805 18015 2839
rect 17957 2799 18015 2805
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 18966 2836 18972 2848
rect 18739 2808 18972 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 18966 2796 18972 2808
rect 19024 2796 19030 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3050 2592 3056 2644
rect 3108 2632 3114 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3108 2604 3801 2632
rect 3108 2592 3114 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 6181 2635 6239 2641
rect 6181 2632 6193 2635
rect 5960 2604 6193 2632
rect 5960 2592 5966 2604
rect 6181 2601 6193 2604
rect 6227 2601 6239 2635
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 6181 2595 6239 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 7834 2632 7840 2644
rect 7699 2604 7840 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8941 2635 8999 2641
rect 8941 2601 8953 2635
rect 8987 2632 8999 2635
rect 9122 2632 9128 2644
rect 8987 2604 9128 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11287 2604 11897 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11885 2601 11897 2604
rect 11931 2632 11943 2635
rect 11931 2604 13317 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 1946 2524 1952 2576
rect 2004 2564 2010 2576
rect 3329 2567 3387 2573
rect 3329 2564 3341 2567
rect 2004 2536 3341 2564
rect 2004 2524 2010 2536
rect 3329 2533 3341 2536
rect 3375 2564 3387 2567
rect 3375 2536 4292 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 3605 2499 3663 2505
rect 3605 2465 3617 2499
rect 3651 2496 3663 2499
rect 4062 2496 4068 2508
rect 3651 2468 4068 2496
rect 3651 2465 3663 2468
rect 3605 2459 3663 2465
rect 3988 2360 4016 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4264 2505 4292 2536
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 9769 2567 9827 2573
rect 9769 2564 9781 2567
rect 7248 2536 9781 2564
rect 7248 2524 7254 2536
rect 9769 2533 9781 2536
rect 9815 2564 9827 2567
rect 11146 2564 11152 2576
rect 9815 2536 11152 2564
rect 9815 2533 9827 2536
rect 9769 2527 9827 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11701 2567 11759 2573
rect 11701 2533 11713 2567
rect 11747 2564 11759 2567
rect 12802 2564 12808 2576
rect 11747 2536 12808 2564
rect 11747 2533 11759 2536
rect 11701 2527 11759 2533
rect 12802 2524 12808 2536
rect 12860 2524 12866 2576
rect 13289 2564 13317 2604
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 14553 2635 14611 2641
rect 14553 2632 14565 2635
rect 13412 2604 14565 2632
rect 13412 2592 13418 2604
rect 14553 2601 14565 2604
rect 14599 2601 14611 2635
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 14553 2595 14611 2601
rect 13538 2564 13544 2576
rect 13289 2536 13544 2564
rect 13538 2524 13544 2536
rect 13596 2564 13602 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 13596 2536 13645 2564
rect 13596 2524 13602 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 4522 2496 4528 2508
rect 4479 2468 4528 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 7282 2496 7288 2508
rect 7055 2468 7288 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 7282 2456 7288 2468
rect 7340 2496 7346 2508
rect 8297 2499 8355 2505
rect 8297 2496 8309 2499
rect 7340 2468 8309 2496
rect 7340 2456 7346 2468
rect 8297 2465 8309 2468
rect 8343 2496 8355 2499
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8343 2468 9505 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 10778 2496 10784 2508
rect 9640 2468 10640 2496
rect 10739 2468 10784 2496
rect 9640 2456 9646 2468
rect 4154 2428 4160 2440
rect 4115 2400 4160 2428
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 5074 2437 5080 2440
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5068 2391 5080 2437
rect 5132 2428 5138 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 5132 2400 5168 2428
rect 6472 2400 8033 2428
rect 4816 2360 4844 2391
rect 5074 2388 5080 2391
rect 5132 2388 5138 2400
rect 3988 2332 4844 2360
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 6472 2369 6500 2400
rect 8021 2397 8033 2400
rect 8067 2428 8079 2431
rect 8386 2428 8392 2440
rect 8067 2400 8392 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 8536 2400 9321 2428
rect 8536 2388 8542 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10612 2437 10640 2468
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2496 12771 2499
rect 12759 2468 13032 2496
rect 12759 2465 12771 2468
rect 12713 2459 12771 2465
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 10008 2400 10057 2428
rect 10008 2388 10014 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11020 2400 11529 2428
rect 11020 2388 11026 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 11517 2391 11575 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13004 2437 13032 2468
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 14274 2496 14280 2508
rect 13504 2468 14280 2496
rect 13504 2456 13510 2468
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14568 2496 14596 2595
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17313 2635 17371 2641
rect 17313 2601 17325 2635
rect 17359 2632 17371 2635
rect 17402 2632 17408 2644
rect 17359 2604 17408 2632
rect 17359 2601 17371 2604
rect 17313 2595 17371 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 17770 2632 17776 2644
rect 17727 2604 17776 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 18138 2632 18144 2644
rect 18095 2604 18144 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18417 2635 18475 2641
rect 18417 2601 18429 2635
rect 18463 2632 18475 2635
rect 18506 2632 18512 2644
rect 18463 2604 18512 2632
rect 18463 2601 18475 2604
rect 18417 2595 18475 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 15470 2564 15476 2576
rect 14967 2536 15476 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 16209 2567 16267 2573
rect 16209 2533 16221 2567
rect 16255 2564 16267 2567
rect 17034 2564 17040 2576
rect 16255 2536 17040 2564
rect 16255 2533 16267 2536
rect 16209 2527 16267 2533
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 14568 2468 14872 2496
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14844 2428 14872 2468
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15252 2468 15853 2496
rect 15252 2456 15258 2468
rect 15488 2437 15516 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 15381 2431 15439 2437
rect 15381 2428 15393 2431
rect 14844 2400 15393 2428
rect 14737 2391 14795 2397
rect 15381 2397 15393 2400
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 6457 2363 6515 2369
rect 6457 2360 6469 2363
rect 5960 2332 6469 2360
rect 5960 2320 5966 2332
rect 6457 2329 6469 2332
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 6638 2320 6644 2372
rect 6696 2360 6702 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6696 2332 6745 2360
rect 6696 2320 6702 2332
rect 6733 2329 6745 2332
rect 6779 2360 6791 2363
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 6779 2332 8125 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 8113 2329 8125 2332
rect 8159 2360 8171 2363
rect 10321 2363 10379 2369
rect 8159 2332 9904 2360
rect 8159 2329 8171 2332
rect 8113 2323 8171 2329
rect 3694 2252 3700 2304
rect 3752 2292 3758 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 3752 2264 4721 2292
rect 3752 2252 3758 2264
rect 4709 2261 4721 2264
rect 4755 2292 4767 2295
rect 7098 2292 7104 2304
rect 4755 2264 7104 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 8478 2292 8484 2304
rect 7248 2264 7293 2292
rect 8439 2264 8484 2292
rect 7248 2252 7254 2264
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 8570 2252 8576 2304
rect 8628 2292 8634 2304
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8628 2264 8677 2292
rect 8628 2252 8634 2264
rect 8665 2261 8677 2264
rect 8711 2292 8723 2295
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 8711 2264 9413 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9876 2292 9904 2332
rect 10321 2329 10333 2363
rect 10367 2360 10379 2363
rect 14752 2360 14780 2391
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 15620 2400 16037 2428
rect 15620 2388 15626 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16172 2400 16865 2428
rect 16172 2388 16178 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18414 2360 18420 2372
rect 10367 2332 14780 2360
rect 17052 2332 18420 2360
rect 10367 2329 10379 2332
rect 10321 2323 10379 2329
rect 11238 2292 11244 2304
rect 9876 2264 11244 2292
rect 9401 2255 9459 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12584 2264 13185 2292
rect 12584 2252 12590 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 15160 2264 15209 2292
rect 15160 2252 15166 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15746 2292 15752 2304
rect 15703 2264 15752 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 17052 2301 17080 2332
rect 18414 2320 18420 2332
rect 18472 2320 18478 2372
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2261 17095 2295
rect 17037 2255 17095 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 2222 2048 2228 2100
rect 2280 2088 2286 2100
rect 3786 2088 3792 2100
rect 2280 2060 3792 2088
rect 2280 2048 2286 2060
rect 3786 2048 3792 2060
rect 3844 2048 3850 2100
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 7190 2088 7196 2100
rect 4028 2060 7196 2088
rect 4028 2048 4034 2060
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 3326 1980 3332 2032
rect 3384 2020 3390 2032
rect 5902 2020 5908 2032
rect 3384 1992 5908 2020
rect 3384 1980 3390 1992
rect 5902 1980 5908 1992
rect 5960 1980 5966 2032
rect 7098 1980 7104 2032
rect 7156 2020 7162 2032
rect 13170 2020 13176 2032
rect 7156 1992 13176 2020
rect 7156 1980 7162 1992
rect 13170 1980 13176 1992
rect 13228 1980 13234 2032
rect 2590 1912 2596 1964
rect 2648 1952 2654 1964
rect 8478 1952 8484 1964
rect 2648 1924 8484 1952
rect 2648 1912 2654 1924
rect 8478 1912 8484 1924
rect 8536 1912 8542 1964
rect 3786 1844 3792 1896
rect 3844 1884 3850 1896
rect 8570 1884 8576 1896
rect 3844 1856 8576 1884
rect 3844 1844 3850 1856
rect 8570 1844 8576 1856
rect 8628 1884 8634 1896
rect 12342 1884 12348 1896
rect 8628 1856 12348 1884
rect 8628 1844 8634 1856
rect 12342 1844 12348 1856
rect 12400 1844 12406 1896
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 9214 1544 9220 1556
rect 8536 1516 9220 1544
rect 8536 1504 8542 1516
rect 9214 1504 9220 1516
rect 9272 1504 9278 1556
rect 5718 1368 5724 1420
rect 5776 1408 5782 1420
rect 6270 1408 6276 1420
rect 5776 1380 6276 1408
rect 5776 1368 5782 1380
rect 6270 1368 6276 1380
rect 6328 1368 6334 1420
<< via1 >>
rect 3884 20952 3936 21004
rect 10968 20952 11020 21004
rect 4068 20748 4120 20800
rect 20536 20748 20588 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 940 20544 992 20596
rect 5816 20587 5868 20596
rect 5816 20553 5825 20587
rect 5825 20553 5859 20587
rect 5859 20553 5868 20587
rect 5816 20544 5868 20553
rect 10876 20544 10928 20596
rect 12348 20544 12400 20596
rect 15292 20544 15344 20596
rect 17132 20544 17184 20596
rect 20444 20544 20496 20596
rect 5080 20476 5132 20528
rect 5540 20408 5592 20460
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 5632 20340 5684 20349
rect 8300 20408 8352 20460
rect 10416 20451 10468 20460
rect 10416 20417 10425 20451
rect 10425 20417 10459 20451
rect 10459 20417 10468 20451
rect 10416 20408 10468 20417
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 1308 20272 1360 20324
rect 7104 20340 7156 20392
rect 20996 20519 21048 20528
rect 11520 20451 11572 20460
rect 11520 20417 11529 20451
rect 11529 20417 11563 20451
rect 11563 20417 11572 20451
rect 11520 20408 11572 20417
rect 14372 20408 14424 20460
rect 14464 20408 14516 20460
rect 17224 20408 17276 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 18972 20408 19024 20460
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 20996 20485 21005 20519
rect 21005 20485 21039 20519
rect 21039 20485 21048 20519
rect 20996 20476 21048 20485
rect 20076 20408 20128 20460
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 5908 20272 5960 20324
rect 10600 20272 10652 20324
rect 11704 20272 11756 20324
rect 12072 20340 12124 20392
rect 18420 20340 18472 20392
rect 21548 20340 21600 20392
rect 16764 20272 16816 20324
rect 17592 20272 17644 20324
rect 19340 20272 19392 20324
rect 19708 20272 19760 20324
rect 3700 20204 3752 20256
rect 4712 20204 4764 20256
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 5448 20204 5500 20256
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7380 20204 7432 20213
rect 7472 20247 7524 20256
rect 7472 20213 7481 20247
rect 7481 20213 7515 20247
rect 7515 20213 7524 20247
rect 7472 20204 7524 20213
rect 11152 20204 11204 20256
rect 12992 20204 13044 20256
rect 14740 20204 14792 20256
rect 15108 20247 15160 20256
rect 15108 20213 15117 20247
rect 15117 20213 15151 20247
rect 15151 20213 15160 20247
rect 15108 20204 15160 20213
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 17224 20204 17276 20256
rect 19892 20204 19944 20256
rect 20168 20204 20220 20256
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1676 20000 1728 20052
rect 5448 20000 5500 20052
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 7104 20043 7156 20052
rect 7104 20009 7113 20043
rect 7113 20009 7147 20043
rect 7147 20009 7156 20043
rect 7104 20000 7156 20009
rect 7656 20000 7708 20052
rect 11796 20000 11848 20052
rect 11980 20043 12032 20052
rect 11980 20009 11989 20043
rect 11989 20009 12023 20043
rect 12023 20009 12032 20043
rect 11980 20000 12032 20009
rect 13084 20000 13136 20052
rect 13544 20000 13596 20052
rect 14280 20000 14332 20052
rect 14648 20000 14700 20052
rect 15200 20000 15252 20052
rect 15660 20000 15712 20052
rect 16948 20000 17000 20052
rect 18604 20000 18656 20052
rect 7012 19932 7064 19984
rect 11060 19932 11112 19984
rect 7288 19907 7340 19916
rect 4160 19796 4212 19848
rect 5264 19796 5316 19848
rect 5632 19796 5684 19848
rect 7288 19873 7297 19907
rect 7297 19873 7331 19907
rect 7331 19873 7340 19907
rect 7288 19864 7340 19873
rect 7380 19864 7432 19916
rect 8668 19864 8720 19916
rect 7748 19796 7800 19848
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 11152 19864 11204 19916
rect 12716 19932 12768 19984
rect 11060 19839 11112 19848
rect 11060 19805 11079 19839
rect 11079 19805 11112 19839
rect 17776 19864 17828 19916
rect 18420 19907 18472 19916
rect 18420 19873 18429 19907
rect 18429 19873 18463 19907
rect 18463 19873 18472 19907
rect 18420 19864 18472 19873
rect 11060 19796 11112 19805
rect 11520 19796 11572 19848
rect 11704 19796 11756 19848
rect 12900 19839 12952 19848
rect 12900 19805 12909 19839
rect 12909 19805 12943 19839
rect 12943 19805 12952 19839
rect 12900 19796 12952 19805
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 3884 19728 3936 19780
rect 4712 19728 4764 19780
rect 2228 19703 2280 19712
rect 2228 19669 2237 19703
rect 2237 19669 2271 19703
rect 2271 19669 2280 19703
rect 2228 19660 2280 19669
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 2780 19660 2832 19712
rect 3056 19660 3108 19712
rect 3148 19660 3200 19712
rect 7196 19660 7248 19712
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8760 19703 8812 19712
rect 8392 19660 8444 19669
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 10508 19728 10560 19780
rect 10600 19728 10652 19780
rect 10784 19728 10836 19780
rect 12072 19728 12124 19780
rect 13176 19728 13228 19780
rect 14280 19796 14332 19848
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15476 19796 15528 19848
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 11796 19660 11848 19712
rect 15660 19796 15712 19848
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 18604 19796 18656 19848
rect 18972 19796 19024 19848
rect 20812 20000 20864 20052
rect 21548 20000 21600 20052
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 19616 19864 19668 19873
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20628 19864 20680 19916
rect 19800 19796 19852 19848
rect 20444 19796 20496 19848
rect 18512 19728 18564 19780
rect 20168 19728 20220 19780
rect 15936 19660 15988 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 3332 19499 3384 19508
rect 2044 19388 2096 19440
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 4712 19456 4764 19508
rect 5816 19499 5868 19508
rect 5816 19465 5825 19499
rect 5825 19465 5859 19499
rect 5859 19465 5868 19499
rect 5816 19456 5868 19465
rect 6460 19456 6512 19508
rect 7196 19499 7248 19508
rect 7196 19465 7205 19499
rect 7205 19465 7239 19499
rect 7239 19465 7248 19499
rect 7196 19456 7248 19465
rect 7472 19456 7524 19508
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 10416 19456 10468 19508
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 13820 19456 13872 19508
rect 15200 19456 15252 19508
rect 16028 19456 16080 19508
rect 16396 19456 16448 19508
rect 17500 19456 17552 19508
rect 17868 19499 17920 19508
rect 17868 19465 17877 19499
rect 17877 19465 17911 19499
rect 17911 19465 17920 19499
rect 17868 19456 17920 19465
rect 3148 19388 3200 19440
rect 2228 19320 2280 19372
rect 2596 19320 2648 19372
rect 2872 19320 2924 19372
rect 3056 19320 3108 19372
rect 4160 19320 4212 19372
rect 5172 19320 5224 19372
rect 5264 19363 5316 19372
rect 5264 19329 5284 19363
rect 5284 19329 5316 19363
rect 5264 19320 5316 19329
rect 5448 19320 5500 19372
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 7196 19320 7248 19372
rect 7748 19388 7800 19440
rect 8760 19388 8812 19440
rect 10968 19388 11020 19440
rect 13728 19388 13780 19440
rect 14464 19431 14516 19440
rect 10600 19363 10652 19372
rect 10600 19329 10609 19363
rect 10609 19329 10643 19363
rect 10643 19329 10652 19363
rect 10600 19320 10652 19329
rect 10876 19320 10928 19372
rect 11244 19320 11296 19372
rect 13176 19363 13228 19372
rect 2412 19184 2464 19236
rect 2872 19159 2924 19168
rect 2872 19125 2881 19159
rect 2881 19125 2915 19159
rect 2915 19125 2924 19159
rect 3240 19184 3292 19236
rect 2872 19116 2924 19125
rect 4160 19116 4212 19168
rect 5540 19184 5592 19236
rect 6000 19184 6052 19236
rect 6368 19184 6420 19236
rect 7104 19184 7156 19236
rect 8484 19252 8536 19304
rect 10784 19295 10836 19304
rect 10784 19261 10793 19295
rect 10793 19261 10827 19295
rect 10827 19261 10836 19295
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13820 19320 13872 19372
rect 14464 19397 14473 19431
rect 14473 19397 14507 19431
rect 14507 19397 14516 19431
rect 14464 19388 14516 19397
rect 15660 19388 15712 19440
rect 17592 19388 17644 19440
rect 18512 19499 18564 19508
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 18236 19388 18288 19440
rect 19708 19431 19760 19440
rect 19708 19397 19717 19431
rect 19717 19397 19751 19431
rect 19751 19397 19760 19431
rect 19708 19388 19760 19397
rect 20260 19431 20312 19440
rect 20260 19397 20269 19431
rect 20269 19397 20303 19431
rect 20303 19397 20312 19431
rect 20260 19388 20312 19397
rect 21180 19388 21232 19440
rect 21456 19388 21508 19440
rect 10784 19252 10836 19261
rect 13084 19252 13136 19304
rect 13544 19184 13596 19236
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 19340 19363 19392 19372
rect 16488 19295 16540 19304
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 19340 19329 19349 19363
rect 19349 19329 19383 19363
rect 19383 19329 19392 19363
rect 19340 19320 19392 19329
rect 16488 19252 16540 19261
rect 18604 19252 18656 19304
rect 19064 19252 19116 19304
rect 20444 19320 20496 19372
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 19892 19252 19944 19304
rect 8024 19116 8076 19168
rect 8300 19116 8352 19168
rect 12808 19116 12860 19168
rect 13636 19116 13688 19168
rect 14372 19116 14424 19168
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 17592 19159 17644 19168
rect 17592 19125 17601 19159
rect 17601 19125 17635 19159
rect 17635 19125 17644 19159
rect 17592 19116 17644 19125
rect 18788 19159 18840 19168
rect 18788 19125 18797 19159
rect 18797 19125 18831 19159
rect 18831 19125 18840 19159
rect 18788 19116 18840 19125
rect 19340 19116 19392 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 3332 18912 3384 18964
rect 4804 18912 4856 18964
rect 3148 18844 3200 18896
rect 3608 18844 3660 18896
rect 4160 18887 4212 18896
rect 4160 18853 4169 18887
rect 4169 18853 4203 18887
rect 4203 18853 4212 18887
rect 4160 18844 4212 18853
rect 4896 18844 4948 18896
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 2964 18776 3016 18828
rect 4528 18776 4580 18828
rect 2136 18708 2188 18760
rect 2872 18708 2924 18760
rect 4712 18819 4764 18828
rect 4712 18785 4721 18819
rect 4721 18785 4755 18819
rect 4755 18785 4764 18819
rect 4712 18776 4764 18785
rect 5540 18776 5592 18828
rect 5724 18819 5776 18828
rect 5724 18785 5733 18819
rect 5733 18785 5767 18819
rect 5767 18785 5776 18819
rect 5724 18776 5776 18785
rect 3240 18640 3292 18692
rect 572 18368 624 18420
rect 2320 18572 2372 18624
rect 3332 18572 3384 18624
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 5356 18640 5408 18692
rect 5908 18776 5960 18828
rect 6368 18819 6420 18828
rect 6368 18785 6377 18819
rect 6377 18785 6411 18819
rect 6411 18785 6420 18819
rect 6368 18776 6420 18785
rect 7196 18912 7248 18964
rect 7288 18912 7340 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 9588 18912 9640 18964
rect 10600 18912 10652 18964
rect 10968 18912 11020 18964
rect 8024 18844 8076 18896
rect 11796 18912 11848 18964
rect 12900 18912 12952 18964
rect 18972 18955 19024 18964
rect 18972 18921 18981 18955
rect 18981 18921 19015 18955
rect 19015 18921 19024 18955
rect 18972 18912 19024 18921
rect 19064 18912 19116 18964
rect 21364 18955 21416 18964
rect 21364 18921 21373 18955
rect 21373 18921 21407 18955
rect 21407 18921 21416 18955
rect 21364 18912 21416 18921
rect 8668 18776 8720 18828
rect 10876 18776 10928 18828
rect 13084 18844 13136 18896
rect 12808 18819 12860 18828
rect 12808 18785 12817 18819
rect 12817 18785 12851 18819
rect 12851 18785 12860 18819
rect 12808 18776 12860 18785
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14372 18819 14424 18828
rect 14372 18785 14381 18819
rect 14381 18785 14415 18819
rect 14415 18785 14424 18819
rect 14372 18776 14424 18785
rect 15568 18776 15620 18828
rect 20720 18844 20772 18896
rect 7012 18708 7064 18760
rect 6460 18683 6512 18692
rect 6460 18649 6469 18683
rect 6469 18649 6503 18683
rect 6503 18649 6512 18683
rect 6460 18640 6512 18649
rect 5724 18572 5776 18624
rect 5908 18572 5960 18624
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 7104 18640 7156 18692
rect 8024 18708 8076 18760
rect 7472 18640 7524 18692
rect 18972 18708 19024 18760
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 20444 18708 20496 18760
rect 21272 18708 21324 18760
rect 11704 18640 11756 18692
rect 11980 18640 12032 18692
rect 7380 18572 7432 18624
rect 9036 18572 9088 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9680 18572 9732 18624
rect 10692 18572 10744 18624
rect 10876 18572 10928 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 12624 18615 12676 18624
rect 12624 18581 12633 18615
rect 12633 18581 12667 18615
rect 12667 18581 12676 18615
rect 13360 18615 13412 18624
rect 12624 18572 12676 18581
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 15752 18572 15804 18624
rect 20996 18640 21048 18692
rect 22284 18572 22336 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2320 18368 2372 18420
rect 1308 18300 1360 18352
rect 3056 18300 3108 18352
rect 2320 18232 2372 18284
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 5264 18232 5316 18284
rect 5540 18343 5592 18352
rect 5540 18309 5558 18343
rect 5558 18309 5592 18343
rect 5540 18300 5592 18309
rect 8392 18368 8444 18420
rect 10048 18411 10100 18420
rect 5908 18232 5960 18284
rect 2872 18207 2924 18216
rect 2872 18173 2881 18207
rect 2881 18173 2915 18207
rect 2915 18173 2924 18207
rect 2872 18164 2924 18173
rect 3056 18207 3108 18216
rect 3056 18173 3065 18207
rect 3065 18173 3099 18207
rect 3099 18173 3108 18207
rect 3056 18164 3108 18173
rect 3792 18207 3844 18216
rect 3792 18173 3801 18207
rect 3801 18173 3835 18207
rect 3835 18173 3844 18207
rect 3792 18164 3844 18173
rect 4528 18164 4580 18216
rect 3976 18096 4028 18148
rect 2136 18028 2188 18080
rect 3608 18028 3660 18080
rect 4712 18096 4764 18148
rect 5172 18028 5224 18080
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 6736 18232 6788 18284
rect 8024 18300 8076 18352
rect 10048 18377 10057 18411
rect 10057 18377 10091 18411
rect 10091 18377 10100 18411
rect 10048 18368 10100 18377
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 11704 18300 11756 18352
rect 13084 18343 13136 18352
rect 7472 18232 7524 18284
rect 8484 18232 8536 18284
rect 12164 18232 12216 18284
rect 13084 18309 13093 18343
rect 13093 18309 13127 18343
rect 13127 18309 13136 18343
rect 13084 18300 13136 18309
rect 13544 18300 13596 18352
rect 14188 18368 14240 18420
rect 14464 18368 14516 18420
rect 15568 18411 15620 18420
rect 15568 18377 15577 18411
rect 15577 18377 15611 18411
rect 15611 18377 15620 18411
rect 15568 18368 15620 18377
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 20536 18411 20588 18420
rect 20536 18377 20545 18411
rect 20545 18377 20579 18411
rect 20579 18377 20588 18411
rect 20536 18368 20588 18377
rect 21456 18411 21508 18420
rect 21456 18377 21465 18411
rect 21465 18377 21499 18411
rect 21499 18377 21508 18411
rect 21456 18368 21508 18377
rect 17040 18300 17092 18352
rect 18328 18300 18380 18352
rect 7104 18164 7156 18216
rect 7288 18164 7340 18216
rect 8300 18164 8352 18216
rect 8668 18164 8720 18216
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 6736 18096 6788 18148
rect 7012 18028 7064 18080
rect 9036 18139 9088 18148
rect 9036 18105 9045 18139
rect 9045 18105 9079 18139
rect 9079 18105 9088 18139
rect 9036 18096 9088 18105
rect 9496 18096 9548 18148
rect 10968 18164 11020 18216
rect 11888 18164 11940 18216
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12808 18232 12860 18284
rect 12716 18207 12768 18216
rect 12716 18173 12725 18207
rect 12725 18173 12759 18207
rect 12759 18173 12768 18207
rect 12716 18164 12768 18173
rect 19524 18232 19576 18284
rect 21640 18300 21692 18352
rect 20444 18232 20496 18284
rect 20076 18164 20128 18216
rect 11980 18096 12032 18148
rect 19800 18096 19852 18148
rect 8392 18028 8444 18080
rect 11612 18028 11664 18080
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1768 17867 1820 17876
rect 1768 17833 1777 17867
rect 1777 17833 1811 17867
rect 1811 17833 1820 17867
rect 1768 17824 1820 17833
rect 4528 17867 4580 17876
rect 4528 17833 4537 17867
rect 4537 17833 4571 17867
rect 4571 17833 4580 17867
rect 4528 17824 4580 17833
rect 5264 17824 5316 17876
rect 5540 17824 5592 17876
rect 5908 17824 5960 17876
rect 6000 17824 6052 17876
rect 6552 17867 6604 17876
rect 6552 17833 6561 17867
rect 6561 17833 6595 17867
rect 6595 17833 6604 17867
rect 6552 17824 6604 17833
rect 6736 17824 6788 17876
rect 5816 17756 5868 17808
rect 6460 17799 6512 17808
rect 4896 17688 4948 17740
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 6460 17765 6469 17799
rect 6469 17765 6503 17799
rect 6503 17765 6512 17799
rect 6460 17756 6512 17765
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 1952 17663 2004 17672
rect 1952 17629 1961 17663
rect 1961 17629 1995 17663
rect 1995 17629 2004 17663
rect 1952 17620 2004 17629
rect 2780 17620 2832 17672
rect 3516 17620 3568 17672
rect 4528 17620 4580 17672
rect 4620 17620 4672 17672
rect 6000 17552 6052 17604
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 4252 17484 4304 17536
rect 5264 17484 5316 17536
rect 5540 17484 5592 17536
rect 5816 17527 5868 17536
rect 5816 17493 5825 17527
rect 5825 17493 5859 17527
rect 5859 17493 5868 17527
rect 6552 17620 6604 17672
rect 9312 17824 9364 17876
rect 9404 17824 9456 17876
rect 12072 17824 12124 17876
rect 12348 17824 12400 17876
rect 20444 17824 20496 17876
rect 21548 17867 21600 17876
rect 21548 17833 21557 17867
rect 21557 17833 21591 17867
rect 21591 17833 21600 17867
rect 21548 17824 21600 17833
rect 8484 17756 8536 17808
rect 9128 17756 9180 17808
rect 13360 17756 13412 17808
rect 19892 17756 19944 17808
rect 8300 17688 8352 17740
rect 9496 17731 9548 17740
rect 9496 17697 9505 17731
rect 9505 17697 9539 17731
rect 9539 17697 9548 17731
rect 9496 17688 9548 17697
rect 10232 17688 10284 17740
rect 10968 17688 11020 17740
rect 11704 17688 11756 17740
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 10692 17552 10744 17604
rect 12716 17620 12768 17672
rect 13084 17620 13136 17672
rect 14464 17663 14516 17672
rect 14464 17629 14498 17663
rect 14498 17629 14516 17663
rect 14464 17620 14516 17629
rect 15476 17620 15528 17672
rect 5816 17484 5868 17493
rect 8024 17484 8076 17536
rect 8208 17484 8260 17536
rect 8576 17484 8628 17536
rect 8760 17484 8812 17536
rect 11060 17484 11112 17536
rect 12532 17552 12584 17604
rect 12992 17552 13044 17604
rect 14740 17552 14792 17604
rect 11888 17527 11940 17536
rect 11888 17493 11897 17527
rect 11897 17493 11931 17527
rect 11931 17493 11940 17527
rect 11888 17484 11940 17493
rect 12716 17527 12768 17536
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 15384 17484 15436 17536
rect 15660 17620 15712 17672
rect 16212 17552 16264 17604
rect 21548 17552 21600 17604
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 16396 17484 16448 17536
rect 19616 17484 19668 17536
rect 20352 17484 20404 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 2872 17280 2924 17332
rect 2044 17212 2096 17264
rect 3608 17212 3660 17264
rect 5724 17280 5776 17332
rect 3884 17212 3936 17264
rect 7288 17280 7340 17332
rect 8208 17323 8260 17332
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 8668 17280 8720 17332
rect 9128 17280 9180 17332
rect 10232 17280 10284 17332
rect 11612 17280 11664 17332
rect 11796 17323 11848 17332
rect 11796 17289 11805 17323
rect 11805 17289 11839 17323
rect 11839 17289 11848 17323
rect 11796 17280 11848 17289
rect 5908 17212 5960 17264
rect 7104 17212 7156 17264
rect 5172 17144 5224 17196
rect 6920 17187 6972 17196
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7656 17144 7708 17196
rect 6092 17076 6144 17128
rect 4988 17008 5040 17060
rect 5356 17008 5408 17060
rect 7012 17076 7064 17128
rect 7196 17076 7248 17128
rect 10692 17144 10744 17196
rect 8392 17076 8444 17128
rect 4620 16940 4672 16992
rect 7472 17008 7524 17060
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 8300 16940 8352 16992
rect 9496 17076 9548 17128
rect 9680 17076 9732 17128
rect 11796 17076 11848 17128
rect 12992 17280 13044 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 15660 17280 15712 17332
rect 15752 17323 15804 17332
rect 15752 17289 15761 17323
rect 15761 17289 15795 17323
rect 15795 17289 15804 17323
rect 16396 17323 16448 17332
rect 15752 17280 15804 17289
rect 16396 17289 16405 17323
rect 16405 17289 16439 17323
rect 16439 17289 16448 17323
rect 16396 17280 16448 17289
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 21088 17280 21140 17332
rect 21364 17323 21416 17332
rect 21364 17289 21373 17323
rect 21373 17289 21407 17323
rect 21407 17289 21416 17323
rect 21364 17280 21416 17289
rect 12164 17212 12216 17264
rect 15292 17144 15344 17196
rect 15660 17144 15712 17196
rect 15844 17187 15896 17196
rect 15844 17153 15853 17187
rect 15853 17153 15887 17187
rect 15887 17153 15896 17187
rect 15844 17144 15896 17153
rect 19984 17187 20036 17196
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 12348 17076 12400 17128
rect 12808 17076 12860 17128
rect 13176 17076 13228 17128
rect 12072 17008 12124 17060
rect 12532 17008 12584 17060
rect 13084 17008 13136 17060
rect 13268 17008 13320 17060
rect 14280 17008 14332 17060
rect 15384 17076 15436 17128
rect 16120 17008 16172 17060
rect 12164 16940 12216 16992
rect 12992 16940 13044 16992
rect 16028 16940 16080 16992
rect 16764 16983 16816 16992
rect 16764 16949 16773 16983
rect 16773 16949 16807 16983
rect 16807 16949 16816 16983
rect 16764 16940 16816 16949
rect 19892 16940 19944 16992
rect 20812 16940 20864 16992
rect 22468 16940 22520 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 4896 16736 4948 16788
rect 5908 16736 5960 16788
rect 7104 16736 7156 16788
rect 7932 16736 7984 16788
rect 8024 16736 8076 16788
rect 2044 16668 2096 16720
rect 5724 16668 5776 16720
rect 6092 16711 6144 16720
rect 6092 16677 6101 16711
rect 6101 16677 6135 16711
rect 6135 16677 6144 16711
rect 6092 16668 6144 16677
rect 4620 16600 4672 16652
rect 7012 16643 7064 16652
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 2596 16575 2648 16584
rect 2596 16541 2605 16575
rect 2605 16541 2639 16575
rect 2639 16541 2648 16575
rect 2596 16532 2648 16541
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 4988 16575 5040 16584
rect 4988 16541 5011 16575
rect 5011 16541 5040 16575
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 7472 16600 7524 16652
rect 8024 16600 8076 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 8576 16736 8628 16788
rect 9404 16736 9456 16788
rect 8484 16668 8536 16720
rect 11244 16668 11296 16720
rect 4988 16532 5040 16541
rect 7288 16532 7340 16584
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10048 16600 10100 16609
rect 11704 16736 11756 16788
rect 11888 16736 11940 16788
rect 14280 16736 14332 16788
rect 15660 16736 15712 16788
rect 15752 16736 15804 16788
rect 19524 16736 19576 16788
rect 21088 16736 21140 16788
rect 17868 16668 17920 16720
rect 11612 16643 11664 16652
rect 10140 16532 10192 16584
rect 11060 16532 11112 16584
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 14464 16600 14516 16652
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 3148 16464 3200 16516
rect 3056 16396 3108 16448
rect 3700 16396 3752 16448
rect 4068 16464 4120 16516
rect 5816 16464 5868 16516
rect 6460 16464 6512 16516
rect 7012 16464 7064 16516
rect 10968 16464 11020 16516
rect 13176 16532 13228 16584
rect 19984 16600 20036 16652
rect 3884 16396 3936 16448
rect 6828 16396 6880 16448
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 11796 16396 11848 16448
rect 13636 16464 13688 16516
rect 15200 16507 15252 16516
rect 15200 16473 15218 16507
rect 15218 16473 15252 16507
rect 15200 16464 15252 16473
rect 15384 16464 15436 16516
rect 17408 16532 17460 16584
rect 16764 16507 16816 16516
rect 16304 16396 16356 16448
rect 16764 16473 16773 16507
rect 16773 16473 16807 16507
rect 16807 16473 16816 16507
rect 16764 16464 16816 16473
rect 17592 16464 17644 16516
rect 20168 16464 20220 16516
rect 22560 16464 22612 16516
rect 17040 16396 17092 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 3884 16192 3936 16244
rect 5540 16192 5592 16244
rect 5816 16235 5868 16244
rect 5816 16201 5825 16235
rect 5825 16201 5859 16235
rect 5859 16201 5868 16235
rect 5816 16192 5868 16201
rect 7288 16192 7340 16244
rect 2228 15895 2280 15904
rect 2228 15861 2237 15895
rect 2237 15861 2271 15895
rect 2271 15861 2280 15895
rect 2228 15852 2280 15861
rect 2872 15988 2924 16040
rect 3424 16056 3476 16108
rect 3884 16056 3936 16108
rect 4252 16031 4304 16040
rect 2688 15852 2740 15904
rect 2964 15852 3016 15904
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 4712 16124 4764 16176
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 6920 16124 6972 16176
rect 9496 16192 9548 16244
rect 9588 16192 9640 16244
rect 12532 16192 12584 16244
rect 13176 16192 13228 16244
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 15752 16192 15804 16244
rect 15844 16192 15896 16244
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 17868 16192 17920 16244
rect 20628 16235 20680 16244
rect 20628 16201 20637 16235
rect 20637 16201 20671 16235
rect 20671 16201 20680 16235
rect 20628 16192 20680 16201
rect 21088 16192 21140 16244
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 5724 16056 5776 16108
rect 4896 15988 4948 16040
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 3700 15920 3752 15972
rect 4804 15920 4856 15972
rect 6828 15988 6880 16040
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 7472 15988 7524 15997
rect 9220 16124 9272 16176
rect 10048 16124 10100 16176
rect 10692 16124 10744 16176
rect 13452 16124 13504 16176
rect 14280 16124 14332 16176
rect 9128 16056 9180 16108
rect 11152 16056 11204 16108
rect 13636 16056 13688 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 12348 16031 12400 16040
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 12348 15997 12357 16031
rect 12357 15997 12391 16031
rect 12391 15997 12400 16031
rect 12348 15988 12400 15997
rect 15200 16124 15252 16176
rect 16304 16124 16356 16176
rect 18236 16124 18288 16176
rect 18512 16124 18564 16176
rect 14740 16056 14792 16108
rect 16120 16056 16172 16108
rect 17132 16056 17184 16108
rect 19984 16056 20036 16108
rect 20904 16056 20956 16108
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 16672 15988 16724 16040
rect 17776 15988 17828 16040
rect 16396 15920 16448 15972
rect 18420 15988 18472 16040
rect 18788 15988 18840 16040
rect 20628 15988 20680 16040
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 17868 15852 17920 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1860 15648 1912 15700
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 4160 15691 4212 15700
rect 2780 15648 2832 15657
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 4620 15648 4672 15700
rect 6000 15691 6052 15700
rect 6000 15657 6009 15691
rect 6009 15657 6043 15691
rect 6043 15657 6052 15691
rect 6000 15648 6052 15657
rect 7472 15648 7524 15700
rect 7656 15648 7708 15700
rect 2228 15444 2280 15496
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3424 15555 3476 15564
rect 3424 15521 3433 15555
rect 3433 15521 3467 15555
rect 3467 15521 3476 15555
rect 3424 15512 3476 15521
rect 6828 15580 6880 15632
rect 8392 15580 8444 15632
rect 9220 15580 9272 15632
rect 12440 15648 12492 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 14464 15648 14516 15700
rect 12716 15580 12768 15632
rect 13912 15580 13964 15632
rect 17040 15648 17092 15700
rect 17776 15648 17828 15700
rect 21364 15691 21416 15700
rect 21364 15657 21373 15691
rect 21373 15657 21407 15691
rect 21407 15657 21416 15691
rect 21364 15648 21416 15657
rect 16304 15580 16356 15632
rect 5172 15444 5224 15496
rect 5724 15444 5776 15496
rect 6920 15512 6972 15564
rect 7288 15555 7340 15564
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12900 15512 12952 15564
rect 14832 15512 14884 15564
rect 15476 15512 15528 15564
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 7380 15444 7432 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10784 15487 10836 15496
rect 10784 15453 10818 15487
rect 10818 15453 10836 15487
rect 10784 15444 10836 15453
rect 12072 15444 12124 15496
rect 4896 15376 4948 15428
rect 6552 15376 6604 15428
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 4804 15308 4856 15360
rect 5540 15308 5592 15360
rect 9220 15376 9272 15428
rect 10600 15376 10652 15428
rect 12256 15376 12308 15428
rect 10876 15308 10928 15360
rect 11888 15308 11940 15360
rect 12440 15308 12492 15360
rect 12900 15308 12952 15360
rect 12992 15308 13044 15360
rect 14740 15376 14792 15428
rect 13452 15308 13504 15360
rect 15016 15444 15068 15496
rect 16672 15487 16724 15496
rect 16672 15453 16706 15487
rect 16706 15453 16724 15487
rect 16672 15444 16724 15453
rect 16948 15444 17000 15496
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 18328 15487 18380 15496
rect 18328 15453 18337 15487
rect 18337 15453 18371 15487
rect 18371 15453 18380 15487
rect 18328 15444 18380 15453
rect 19616 15487 19668 15496
rect 19616 15453 19625 15487
rect 19625 15453 19659 15487
rect 19659 15453 19668 15487
rect 19616 15444 19668 15453
rect 15384 15419 15436 15428
rect 15384 15385 15393 15419
rect 15393 15385 15427 15419
rect 15427 15385 15436 15419
rect 15384 15376 15436 15385
rect 17500 15376 17552 15428
rect 16120 15308 16172 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 21088 15308 21140 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 5632 15104 5684 15156
rect 6920 15104 6972 15156
rect 7472 15104 7524 15156
rect 8116 15104 8168 15156
rect 9128 15104 9180 15156
rect 9404 15104 9456 15156
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 3056 15036 3108 15088
rect 3148 15036 3200 15088
rect 7748 15036 7800 15088
rect 11244 15104 11296 15156
rect 11888 15104 11940 15156
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 16580 15104 16632 15156
rect 16948 15104 17000 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 10416 15079 10468 15088
rect 10416 15045 10425 15079
rect 10425 15045 10459 15079
rect 10459 15045 10468 15079
rect 10416 15036 10468 15045
rect 16212 15036 16264 15088
rect 16304 15036 16356 15088
rect 3976 14968 4028 15020
rect 5172 14968 5224 15020
rect 5632 14968 5684 15020
rect 6828 14968 6880 15020
rect 3884 14900 3936 14952
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 7012 14900 7064 14952
rect 7840 14900 7892 14952
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 9588 14900 9640 14952
rect 2780 14764 2832 14816
rect 6368 14832 6420 14884
rect 7288 14832 7340 14884
rect 7380 14832 7432 14884
rect 10048 14832 10100 14884
rect 4344 14764 4396 14816
rect 4528 14764 4580 14816
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 8668 14764 8720 14816
rect 9404 14764 9456 14816
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 16396 14968 16448 15020
rect 17776 15036 17828 15088
rect 19984 15079 20036 15088
rect 19984 15045 19993 15079
rect 19993 15045 20027 15079
rect 20027 15045 20036 15079
rect 19984 15036 20036 15045
rect 17316 14968 17368 15020
rect 18880 14968 18932 15020
rect 19708 15011 19760 15020
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 12532 14900 12584 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 14280 14900 14332 14952
rect 14464 14900 14516 14952
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 15844 14764 15896 14816
rect 16212 14764 16264 14816
rect 17224 14764 17276 14816
rect 19800 14832 19852 14884
rect 18236 14764 18288 14816
rect 21180 14764 21232 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 2872 14603 2924 14612
rect 2872 14569 2881 14603
rect 2881 14569 2915 14603
rect 2915 14569 2924 14603
rect 2872 14560 2924 14569
rect 1584 14535 1636 14544
rect 1584 14501 1593 14535
rect 1593 14501 1627 14535
rect 1627 14501 1636 14535
rect 1584 14492 1636 14501
rect 2780 14492 2832 14544
rect 3332 14492 3384 14544
rect 4068 14492 4120 14544
rect 2596 14424 2648 14476
rect 5724 14560 5776 14612
rect 7748 14560 7800 14612
rect 9864 14603 9916 14612
rect 9588 14492 9640 14544
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 11888 14560 11940 14612
rect 12532 14560 12584 14612
rect 14004 14560 14056 14612
rect 15200 14560 15252 14612
rect 19984 14560 20036 14612
rect 20904 14560 20956 14612
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 4988 14424 5040 14476
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 5540 14356 5592 14408
rect 7288 14356 7340 14408
rect 3332 14288 3384 14340
rect 3424 14331 3476 14340
rect 3424 14297 3433 14331
rect 3433 14297 3467 14331
rect 3467 14297 3476 14331
rect 3424 14288 3476 14297
rect 7840 14288 7892 14340
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 9864 14424 9916 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 10324 14424 10376 14476
rect 13820 14424 13872 14476
rect 15844 14467 15896 14476
rect 8116 14356 8168 14408
rect 8668 14356 8720 14408
rect 9588 14356 9640 14408
rect 10508 14356 10560 14408
rect 12532 14399 12584 14408
rect 12532 14365 12566 14399
rect 12566 14365 12584 14399
rect 10692 14288 10744 14340
rect 11060 14331 11112 14340
rect 11060 14297 11094 14331
rect 11094 14297 11112 14331
rect 12532 14356 12584 14365
rect 11060 14288 11112 14297
rect 12440 14288 12492 14340
rect 14648 14356 14700 14408
rect 15844 14433 15853 14467
rect 15853 14433 15887 14467
rect 15887 14433 15896 14467
rect 15844 14424 15896 14433
rect 16580 14467 16632 14476
rect 16580 14433 16589 14467
rect 16589 14433 16623 14467
rect 16623 14433 16632 14467
rect 16580 14424 16632 14433
rect 15936 14356 15988 14408
rect 2504 14263 2556 14272
rect 2504 14229 2513 14263
rect 2513 14229 2547 14263
rect 2547 14229 2556 14263
rect 2504 14220 2556 14229
rect 3976 14263 4028 14272
rect 3976 14229 3985 14263
rect 3985 14229 4019 14263
rect 4019 14229 4028 14263
rect 3976 14220 4028 14229
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 5816 14220 5868 14272
rect 6736 14220 6788 14272
rect 8944 14263 8996 14272
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9680 14220 9732 14272
rect 10876 14220 10928 14272
rect 12808 14220 12860 14272
rect 17040 14288 17092 14340
rect 21088 14492 21140 14544
rect 17316 14424 17368 14476
rect 17592 14424 17644 14476
rect 18420 14356 18472 14408
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 17316 14288 17368 14340
rect 18144 14288 18196 14340
rect 18696 14288 18748 14340
rect 14924 14220 14976 14272
rect 15660 14220 15712 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 16948 14220 17000 14272
rect 17776 14220 17828 14272
rect 18788 14220 18840 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1676 14016 1728 14068
rect 5540 14016 5592 14068
rect 6552 14016 6604 14068
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 7012 14016 7064 14068
rect 9864 14059 9916 14068
rect 3056 13948 3108 14000
rect 3148 13948 3200 14000
rect 4160 13948 4212 14000
rect 4988 13948 5040 14000
rect 9220 13948 9272 14000
rect 4068 13855 4120 13864
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 3976 13744 4028 13796
rect 1952 13676 2004 13728
rect 5816 13880 5868 13932
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 7288 13880 7340 13932
rect 6828 13812 6880 13864
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 10324 14016 10376 14068
rect 11336 14016 11388 14068
rect 12900 14016 12952 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 17040 14016 17092 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 10048 13948 10100 14000
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 12072 13880 12124 13932
rect 9496 13812 9548 13864
rect 9588 13812 9640 13864
rect 9864 13812 9916 13864
rect 10600 13812 10652 13864
rect 10876 13855 10928 13864
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 11060 13812 11112 13864
rect 11796 13812 11848 13864
rect 7012 13744 7064 13796
rect 11244 13744 11296 13796
rect 11612 13744 11664 13796
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 16304 13948 16356 14000
rect 21088 14016 21140 14068
rect 19616 13948 19668 14000
rect 15384 13880 15436 13932
rect 15936 13923 15988 13932
rect 15936 13889 15954 13923
rect 15954 13889 15988 13923
rect 15936 13880 15988 13889
rect 16856 13880 16908 13932
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 19524 13880 19576 13932
rect 14004 13812 14056 13864
rect 14280 13812 14332 13864
rect 14556 13855 14608 13864
rect 14556 13821 14565 13855
rect 14565 13821 14599 13855
rect 14599 13821 14608 13855
rect 14556 13812 14608 13821
rect 14648 13744 14700 13796
rect 15200 13812 15252 13864
rect 17684 13855 17736 13864
rect 16396 13744 16448 13796
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 17776 13812 17828 13864
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 19064 13744 19116 13796
rect 19708 13812 19760 13864
rect 19800 13744 19852 13796
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 6368 13676 6420 13685
rect 8392 13676 8444 13728
rect 9128 13676 9180 13728
rect 9220 13676 9272 13728
rect 10968 13676 11020 13728
rect 12164 13676 12216 13728
rect 15844 13676 15896 13728
rect 16212 13676 16264 13728
rect 18512 13676 18564 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2320 13472 2372 13524
rect 4252 13472 4304 13524
rect 5448 13472 5500 13524
rect 5724 13472 5776 13524
rect 7380 13472 7432 13524
rect 12164 13472 12216 13524
rect 13728 13472 13780 13524
rect 15200 13472 15252 13524
rect 4068 13404 4120 13456
rect 1952 13336 2004 13388
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2596 13268 2648 13320
rect 4160 13336 4212 13388
rect 4344 13336 4396 13388
rect 5356 13336 5408 13388
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 6368 13336 6420 13388
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 6828 13336 6880 13388
rect 7748 13336 7800 13388
rect 10324 13404 10376 13456
rect 15936 13447 15988 13456
rect 9220 13336 9272 13388
rect 4528 13268 4580 13320
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 8208 13268 8260 13320
rect 9496 13268 9548 13320
rect 9588 13268 9640 13320
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13728 13336 13780 13388
rect 15936 13413 15945 13447
rect 15945 13413 15979 13447
rect 15979 13413 15988 13447
rect 15936 13404 15988 13413
rect 16396 13472 16448 13524
rect 16948 13472 17000 13524
rect 18880 13472 18932 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 16856 13447 16908 13456
rect 16856 13413 16865 13447
rect 16865 13413 16899 13447
rect 16899 13413 16908 13447
rect 16856 13404 16908 13413
rect 18972 13404 19024 13456
rect 11152 13268 11204 13320
rect 13360 13268 13412 13320
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 16948 13336 17000 13388
rect 17592 13336 17644 13388
rect 3148 13200 3200 13252
rect 3332 13243 3384 13252
rect 3332 13209 3372 13243
rect 3372 13209 3384 13243
rect 3332 13200 3384 13209
rect 4160 13200 4212 13252
rect 7380 13243 7432 13252
rect 3056 13132 3108 13184
rect 3240 13132 3292 13184
rect 4344 13132 4396 13184
rect 4620 13132 4672 13184
rect 5448 13132 5500 13184
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 5816 13132 5868 13184
rect 6644 13132 6696 13184
rect 7380 13209 7389 13243
rect 7389 13209 7423 13243
rect 7423 13209 7432 13243
rect 7380 13200 7432 13209
rect 7932 13132 7984 13184
rect 9036 13132 9088 13184
rect 10600 13200 10652 13252
rect 10692 13132 10744 13184
rect 13820 13200 13872 13252
rect 17040 13268 17092 13320
rect 18788 13268 18840 13320
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 14648 13200 14700 13252
rect 15200 13200 15252 13252
rect 15844 13200 15896 13252
rect 17776 13200 17828 13252
rect 17868 13200 17920 13252
rect 11152 13132 11204 13184
rect 12348 13132 12400 13184
rect 14740 13132 14792 13184
rect 19984 13200 20036 13252
rect 18972 13132 19024 13184
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 20168 13132 20220 13184
rect 20444 13175 20496 13184
rect 20444 13141 20453 13175
rect 20453 13141 20487 13175
rect 20487 13141 20496 13175
rect 20444 13132 20496 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 3056 12928 3108 12980
rect 3976 12928 4028 12980
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 1952 12860 2004 12912
rect 4712 12860 4764 12912
rect 6000 12860 6052 12912
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 4068 12792 4120 12844
rect 4896 12792 4948 12844
rect 5356 12792 5408 12844
rect 7288 12928 7340 12980
rect 7472 12928 7524 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 9128 12971 9180 12980
rect 4252 12724 4304 12776
rect 5724 12724 5776 12776
rect 6000 12724 6052 12776
rect 6828 12860 6880 12912
rect 7012 12860 7064 12912
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 12532 12928 12584 12980
rect 13728 12928 13780 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 17040 12928 17092 12980
rect 17960 12928 18012 12980
rect 19432 12928 19484 12980
rect 19524 12928 19576 12980
rect 19800 12928 19852 12980
rect 20444 12928 20496 12980
rect 6644 12835 6696 12844
rect 6644 12801 6667 12835
rect 6667 12801 6696 12835
rect 6644 12792 6696 12801
rect 7748 12792 7800 12844
rect 7840 12724 7892 12776
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 3884 12588 3936 12640
rect 4252 12588 4304 12640
rect 5080 12588 5132 12640
rect 5448 12588 5500 12640
rect 6736 12588 6788 12640
rect 9496 12792 9548 12844
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 9588 12724 9640 12776
rect 10140 12724 10192 12776
rect 10692 12656 10744 12708
rect 9036 12588 9088 12640
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 11152 12792 11204 12844
rect 12348 12792 12400 12844
rect 14648 12860 14700 12912
rect 14740 12792 14792 12844
rect 14832 12792 14884 12844
rect 15936 12860 15988 12912
rect 16948 12860 17000 12912
rect 17132 12903 17184 12912
rect 17132 12869 17141 12903
rect 17141 12869 17175 12903
rect 17175 12869 17184 12903
rect 17132 12860 17184 12869
rect 17224 12860 17276 12912
rect 13544 12656 13596 12708
rect 17040 12792 17092 12844
rect 18972 12860 19024 12912
rect 20536 12860 20588 12912
rect 21272 12860 21324 12912
rect 18236 12792 18288 12844
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 18052 12724 18104 12776
rect 16212 12656 16264 12708
rect 12992 12588 13044 12640
rect 13452 12588 13504 12640
rect 15200 12588 15252 12640
rect 15568 12588 15620 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 17224 12588 17276 12640
rect 17592 12588 17644 12640
rect 17960 12588 18012 12640
rect 18328 12588 18380 12640
rect 18696 12588 18748 12640
rect 19064 12588 19116 12640
rect 20904 12588 20956 12640
rect 22376 12588 22428 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 1860 12384 1912 12436
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 3148 12384 3200 12436
rect 4804 12384 4856 12436
rect 6000 12384 6052 12436
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 7656 12384 7708 12436
rect 2504 12316 2556 12368
rect 3332 12248 3384 12300
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 3240 12223 3292 12232
rect 2228 12180 2280 12189
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3884 12316 3936 12368
rect 3976 12316 4028 12368
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 6644 12316 6696 12368
rect 4528 12248 4580 12300
rect 9956 12316 10008 12368
rect 12348 12384 12400 12436
rect 12992 12384 13044 12436
rect 15292 12316 15344 12368
rect 15752 12316 15804 12368
rect 16304 12384 16356 12436
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 19708 12384 19760 12436
rect 20628 12384 20680 12436
rect 20444 12316 20496 12368
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 8208 12248 8260 12300
rect 8300 12248 8352 12300
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 13728 12248 13780 12300
rect 14188 12291 14240 12300
rect 14188 12257 14197 12291
rect 14197 12257 14231 12291
rect 14231 12257 14240 12291
rect 14188 12248 14240 12257
rect 14648 12248 14700 12300
rect 15200 12248 15252 12300
rect 16948 12291 17000 12300
rect 3332 12112 3384 12164
rect 2412 12044 2464 12096
rect 6552 12180 6604 12232
rect 7288 12180 7340 12232
rect 11152 12180 11204 12232
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 5540 12112 5592 12164
rect 6920 12112 6972 12164
rect 7748 12112 7800 12164
rect 12164 12112 12216 12164
rect 14556 12180 14608 12232
rect 15752 12180 15804 12232
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 18144 12248 18196 12300
rect 18788 12248 18840 12300
rect 19984 12248 20036 12300
rect 20720 12248 20772 12300
rect 16672 12180 16724 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 4252 12044 4304 12096
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7012 12044 7064 12096
rect 9404 12044 9456 12096
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 11060 12044 11112 12096
rect 11152 12044 11204 12096
rect 12256 12044 12308 12096
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 16764 12155 16816 12164
rect 15292 12044 15344 12096
rect 16764 12121 16773 12155
rect 16773 12121 16807 12155
rect 16807 12121 16816 12155
rect 16764 12112 16816 12121
rect 17224 12112 17276 12164
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 17776 12044 17828 12096
rect 18604 12044 18656 12096
rect 19064 12044 19116 12096
rect 21364 12044 21416 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2228 11840 2280 11892
rect 4712 11883 4764 11892
rect 2504 11772 2556 11824
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 4804 11840 4856 11892
rect 5448 11840 5500 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 3240 11772 3292 11824
rect 4068 11772 4120 11824
rect 4252 11772 4304 11824
rect 4528 11772 4580 11824
rect 4896 11815 4948 11824
rect 4896 11781 4905 11815
rect 4905 11781 4939 11815
rect 4939 11781 4948 11815
rect 4896 11772 4948 11781
rect 8668 11840 8720 11892
rect 11244 11840 11296 11892
rect 11428 11840 11480 11892
rect 8300 11772 8352 11824
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 4712 11704 4764 11756
rect 4988 11704 5040 11756
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 8576 11747 8628 11756
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2964 11679 3016 11688
rect 2780 11636 2832 11645
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 6552 11636 6604 11688
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 3976 11568 4028 11620
rect 5080 11500 5132 11552
rect 6736 11568 6788 11620
rect 6920 11568 6972 11620
rect 7932 11500 7984 11552
rect 9772 11704 9824 11756
rect 10508 11704 10560 11756
rect 12164 11840 12216 11892
rect 14740 11840 14792 11892
rect 15752 11840 15804 11892
rect 16028 11840 16080 11892
rect 17776 11840 17828 11892
rect 18972 11840 19024 11892
rect 12808 11815 12860 11824
rect 12808 11781 12817 11815
rect 12817 11781 12851 11815
rect 12851 11781 12860 11815
rect 12808 11772 12860 11781
rect 13452 11772 13504 11824
rect 13820 11772 13872 11824
rect 17500 11772 17552 11824
rect 17960 11772 18012 11824
rect 11520 11704 11572 11756
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 12256 11704 12308 11756
rect 12532 11704 12584 11756
rect 14188 11747 14240 11756
rect 11060 11568 11112 11620
rect 11336 11611 11388 11620
rect 11336 11577 11345 11611
rect 11345 11577 11379 11611
rect 11379 11577 11388 11611
rect 13176 11636 13228 11688
rect 13452 11636 13504 11688
rect 11336 11568 11388 11577
rect 9312 11500 9364 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 14464 11747 14516 11756
rect 14464 11713 14498 11747
rect 14498 11713 14516 11747
rect 14464 11704 14516 11713
rect 15568 11704 15620 11756
rect 16212 11704 16264 11756
rect 21180 11772 21232 11824
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 19616 11704 19668 11756
rect 16304 11679 16356 11688
rect 16304 11645 16313 11679
rect 16313 11645 16347 11679
rect 16347 11645 16356 11679
rect 16304 11636 16356 11645
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 17776 11679 17828 11688
rect 16856 11568 16908 11620
rect 17776 11645 17785 11679
rect 17785 11645 17819 11679
rect 17819 11645 17828 11679
rect 17776 11636 17828 11645
rect 17868 11568 17920 11620
rect 17960 11568 18012 11620
rect 15568 11500 15620 11552
rect 15844 11500 15896 11552
rect 17316 11500 17368 11552
rect 18052 11500 18104 11552
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 18972 11500 19024 11552
rect 21364 11704 21416 11756
rect 22100 11704 22152 11756
rect 21640 11636 21692 11688
rect 21180 11568 21232 11620
rect 21272 11568 21324 11620
rect 20444 11543 20496 11552
rect 20444 11509 20453 11543
rect 20453 11509 20487 11543
rect 20487 11509 20496 11543
rect 20444 11500 20496 11509
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2964 11296 3016 11348
rect 3516 11296 3568 11348
rect 4252 11296 4304 11348
rect 2872 11228 2924 11280
rect 5264 11296 5316 11348
rect 5540 11296 5592 11348
rect 5816 11296 5868 11348
rect 8208 11296 8260 11348
rect 9404 11296 9456 11348
rect 3884 11160 3936 11212
rect 1492 11092 1544 11144
rect 3516 11092 3568 11144
rect 4252 11092 4304 11144
rect 2596 11024 2648 11076
rect 6552 11160 6604 11212
rect 8576 11160 8628 11212
rect 4528 11024 4580 11076
rect 5264 11024 5316 11076
rect 6000 10956 6052 11008
rect 7012 10956 7064 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7472 11024 7524 11076
rect 8024 11024 8076 11076
rect 8668 11092 8720 11144
rect 9220 11092 9272 11144
rect 11428 11296 11480 11348
rect 13820 11296 13872 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16304 11296 16356 11348
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 18604 11339 18656 11348
rect 18604 11305 18613 11339
rect 18613 11305 18647 11339
rect 18647 11305 18656 11339
rect 18604 11296 18656 11305
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 11888 11160 11940 11212
rect 12256 11228 12308 11280
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13820 11203 13872 11212
rect 13452 11160 13504 11169
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 15568 11228 15620 11280
rect 15844 11203 15896 11212
rect 15844 11169 15853 11203
rect 15853 11169 15887 11203
rect 15887 11169 15896 11203
rect 15844 11160 15896 11169
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 11060 11092 11112 11144
rect 9956 11024 10008 11076
rect 10784 11024 10836 11076
rect 12256 11024 12308 11076
rect 12624 11092 12676 11144
rect 16120 11092 16172 11144
rect 17040 11092 17092 11144
rect 17316 11228 17368 11280
rect 18144 11160 18196 11212
rect 17960 11092 18012 11144
rect 19892 11296 19944 11348
rect 20536 11296 20588 11348
rect 14556 11024 14608 11076
rect 15108 11024 15160 11076
rect 16948 11024 17000 11076
rect 19064 11024 19116 11076
rect 19156 11024 19208 11076
rect 19708 11024 19760 11076
rect 20444 11024 20496 11076
rect 21088 11092 21140 11144
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 21640 11024 21692 11076
rect 22192 11024 22244 11076
rect 7196 10956 7248 10965
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 10140 10956 10192 11008
rect 10508 10999 10560 11008
rect 10508 10965 10517 10999
rect 10517 10965 10551 10999
rect 10551 10965 10560 10999
rect 10508 10956 10560 10965
rect 10600 10999 10652 11008
rect 10600 10965 10609 10999
rect 10609 10965 10643 10999
rect 10643 10965 10652 10999
rect 10600 10956 10652 10965
rect 11704 10956 11756 11008
rect 11980 10999 12032 11008
rect 11980 10965 11989 10999
rect 11989 10965 12023 10999
rect 12023 10965 12032 10999
rect 11980 10956 12032 10965
rect 12900 10999 12952 11008
rect 12900 10965 12909 10999
rect 12909 10965 12943 10999
rect 12943 10965 12952 10999
rect 13268 10999 13320 11008
rect 12900 10956 12952 10965
rect 13268 10965 13277 10999
rect 13277 10965 13311 10999
rect 13311 10965 13320 10999
rect 13268 10956 13320 10965
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 15384 10956 15436 11008
rect 15844 10956 15896 11008
rect 15936 10956 15988 11008
rect 16396 10956 16448 11008
rect 17684 10956 17736 11008
rect 17960 10956 18012 11008
rect 18972 10956 19024 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2964 10684 3016 10736
rect 1492 10616 1544 10668
rect 1676 10659 1728 10668
rect 1676 10625 1710 10659
rect 1710 10625 1728 10659
rect 1676 10616 1728 10625
rect 3516 10616 3568 10668
rect 4528 10752 4580 10804
rect 6552 10752 6604 10804
rect 7196 10752 7248 10804
rect 5080 10684 5132 10736
rect 5356 10684 5408 10736
rect 6000 10684 6052 10736
rect 6460 10684 6512 10736
rect 9220 10752 9272 10804
rect 4252 10548 4304 10600
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 5724 10480 5776 10532
rect 6460 10548 6512 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 2596 10412 2648 10464
rect 4068 10412 4120 10464
rect 7472 10480 7524 10532
rect 8300 10616 8352 10668
rect 8024 10548 8076 10600
rect 9404 10684 9456 10736
rect 9588 10684 9640 10736
rect 8576 10616 8628 10668
rect 9772 10752 9824 10804
rect 10600 10752 10652 10804
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 12808 10752 12860 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 14372 10752 14424 10804
rect 14924 10752 14976 10804
rect 10324 10727 10376 10736
rect 10324 10693 10333 10727
rect 10333 10693 10367 10727
rect 10367 10693 10376 10727
rect 10324 10684 10376 10693
rect 11796 10684 11848 10736
rect 13452 10684 13504 10736
rect 16212 10752 16264 10804
rect 16396 10752 16448 10804
rect 16672 10752 16724 10804
rect 19616 10752 19668 10804
rect 20168 10752 20220 10804
rect 21272 10795 21324 10804
rect 21272 10761 21281 10795
rect 21281 10761 21315 10795
rect 21315 10761 21324 10795
rect 21272 10752 21324 10761
rect 10968 10616 11020 10668
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 15660 10684 15712 10736
rect 7656 10412 7708 10464
rect 8392 10412 8444 10464
rect 8668 10412 8720 10464
rect 10600 10548 10652 10600
rect 11336 10548 11388 10600
rect 13360 10548 13412 10600
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 15016 10548 15068 10600
rect 17316 10616 17368 10668
rect 19156 10684 19208 10736
rect 18604 10616 18656 10668
rect 20076 10616 20128 10668
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 14464 10480 14516 10532
rect 16212 10480 16264 10532
rect 9588 10412 9640 10464
rect 9772 10412 9824 10464
rect 9956 10412 10008 10464
rect 10324 10412 10376 10464
rect 10784 10412 10836 10464
rect 11704 10412 11756 10464
rect 12072 10412 12124 10464
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 16948 10480 17000 10532
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 20812 10591 20864 10600
rect 17316 10480 17368 10532
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18972 10480 19024 10532
rect 19156 10480 19208 10532
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 21640 10480 21692 10532
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2688 10208 2740 10260
rect 2780 10208 2832 10260
rect 3884 10208 3936 10260
rect 2596 10072 2648 10124
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 5540 10140 5592 10192
rect 6644 10208 6696 10260
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 9036 10208 9088 10260
rect 9220 10208 9272 10260
rect 9312 10208 9364 10260
rect 11704 10208 11756 10260
rect 13268 10208 13320 10260
rect 13360 10208 13412 10260
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 16672 10208 16724 10260
rect 18144 10208 18196 10260
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20812 10208 20864 10260
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 4344 10004 4396 10056
rect 5908 10004 5960 10056
rect 6000 10004 6052 10056
rect 7012 10140 7064 10192
rect 8208 10140 8260 10192
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 8576 10115 8628 10124
rect 8576 10081 8585 10115
rect 8585 10081 8619 10115
rect 8619 10081 8628 10115
rect 8576 10072 8628 10081
rect 10140 10140 10192 10192
rect 10784 10183 10836 10192
rect 10784 10149 10793 10183
rect 10793 10149 10827 10183
rect 10827 10149 10836 10183
rect 10784 10140 10836 10149
rect 10968 10140 11020 10192
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 9772 10072 9824 10124
rect 10324 10072 10376 10124
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 11336 10072 11388 10124
rect 11888 10115 11940 10124
rect 4528 9936 4580 9988
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 2136 9911 2188 9920
rect 2136 9877 2145 9911
rect 2145 9877 2179 9911
rect 2179 9877 2188 9911
rect 2136 9868 2188 9877
rect 3056 9868 3108 9920
rect 6920 9936 6972 9988
rect 7564 9936 7616 9988
rect 9036 9936 9088 9988
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 8392 9911 8444 9920
rect 7288 9868 7340 9877
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 10048 10004 10100 10056
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 11980 10072 12032 10124
rect 12164 10004 12216 10056
rect 13636 10140 13688 10192
rect 16764 10140 16816 10192
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 14188 10115 14240 10124
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 14188 10072 14240 10081
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 13176 10004 13228 10056
rect 13544 10004 13596 10056
rect 16212 10072 16264 10124
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 19616 10072 19668 10124
rect 20444 10140 20496 10192
rect 16764 10004 16816 10056
rect 14924 9936 14976 9988
rect 17132 10004 17184 10056
rect 17316 10004 17368 10056
rect 18236 10004 18288 10056
rect 17500 9979 17552 9988
rect 17500 9945 17512 9979
rect 17512 9945 17552 9979
rect 17500 9936 17552 9945
rect 17776 9936 17828 9988
rect 20812 9936 20864 9988
rect 8484 9868 8536 9877
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 13268 9868 13320 9920
rect 13820 9868 13872 9920
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 14740 9868 14792 9920
rect 16672 9868 16724 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 20904 9868 20956 9920
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 21640 9868 21692 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 2044 9664 2096 9716
rect 2596 9596 2648 9648
rect 2044 9528 2096 9580
rect 4436 9664 4488 9716
rect 4528 9664 4580 9716
rect 5080 9707 5132 9716
rect 5080 9673 5089 9707
rect 5089 9673 5123 9707
rect 5123 9673 5132 9707
rect 5080 9664 5132 9673
rect 5540 9664 5592 9716
rect 5724 9664 5776 9716
rect 2228 9503 2280 9512
rect 2228 9469 2237 9503
rect 2237 9469 2271 9503
rect 2271 9469 2280 9503
rect 2228 9460 2280 9469
rect 1676 9392 1728 9444
rect 6000 9596 6052 9648
rect 6552 9596 6604 9648
rect 8300 9707 8352 9716
rect 8300 9673 8309 9707
rect 8309 9673 8343 9707
rect 8343 9673 8352 9707
rect 8300 9664 8352 9673
rect 8576 9664 8628 9716
rect 10600 9664 10652 9716
rect 10784 9664 10836 9716
rect 11704 9664 11756 9716
rect 13452 9664 13504 9716
rect 4988 9392 5040 9444
rect 7012 9528 7064 9580
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 7380 9460 7432 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 8668 9639 8720 9648
rect 8668 9605 8702 9639
rect 8702 9605 8720 9639
rect 10416 9639 10468 9648
rect 8668 9596 8720 9605
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 14188 9664 14240 9716
rect 16304 9664 16356 9716
rect 8024 9528 8076 9580
rect 7472 9460 7524 9469
rect 8300 9460 8352 9512
rect 3976 9367 4028 9376
rect 3976 9333 3985 9367
rect 3985 9333 4019 9367
rect 4019 9333 4028 9367
rect 3976 9324 4028 9333
rect 4436 9324 4488 9376
rect 4896 9324 4948 9376
rect 5080 9324 5132 9376
rect 6920 9324 6972 9376
rect 7748 9324 7800 9376
rect 11888 9571 11940 9580
rect 10508 9460 10560 9512
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 13636 9596 13688 9648
rect 14924 9639 14976 9648
rect 14924 9605 14933 9639
rect 14933 9605 14967 9639
rect 14967 9605 14976 9639
rect 14924 9596 14976 9605
rect 16488 9634 16540 9686
rect 16856 9664 16908 9716
rect 17960 9664 18012 9716
rect 18696 9664 18748 9716
rect 18972 9664 19024 9716
rect 19708 9664 19760 9716
rect 20812 9664 20864 9716
rect 16580 9596 16632 9648
rect 17040 9596 17092 9648
rect 17224 9596 17276 9648
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 14556 9528 14608 9580
rect 9404 9324 9456 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 11704 9392 11756 9444
rect 12348 9392 12400 9444
rect 12256 9324 12308 9376
rect 13360 9460 13412 9512
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 15660 9460 15712 9512
rect 15292 9392 15344 9444
rect 15016 9324 15068 9376
rect 15200 9324 15252 9376
rect 15476 9324 15528 9376
rect 16028 9324 16080 9376
rect 16304 9324 16356 9376
rect 17500 9528 17552 9580
rect 17868 9596 17920 9648
rect 19524 9639 19576 9648
rect 19524 9605 19542 9639
rect 19542 9605 19576 9639
rect 19524 9596 19576 9605
rect 20260 9571 20312 9580
rect 16488 9460 16540 9512
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 17868 9460 17920 9512
rect 20444 9503 20496 9512
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 16764 9324 16816 9376
rect 18696 9392 18748 9444
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 18512 9324 18564 9376
rect 20444 9469 20453 9503
rect 20453 9469 20487 9503
rect 20487 9469 20496 9503
rect 20444 9460 20496 9469
rect 21180 9596 21232 9648
rect 20628 9528 20680 9580
rect 20812 9460 20864 9512
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2228 9120 2280 9172
rect 4344 9120 4396 9172
rect 5816 9120 5868 9172
rect 6092 9163 6144 9172
rect 3424 9052 3476 9104
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 7012 9120 7064 9172
rect 7288 9163 7340 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 2596 8916 2648 8968
rect 3332 9027 3384 9036
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 3332 8984 3384 8993
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 1584 8848 1636 8900
rect 2872 8848 2924 8900
rect 3240 8848 3292 8900
rect 3516 8848 3568 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2136 8780 2188 8832
rect 4344 8984 4396 9036
rect 4804 8984 4856 9036
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5080 8984 5132 9036
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 6460 9052 6512 9104
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 8024 9120 8076 9172
rect 8392 9120 8444 9172
rect 9128 9120 9180 9172
rect 10508 9163 10560 9172
rect 10508 9129 10517 9163
rect 10517 9129 10551 9163
rect 10551 9129 10560 9163
rect 10508 9120 10560 9129
rect 8668 9052 8720 9104
rect 9680 9052 9732 9104
rect 11980 9120 12032 9172
rect 12256 9163 12308 9172
rect 12256 9129 12265 9163
rect 12265 9129 12299 9163
rect 12299 9129 12308 9163
rect 12256 9120 12308 9129
rect 12808 9120 12860 9172
rect 14372 9120 14424 9172
rect 11888 9052 11940 9104
rect 5908 8984 5960 9036
rect 6552 8984 6604 9036
rect 7288 8984 7340 9036
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 3976 8916 4028 8968
rect 4436 8916 4488 8968
rect 6828 8916 6880 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 4620 8848 4672 8900
rect 5080 8848 5132 8900
rect 5356 8848 5408 8900
rect 8208 8848 8260 8900
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 4988 8780 5040 8832
rect 5724 8780 5776 8832
rect 6460 8780 6512 8832
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 8392 8780 8444 8832
rect 13176 9052 13228 9104
rect 17960 9120 18012 9172
rect 20720 9163 20772 9172
rect 12992 9027 13044 9036
rect 11152 8916 11204 8968
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 13084 8984 13136 9036
rect 14556 8984 14608 9036
rect 15108 9027 15160 9036
rect 14648 8916 14700 8968
rect 8668 8848 8720 8900
rect 9772 8848 9824 8900
rect 12164 8848 12216 8900
rect 12532 8848 12584 8900
rect 15108 8993 15117 9027
rect 15117 8993 15151 9027
rect 15151 8993 15160 9027
rect 15108 8984 15160 8993
rect 16764 8959 16816 8968
rect 11796 8780 11848 8832
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 13360 8780 13412 8832
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 14464 8780 14516 8832
rect 15476 8848 15528 8900
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 17776 8984 17828 9036
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 20812 9052 20864 9104
rect 18512 8916 18564 8968
rect 18696 8916 18748 8968
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 20444 8984 20496 9036
rect 19892 8916 19944 8968
rect 21364 8916 21416 8968
rect 15936 8780 15988 8832
rect 16580 8780 16632 8832
rect 18420 8848 18472 8900
rect 17224 8780 17276 8832
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1768 8576 1820 8628
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 4528 8619 4580 8628
rect 2504 8576 2556 8585
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 4804 8576 4856 8628
rect 5356 8576 5408 8628
rect 5816 8576 5868 8628
rect 1860 8508 1912 8560
rect 2596 8508 2648 8560
rect 2872 8440 2924 8492
rect 3240 8483 3292 8492
rect 3240 8449 3274 8483
rect 3274 8449 3292 8483
rect 3240 8440 3292 8449
rect 4160 8440 4212 8492
rect 4620 8440 4672 8492
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 1676 8372 1728 8424
rect 2504 8372 2556 8424
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 1216 8304 1268 8356
rect 2780 8304 2832 8356
rect 2136 8236 2188 8288
rect 4528 8372 4580 8424
rect 5356 8372 5408 8424
rect 6000 8508 6052 8560
rect 8484 8576 8536 8628
rect 9128 8576 9180 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 5724 8440 5776 8492
rect 6276 8440 6328 8492
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 4068 8304 4120 8356
rect 4804 8304 4856 8356
rect 6552 8304 6604 8356
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 9496 8508 9548 8560
rect 10508 8508 10560 8560
rect 8208 8440 8260 8492
rect 11060 8440 11112 8492
rect 12992 8576 13044 8628
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 14280 8576 14332 8628
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 18696 8576 18748 8628
rect 20076 8576 20128 8628
rect 20536 8576 20588 8628
rect 21732 8576 21784 8628
rect 11704 8508 11756 8560
rect 13360 8508 13412 8560
rect 12256 8483 12308 8492
rect 9588 8415 9640 8424
rect 7012 8236 7064 8288
rect 7380 8236 7432 8288
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 8484 8236 8536 8288
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 12900 8440 12952 8492
rect 12164 8372 12216 8424
rect 13728 8440 13780 8492
rect 13544 8372 13596 8424
rect 15476 8508 15528 8560
rect 16120 8483 16172 8492
rect 13728 8304 13780 8356
rect 14556 8304 14608 8356
rect 9404 8236 9456 8288
rect 11152 8236 11204 8288
rect 11796 8236 11848 8288
rect 11980 8236 12032 8288
rect 12808 8236 12860 8288
rect 12992 8279 13044 8288
rect 12992 8245 13001 8279
rect 13001 8245 13035 8279
rect 13035 8245 13044 8279
rect 12992 8236 13044 8245
rect 13084 8236 13136 8288
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 14648 8236 14700 8288
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16948 8440 17000 8492
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 15936 8415 15988 8424
rect 15936 8381 15945 8415
rect 15945 8381 15979 8415
rect 15979 8381 15988 8415
rect 15936 8372 15988 8381
rect 17224 8372 17276 8424
rect 17684 8372 17736 8424
rect 18512 8440 18564 8492
rect 21364 8508 21416 8560
rect 19524 8483 19576 8492
rect 19524 8449 19542 8483
rect 19542 8449 19576 8483
rect 19524 8440 19576 8449
rect 19708 8440 19760 8492
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 22284 8372 22336 8424
rect 17132 8304 17184 8356
rect 17316 8304 17368 8356
rect 19892 8347 19944 8356
rect 19892 8313 19901 8347
rect 19901 8313 19935 8347
rect 19935 8313 19944 8347
rect 19892 8304 19944 8313
rect 20076 8304 20128 8356
rect 21640 8304 21692 8356
rect 15108 8236 15160 8288
rect 15660 8236 15712 8288
rect 16212 8236 16264 8288
rect 18788 8236 18840 8288
rect 19432 8236 19484 8288
rect 19616 8236 19668 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 6368 8032 6420 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 3240 7964 3292 8016
rect 6276 7964 6328 8016
rect 6828 8032 6880 8084
rect 6920 8032 6972 8084
rect 7380 8007 7432 8016
rect 2228 7939 2280 7948
rect 2228 7905 2237 7939
rect 2237 7905 2271 7939
rect 2271 7905 2280 7939
rect 2228 7896 2280 7905
rect 4160 7896 4212 7948
rect 4896 7939 4948 7948
rect 4896 7905 4905 7939
rect 4905 7905 4939 7939
rect 4939 7905 4948 7939
rect 4896 7896 4948 7905
rect 7380 7973 7389 8007
rect 7389 7973 7423 8007
rect 7423 7973 7432 8007
rect 7380 7964 7432 7973
rect 2964 7828 3016 7880
rect 4436 7828 4488 7880
rect 3056 7760 3108 7812
rect 4988 7828 5040 7880
rect 1768 7692 1820 7744
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 2504 7692 2556 7744
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 3608 7692 3660 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 5080 7692 5132 7744
rect 5356 7760 5408 7812
rect 5724 7760 5776 7812
rect 6736 7760 6788 7812
rect 6920 7896 6972 7948
rect 7288 7896 7340 7948
rect 8300 8032 8352 8084
rect 7748 7964 7800 8016
rect 10692 7964 10744 8016
rect 12164 8032 12216 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 13452 8032 13504 8084
rect 11704 7964 11756 8016
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 9588 7939 9640 7948
rect 9588 7905 9597 7939
rect 9597 7905 9631 7939
rect 9631 7905 9640 7939
rect 9588 7896 9640 7905
rect 9772 7896 9824 7948
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8484 7828 8536 7880
rect 10600 7828 10652 7880
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8208 7692 8260 7744
rect 10968 7896 11020 7948
rect 11796 7828 11848 7880
rect 12900 7896 12952 7948
rect 14740 8032 14792 8084
rect 14832 8032 14884 8084
rect 16120 8032 16172 8084
rect 17684 7964 17736 8016
rect 19524 8032 19576 8084
rect 20260 8032 20312 8084
rect 15660 7896 15712 7948
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 16396 7896 16448 7948
rect 20444 7939 20496 7948
rect 9864 7692 9916 7744
rect 10324 7692 10376 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 13728 7760 13780 7812
rect 15016 7760 15068 7812
rect 17316 7828 17368 7880
rect 20444 7905 20453 7939
rect 20453 7905 20487 7939
rect 20487 7905 20496 7939
rect 20444 7896 20496 7905
rect 20720 7896 20772 7948
rect 21364 7939 21416 7948
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 18512 7828 18564 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20904 7828 20956 7880
rect 12992 7692 13044 7744
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 15476 7735 15528 7744
rect 13360 7692 13412 7701
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 15568 7735 15620 7744
rect 15568 7701 15577 7735
rect 15577 7701 15611 7735
rect 15611 7701 15620 7735
rect 15568 7692 15620 7701
rect 15844 7692 15896 7744
rect 17224 7692 17276 7744
rect 18880 7760 18932 7812
rect 21088 7760 21140 7812
rect 18144 7692 18196 7744
rect 19340 7735 19392 7744
rect 19340 7701 19349 7735
rect 19349 7701 19383 7735
rect 19383 7701 19392 7735
rect 19340 7692 19392 7701
rect 19616 7692 19668 7744
rect 20904 7692 20956 7744
rect 21272 7828 21324 7880
rect 21364 7760 21416 7812
rect 21732 7760 21784 7812
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 21640 7692 21692 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 2780 7488 2832 7540
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3608 7488 3660 7497
rect 4712 7488 4764 7540
rect 1492 7420 1544 7472
rect 2136 7420 2188 7472
rect 2504 7463 2556 7472
rect 2504 7429 2513 7463
rect 2513 7429 2547 7463
rect 2547 7429 2556 7463
rect 2504 7420 2556 7429
rect 4252 7420 4304 7472
rect 4436 7420 4488 7472
rect 4896 7420 4948 7472
rect 4988 7420 5040 7472
rect 5816 7463 5868 7472
rect 5816 7429 5825 7463
rect 5825 7429 5859 7463
rect 5859 7429 5868 7463
rect 5816 7420 5868 7429
rect 2872 7352 2924 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 2596 7327 2648 7336
rect 2596 7293 2605 7327
rect 2605 7293 2639 7327
rect 2639 7293 2648 7327
rect 2596 7284 2648 7293
rect 2412 7216 2464 7268
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 7380 7420 7432 7472
rect 5908 7327 5960 7336
rect 5908 7293 5917 7327
rect 5917 7293 5951 7327
rect 5951 7293 5960 7327
rect 5908 7284 5960 7293
rect 3424 7216 3476 7268
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 2596 7148 2648 7200
rect 4160 7148 4212 7200
rect 4804 7148 4856 7200
rect 7564 7352 7616 7404
rect 8576 7420 8628 7472
rect 8668 7352 8720 7404
rect 9404 7352 9456 7404
rect 9864 7463 9916 7472
rect 9864 7429 9873 7463
rect 9873 7429 9907 7463
rect 9907 7429 9916 7463
rect 9864 7420 9916 7429
rect 10232 7488 10284 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 10968 7488 11020 7540
rect 12256 7488 12308 7540
rect 12808 7488 12860 7540
rect 10324 7463 10376 7472
rect 10324 7429 10333 7463
rect 10333 7429 10367 7463
rect 10367 7429 10376 7463
rect 10324 7420 10376 7429
rect 11152 7420 11204 7472
rect 11244 7420 11296 7472
rect 15292 7488 15344 7540
rect 15568 7488 15620 7540
rect 15660 7488 15712 7540
rect 16212 7488 16264 7540
rect 17224 7488 17276 7540
rect 18604 7488 18656 7540
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 20536 7488 20588 7540
rect 21180 7531 21232 7540
rect 10968 7352 11020 7404
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12992 7352 13044 7404
rect 17960 7420 18012 7472
rect 15108 7352 15160 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 17500 7352 17552 7404
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 9128 7216 9180 7268
rect 12532 7216 12584 7268
rect 12624 7216 12676 7268
rect 12992 7216 13044 7268
rect 14464 7284 14516 7336
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 15476 7284 15528 7336
rect 16948 7327 17000 7336
rect 14740 7216 14792 7268
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 17776 7284 17828 7336
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 19524 7420 19576 7472
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 19156 7352 19208 7404
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 20904 7352 20956 7404
rect 21088 7352 21140 7404
rect 6736 7148 6788 7200
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 10968 7191 11020 7200
rect 9496 7148 9548 7157
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 11888 7148 11940 7200
rect 12164 7148 12216 7200
rect 13176 7148 13228 7200
rect 13728 7191 13780 7200
rect 13728 7157 13737 7191
rect 13737 7157 13771 7191
rect 13771 7157 13780 7191
rect 13728 7148 13780 7157
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 17316 7148 17368 7200
rect 18604 7191 18656 7200
rect 18604 7157 18613 7191
rect 18613 7157 18647 7191
rect 18647 7157 18656 7191
rect 18604 7148 18656 7157
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 20720 7284 20772 7336
rect 21364 7216 21416 7268
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2228 6944 2280 6996
rect 2872 6944 2924 6996
rect 3056 6987 3108 6996
rect 3056 6953 3065 6987
rect 3065 6953 3099 6987
rect 3099 6953 3108 6987
rect 3056 6944 3108 6953
rect 3792 6944 3844 6996
rect 4068 6944 4120 6996
rect 9128 6944 9180 6996
rect 11980 6944 12032 6996
rect 12532 6944 12584 6996
rect 14832 6944 14884 6996
rect 15568 6944 15620 6996
rect 18880 6987 18932 6996
rect 18880 6953 18889 6987
rect 18889 6953 18923 6987
rect 18923 6953 18932 6987
rect 18880 6944 18932 6953
rect 19064 6944 19116 6996
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 3516 6808 3568 6860
rect 3792 6851 3844 6860
rect 3792 6817 3801 6851
rect 3801 6817 3835 6851
rect 3835 6817 3844 6851
rect 3792 6808 3844 6817
rect 4436 6740 4488 6792
rect 4988 6808 5040 6860
rect 5264 6808 5316 6860
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 5908 6876 5960 6928
rect 7196 6876 7248 6928
rect 7564 6876 7616 6928
rect 9588 6919 9640 6928
rect 9588 6885 9597 6919
rect 9597 6885 9631 6919
rect 9631 6885 9640 6919
rect 9588 6876 9640 6885
rect 11060 6876 11112 6928
rect 13636 6876 13688 6928
rect 13820 6876 13872 6928
rect 15292 6876 15344 6928
rect 2136 6672 2188 6724
rect 2228 6604 2280 6656
rect 3700 6672 3752 6724
rect 3056 6604 3108 6656
rect 4712 6604 4764 6656
rect 5356 6740 5408 6792
rect 6828 6808 6880 6860
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 5080 6672 5132 6724
rect 7012 6740 7064 6792
rect 7748 6740 7800 6792
rect 8208 6808 8260 6860
rect 8392 6808 8444 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9128 6808 9180 6860
rect 9680 6808 9732 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 15016 6851 15068 6860
rect 14280 6808 14332 6817
rect 9404 6740 9456 6792
rect 5816 6672 5868 6724
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 6276 6647 6328 6656
rect 5264 6604 5316 6613
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 6644 6672 6696 6724
rect 7196 6672 7248 6724
rect 12164 6740 12216 6792
rect 14372 6740 14424 6792
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15108 6808 15160 6860
rect 15476 6740 15528 6792
rect 10416 6672 10468 6724
rect 6460 6604 6512 6656
rect 7564 6604 7616 6656
rect 8300 6604 8352 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 8852 6604 8904 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9404 6604 9456 6656
rect 18604 6808 18656 6860
rect 20076 6876 20128 6928
rect 20352 6808 20404 6860
rect 17132 6783 17184 6792
rect 17132 6749 17150 6783
rect 17150 6749 17184 6783
rect 17132 6740 17184 6749
rect 17316 6740 17368 6792
rect 17776 6783 17828 6792
rect 17776 6749 17810 6783
rect 17810 6749 17828 6783
rect 17776 6740 17828 6749
rect 19432 6740 19484 6792
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 17960 6672 18012 6724
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11244 6604 11296 6656
rect 11796 6604 11848 6656
rect 12716 6604 12768 6656
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 15660 6604 15712 6656
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 16212 6604 16264 6656
rect 17040 6604 17092 6656
rect 18880 6604 18932 6656
rect 19524 6604 19576 6656
rect 19708 6604 19760 6656
rect 21548 6604 21600 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 2964 6400 3016 6452
rect 3240 6400 3292 6452
rect 3792 6400 3844 6452
rect 8116 6400 8168 6452
rect 8760 6400 8812 6452
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 11980 6443 12032 6452
rect 3608 6332 3660 6384
rect 4436 6332 4488 6384
rect 4528 6332 4580 6384
rect 6644 6332 6696 6384
rect 7748 6332 7800 6384
rect 9496 6332 9548 6384
rect 10048 6332 10100 6384
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 14372 6400 14424 6452
rect 15936 6400 15988 6452
rect 16948 6400 17000 6452
rect 17500 6443 17552 6452
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 17776 6400 17828 6452
rect 2412 6196 2464 6248
rect 2872 6264 2924 6316
rect 2780 6196 2832 6248
rect 3516 6196 3568 6248
rect 3700 6196 3752 6248
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 4252 6128 4304 6180
rect 6552 6264 6604 6316
rect 7656 6264 7708 6316
rect 1492 6060 1544 6069
rect 3332 6060 3384 6112
rect 4068 6060 4120 6112
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 7380 6239 7432 6248
rect 6920 6196 6972 6205
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 6184 6171 6236 6180
rect 6184 6137 6193 6171
rect 6193 6137 6227 6171
rect 6227 6137 6236 6171
rect 8116 6239 8168 6248
rect 8116 6205 8125 6239
rect 8125 6205 8159 6239
rect 8159 6205 8168 6239
rect 8116 6196 8168 6205
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 12164 6332 12216 6384
rect 13084 6375 13136 6384
rect 13084 6341 13093 6375
rect 13093 6341 13127 6375
rect 13127 6341 13136 6375
rect 13084 6332 13136 6341
rect 14280 6332 14332 6384
rect 14832 6332 14884 6384
rect 19892 6400 19944 6452
rect 20352 6332 20404 6384
rect 20536 6332 20588 6384
rect 22468 6332 22520 6384
rect 6184 6128 6236 6137
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 7656 6060 7708 6112
rect 8576 6060 8628 6112
rect 9588 6060 9640 6112
rect 10048 6060 10100 6112
rect 10416 6128 10468 6180
rect 11152 6128 11204 6180
rect 11612 6128 11664 6180
rect 11704 6060 11756 6112
rect 12900 6196 12952 6248
rect 15016 6264 15068 6316
rect 15108 6264 15160 6316
rect 17500 6264 17552 6316
rect 12164 6128 12216 6180
rect 13084 6128 13136 6180
rect 13820 6128 13872 6180
rect 15384 6128 15436 6180
rect 15936 6196 15988 6248
rect 15752 6128 15804 6180
rect 17408 6196 17460 6248
rect 17776 6196 17828 6248
rect 19892 6264 19944 6316
rect 19708 6239 19760 6248
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 20260 6239 20312 6248
rect 20260 6205 20269 6239
rect 20269 6205 20303 6239
rect 20303 6205 20312 6239
rect 20260 6196 20312 6205
rect 20812 6264 20864 6316
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21548 6264 21600 6316
rect 15844 6060 15896 6112
rect 19892 6128 19944 6180
rect 17316 6060 17368 6112
rect 17500 6060 17552 6112
rect 21364 6060 21416 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1400 5856 1452 5908
rect 3148 5856 3200 5908
rect 4436 5856 4488 5908
rect 5540 5831 5592 5840
rect 5540 5797 5549 5831
rect 5549 5797 5583 5831
rect 5583 5797 5592 5831
rect 5540 5788 5592 5797
rect 2136 5720 2188 5772
rect 3332 5763 3384 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 4068 5720 4120 5772
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 5724 5720 5776 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 6736 5856 6788 5908
rect 9128 5856 9180 5908
rect 10324 5856 10376 5908
rect 11428 5856 11480 5908
rect 11704 5856 11756 5908
rect 11980 5856 12032 5908
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 8668 5788 8720 5840
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 8116 5720 8168 5772
rect 8852 5720 8904 5772
rect 6368 5652 6420 5704
rect 7288 5652 7340 5704
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 8300 5652 8352 5704
rect 8484 5652 8536 5704
rect 8760 5652 8812 5704
rect 1584 5584 1636 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 4068 5584 4120 5636
rect 4712 5584 4764 5636
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 4344 5516 4396 5568
rect 4988 5516 5040 5568
rect 6552 5584 6604 5636
rect 9496 5652 9548 5704
rect 13636 5720 13688 5772
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11612 5652 11664 5704
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 6828 5516 6880 5525
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 8392 5516 8444 5568
rect 8484 5516 8536 5568
rect 9588 5584 9640 5636
rect 10140 5584 10192 5636
rect 10416 5516 10468 5568
rect 11152 5584 11204 5636
rect 12164 5652 12216 5704
rect 12256 5652 12308 5704
rect 17040 5856 17092 5908
rect 19892 5856 19944 5908
rect 18144 5788 18196 5840
rect 20260 5856 20312 5908
rect 21088 5856 21140 5908
rect 22100 5856 22152 5908
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16764 5763 16816 5772
rect 16764 5729 16773 5763
rect 16773 5729 16807 5763
rect 16807 5729 16816 5763
rect 16764 5720 16816 5729
rect 15384 5695 15436 5704
rect 15384 5661 15402 5695
rect 15402 5661 15436 5695
rect 15384 5652 15436 5661
rect 12808 5584 12860 5636
rect 15752 5652 15804 5704
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 18052 5720 18104 5772
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17776 5652 17828 5704
rect 16580 5584 16632 5636
rect 17500 5584 17552 5636
rect 11244 5559 11296 5568
rect 11244 5525 11253 5559
rect 11253 5525 11287 5559
rect 11287 5525 11296 5559
rect 11244 5516 11296 5525
rect 11428 5516 11480 5568
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 14280 5559 14332 5568
rect 12716 5516 12768 5525
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 15384 5516 15436 5568
rect 15568 5516 15620 5568
rect 17316 5559 17368 5568
rect 17316 5525 17325 5559
rect 17325 5525 17359 5559
rect 17359 5525 17368 5559
rect 17316 5516 17368 5525
rect 18880 5516 18932 5568
rect 22284 5652 22336 5704
rect 19524 5627 19576 5636
rect 19524 5593 19558 5627
rect 19558 5593 19576 5627
rect 19524 5584 19576 5593
rect 21364 5584 21416 5636
rect 22192 5584 22244 5636
rect 20076 5516 20128 5568
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 21272 5516 21324 5568
rect 21640 5516 21692 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2044 5312 2096 5364
rect 3240 5312 3292 5364
rect 4252 5312 4304 5364
rect 5356 5312 5408 5364
rect 5540 5312 5592 5364
rect 6552 5312 6604 5364
rect 7288 5312 7340 5364
rect 7840 5312 7892 5364
rect 8484 5312 8536 5364
rect 1676 5287 1728 5296
rect 1676 5253 1685 5287
rect 1685 5253 1719 5287
rect 1719 5253 1728 5287
rect 1676 5244 1728 5253
rect 1768 5244 1820 5296
rect 2596 5244 2648 5296
rect 5080 5287 5132 5296
rect 5080 5253 5089 5287
rect 5089 5253 5123 5287
rect 5123 5253 5132 5287
rect 5080 5244 5132 5253
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 7564 5244 7616 5296
rect 8852 5244 8904 5296
rect 9588 5312 9640 5364
rect 10324 5312 10376 5364
rect 10784 5312 10836 5364
rect 10876 5312 10928 5364
rect 12716 5312 12768 5364
rect 15568 5355 15620 5364
rect 15568 5321 15577 5355
rect 15577 5321 15611 5355
rect 15611 5321 15620 5355
rect 15568 5312 15620 5321
rect 16396 5355 16448 5364
rect 16396 5321 16405 5355
rect 16405 5321 16439 5355
rect 16439 5321 16448 5355
rect 16396 5312 16448 5321
rect 17316 5312 17368 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 20812 5312 20864 5364
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 4252 5176 4304 5228
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5172 5176 5224 5228
rect 5540 5176 5592 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8668 5176 8720 5228
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 4068 5108 4120 5160
rect 4436 5040 4488 5092
rect 4896 5108 4948 5160
rect 5724 5108 5776 5160
rect 6552 5108 6604 5160
rect 6920 5108 6972 5160
rect 7288 5108 7340 5160
rect 8760 5108 8812 5160
rect 8944 5176 8996 5228
rect 9496 5176 9548 5228
rect 9864 5244 9916 5296
rect 10692 5244 10744 5296
rect 13636 5244 13688 5296
rect 16028 5244 16080 5296
rect 16120 5244 16172 5296
rect 8668 5040 8720 5092
rect 4344 4972 4396 5024
rect 6000 4972 6052 5024
rect 7656 4972 7708 5024
rect 8300 4972 8352 5024
rect 10140 4972 10192 5024
rect 11704 5176 11756 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 17040 5176 17092 5228
rect 18880 5244 18932 5296
rect 18972 5244 19024 5296
rect 18236 5176 18288 5228
rect 19616 5176 19668 5228
rect 10324 5108 10376 5160
rect 11336 5108 11388 5160
rect 10692 4972 10744 5024
rect 11152 4972 11204 5024
rect 12164 5040 12216 5092
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 15384 5108 15436 5160
rect 15936 5108 15988 5160
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 16396 5108 16448 5160
rect 16764 5151 16816 5160
rect 16764 5117 16773 5151
rect 16773 5117 16807 5151
rect 16807 5117 16816 5151
rect 16764 5108 16816 5117
rect 16856 5108 16908 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 19524 5108 19576 5160
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 16212 5040 16264 5092
rect 20904 5244 20956 5296
rect 14372 4972 14424 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14648 5015 14700 5024
rect 14464 4972 14516 4981
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 14924 4972 14976 5024
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 18880 4972 18932 5024
rect 21548 5015 21600 5024
rect 21548 4981 21557 5015
rect 21557 4981 21591 5015
rect 21591 4981 21600 5015
rect 21548 4972 21600 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 2504 4768 2556 4820
rect 4436 4768 4488 4820
rect 4620 4768 4672 4820
rect 4252 4700 4304 4752
rect 5632 4700 5684 4752
rect 6092 4768 6144 4820
rect 7104 4768 7156 4820
rect 8208 4811 8260 4820
rect 8208 4777 8217 4811
rect 8217 4777 8251 4811
rect 8251 4777 8260 4811
rect 8208 4768 8260 4777
rect 8392 4768 8444 4820
rect 9772 4768 9824 4820
rect 10968 4768 11020 4820
rect 11244 4768 11296 4820
rect 11612 4768 11664 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 12532 4768 12584 4820
rect 13728 4768 13780 4820
rect 15660 4768 15712 4820
rect 15936 4768 15988 4820
rect 2964 4496 3016 4548
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 6000 4675 6052 4684
rect 4988 4632 5040 4641
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 7104 4632 7156 4684
rect 7288 4632 7340 4684
rect 7472 4700 7524 4752
rect 8760 4743 8812 4752
rect 8760 4709 8769 4743
rect 8769 4709 8803 4743
rect 8803 4709 8812 4743
rect 8760 4700 8812 4709
rect 9404 4700 9456 4752
rect 10692 4700 10744 4752
rect 7564 4632 7616 4684
rect 7932 4632 7984 4684
rect 8116 4632 8168 4684
rect 8392 4632 8444 4684
rect 9496 4675 9548 4684
rect 7840 4564 7892 4616
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 10600 4632 10652 4684
rect 12164 4700 12216 4752
rect 14280 4700 14332 4752
rect 16856 4768 16908 4820
rect 17132 4768 17184 4820
rect 17868 4768 17920 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 19708 4768 19760 4820
rect 22560 4768 22612 4820
rect 20076 4743 20128 4752
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 10140 4564 10192 4616
rect 11060 4564 11112 4616
rect 11612 4632 11664 4684
rect 11888 4632 11940 4684
rect 11704 4564 11756 4616
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 20076 4709 20085 4743
rect 20085 4709 20119 4743
rect 20119 4709 20128 4743
rect 20076 4700 20128 4709
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 16028 4632 16080 4684
rect 16120 4632 16172 4684
rect 16672 4632 16724 4684
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 17868 4632 17920 4684
rect 13268 4564 13320 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2688 4428 2740 4480
rect 4068 4428 4120 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 7380 4471 7432 4480
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 7564 4428 7616 4480
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 8484 4496 8536 4548
rect 8760 4496 8812 4548
rect 8852 4496 8904 4548
rect 12440 4496 12492 4548
rect 13728 4564 13780 4616
rect 14648 4564 14700 4616
rect 15752 4564 15804 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 7840 4428 7892 4437
rect 10416 4428 10468 4480
rect 10600 4428 10652 4480
rect 10876 4471 10928 4480
rect 10876 4437 10885 4471
rect 10885 4437 10919 4471
rect 10919 4437 10928 4471
rect 10876 4428 10928 4437
rect 11060 4428 11112 4480
rect 11980 4471 12032 4480
rect 11980 4437 11989 4471
rect 11989 4437 12023 4471
rect 12023 4437 12032 4471
rect 11980 4428 12032 4437
rect 12532 4428 12584 4480
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 14648 4471 14700 4480
rect 14648 4437 14657 4471
rect 14657 4437 14691 4471
rect 14691 4437 14700 4471
rect 14648 4428 14700 4437
rect 14832 4428 14884 4480
rect 18052 4564 18104 4616
rect 22376 4564 22428 4616
rect 15200 4471 15252 4480
rect 15200 4437 15209 4471
rect 15209 4437 15243 4471
rect 15243 4437 15252 4471
rect 15200 4428 15252 4437
rect 16212 4428 16264 4480
rect 16764 4428 16816 4480
rect 16948 4428 17000 4480
rect 21640 4496 21692 4548
rect 17868 4428 17920 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 18880 4428 18932 4480
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 19708 4471 19760 4480
rect 19708 4437 19717 4471
rect 19717 4437 19751 4471
rect 19751 4437 19760 4471
rect 19708 4428 19760 4437
rect 21180 4471 21232 4480
rect 21180 4437 21189 4471
rect 21189 4437 21223 4471
rect 21223 4437 21232 4471
rect 21180 4428 21232 4437
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 2412 4224 2464 4276
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 5540 4224 5592 4276
rect 6552 4224 6604 4276
rect 6920 4224 6972 4276
rect 7288 4224 7340 4276
rect 8576 4267 8628 4276
rect 2780 4156 2832 4208
rect 4896 4156 4948 4208
rect 7932 4156 7984 4208
rect 8576 4233 8585 4267
rect 8585 4233 8619 4267
rect 8619 4233 8628 4267
rect 8576 4224 8628 4233
rect 8668 4224 8720 4276
rect 9128 4267 9180 4276
rect 9128 4233 9137 4267
rect 9137 4233 9171 4267
rect 9171 4233 9180 4267
rect 9128 4224 9180 4233
rect 11612 4224 11664 4276
rect 11980 4224 12032 4276
rect 12256 4224 12308 4276
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 3332 4088 3384 4140
rect 2136 4063 2188 4072
rect 2136 4029 2145 4063
rect 2145 4029 2179 4063
rect 2179 4029 2188 4063
rect 2136 4020 2188 4029
rect 1492 3884 1544 3936
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 4436 4020 4488 4072
rect 5080 4088 5132 4140
rect 6184 4088 6236 4140
rect 6920 4088 6972 4140
rect 8668 4131 8720 4140
rect 6092 4020 6144 4072
rect 6644 3952 6696 4004
rect 4528 3927 4580 3936
rect 1768 3884 1820 3893
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 4528 3884 4580 3893
rect 6000 3884 6052 3936
rect 7104 3884 7156 3936
rect 8300 3884 8352 3936
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 9680 4156 9732 4208
rect 9036 4088 9088 4140
rect 9588 4088 9640 4140
rect 10048 4131 10100 4140
rect 10048 4097 10057 4131
rect 10057 4097 10091 4131
rect 10091 4097 10100 4131
rect 10048 4088 10100 4097
rect 10876 4088 10928 4140
rect 9220 3952 9272 4004
rect 11336 4088 11388 4140
rect 12164 4088 12216 4140
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 12440 4088 12492 4140
rect 14464 4156 14516 4208
rect 15200 4224 15252 4276
rect 15752 4224 15804 4276
rect 17132 4224 17184 4276
rect 17408 4224 17460 4276
rect 18328 4224 18380 4276
rect 19248 4224 19300 4276
rect 20076 4224 20128 4276
rect 22100 4224 22152 4276
rect 14924 4156 14976 4208
rect 15660 4156 15712 4208
rect 17224 4156 17276 4208
rect 13820 4088 13872 4140
rect 16120 4088 16172 4140
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17684 4131 17736 4140
rect 17040 4088 17092 4097
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 11612 4063 11664 4072
rect 10324 3884 10376 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 10968 3952 11020 4004
rect 11612 4029 11621 4063
rect 11621 4029 11655 4063
rect 11655 4029 11664 4063
rect 11612 4020 11664 4029
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 12256 4063 12308 4072
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 12256 4020 12308 4029
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13728 4020 13780 4072
rect 14464 4020 14516 4072
rect 14556 4020 14608 4072
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 14740 4020 14792 4029
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 17132 4020 17184 4072
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 19892 4156 19944 4208
rect 19800 4088 19852 4140
rect 19524 4063 19576 4072
rect 11428 3952 11480 4004
rect 12164 3952 12216 4004
rect 16856 3952 16908 4004
rect 11520 3884 11572 3936
rect 12440 3884 12492 3936
rect 12900 3884 12952 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 14556 3884 14608 3936
rect 15016 3884 15068 3936
rect 17960 3952 18012 4004
rect 19524 4029 19533 4063
rect 19533 4029 19567 4063
rect 19567 4029 19576 4063
rect 19524 4020 19576 4029
rect 19616 3952 19668 4004
rect 20352 3952 20404 4004
rect 18972 3927 19024 3936
rect 18972 3893 18981 3927
rect 18981 3893 19015 3927
rect 19015 3893 19024 3927
rect 20076 3927 20128 3936
rect 18972 3884 19024 3893
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1952 3680 2004 3732
rect 4252 3680 4304 3732
rect 8668 3723 8720 3732
rect 2504 3587 2556 3596
rect 2504 3553 2513 3587
rect 2513 3553 2547 3587
rect 2547 3553 2556 3587
rect 2504 3544 2556 3553
rect 2596 3587 2648 3596
rect 2596 3553 2605 3587
rect 2605 3553 2639 3587
rect 2639 3553 2648 3587
rect 2596 3544 2648 3553
rect 2780 3476 2832 3528
rect 3332 3544 3384 3596
rect 4160 3612 4212 3664
rect 4436 3612 4488 3664
rect 5908 3612 5960 3664
rect 4528 3544 4580 3596
rect 4896 3544 4948 3596
rect 5632 3587 5684 3596
rect 5632 3553 5641 3587
rect 5641 3553 5675 3587
rect 5675 3553 5684 3587
rect 5632 3544 5684 3553
rect 6000 3544 6052 3596
rect 4160 3476 4212 3528
rect 8668 3689 8677 3723
rect 8677 3689 8711 3723
rect 8711 3689 8720 3723
rect 8668 3680 8720 3689
rect 10600 3680 10652 3732
rect 11612 3680 11664 3732
rect 10416 3655 10468 3664
rect 10416 3621 10425 3655
rect 10425 3621 10459 3655
rect 10459 3621 10468 3655
rect 10416 3612 10468 3621
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 3884 3408 3936 3460
rect 5908 3408 5960 3460
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 3148 3340 3200 3392
rect 3240 3340 3292 3392
rect 7472 3340 7524 3392
rect 8208 3544 8260 3596
rect 12256 3680 12308 3732
rect 14740 3680 14792 3732
rect 16120 3680 16172 3732
rect 8300 3476 8352 3528
rect 8576 3408 8628 3460
rect 9036 3476 9088 3528
rect 9496 3476 9548 3528
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 12348 3476 12400 3528
rect 12808 3476 12860 3528
rect 13820 3476 13872 3528
rect 13912 3519 13964 3528
rect 13912 3485 13921 3519
rect 13921 3485 13955 3519
rect 13955 3485 13964 3519
rect 13912 3476 13964 3485
rect 9772 3408 9824 3460
rect 9036 3340 9088 3392
rect 10324 3383 10376 3392
rect 10324 3349 10333 3383
rect 10333 3349 10367 3383
rect 10367 3349 10376 3383
rect 10324 3340 10376 3349
rect 10692 3340 10744 3392
rect 12072 3408 12124 3460
rect 13452 3408 13504 3460
rect 13728 3408 13780 3460
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 14924 3544 14976 3596
rect 14464 3476 14516 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 16488 3612 16540 3664
rect 16028 3544 16080 3596
rect 17684 3680 17736 3732
rect 17960 3680 18012 3732
rect 19064 3680 19116 3732
rect 17592 3612 17644 3664
rect 18972 3612 19024 3664
rect 15384 3476 15436 3485
rect 16396 3476 16448 3528
rect 17408 3476 17460 3528
rect 17868 3587 17920 3596
rect 17868 3553 17877 3587
rect 17877 3553 17911 3587
rect 17911 3553 17920 3587
rect 17868 3544 17920 3553
rect 19524 3544 19576 3596
rect 19064 3476 19116 3528
rect 17960 3408 18012 3460
rect 18420 3408 18472 3460
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 14372 3340 14424 3392
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 16212 3383 16264 3392
rect 16212 3349 16221 3383
rect 16221 3349 16255 3383
rect 16255 3349 16264 3383
rect 16212 3340 16264 3349
rect 16488 3340 16540 3392
rect 19708 3340 19760 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 2412 3136 2464 3188
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 3240 3136 3292 3188
rect 3516 3136 3568 3188
rect 7380 3136 7432 3188
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 9220 3136 9272 3188
rect 12624 3136 12676 3188
rect 12808 3136 12860 3188
rect 14924 3136 14976 3188
rect 15108 3136 15160 3188
rect 2964 3068 3016 3120
rect 6644 3068 6696 3120
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 1860 2932 1912 2984
rect 4436 3000 4488 3052
rect 7656 3068 7708 3120
rect 7196 3000 7248 3052
rect 6920 2975 6972 2984
rect 2872 2864 2924 2916
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 7288 2932 7340 2984
rect 7472 2932 7524 2984
rect 8024 2932 8076 2984
rect 10324 3068 10376 3120
rect 10508 3068 10560 3120
rect 6552 2864 6604 2916
rect 9496 3000 9548 3052
rect 10784 3000 10836 3052
rect 12164 3068 12216 3120
rect 12532 3068 12584 3120
rect 13544 3068 13596 3120
rect 13544 2975 13596 2984
rect 13544 2941 13553 2975
rect 13553 2941 13587 2975
rect 13587 2941 13596 2975
rect 13544 2932 13596 2941
rect 13912 2932 13964 2984
rect 14648 3000 14700 3052
rect 16212 3068 16264 3120
rect 15108 3043 15160 3052
rect 14280 2932 14332 2984
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15292 3043 15344 3052
rect 15292 3009 15301 3043
rect 15301 3009 15335 3043
rect 15335 3009 15344 3043
rect 15292 3000 15344 3009
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 16304 3000 16356 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17592 3068 17644 3120
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17776 3043 17828 3052
rect 17408 3000 17460 3009
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 18788 3000 18840 3052
rect 15568 2975 15620 2984
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 16120 2975 16172 2984
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 5080 2796 5132 2848
rect 9772 2864 9824 2916
rect 9588 2796 9640 2848
rect 12072 2796 12124 2848
rect 14372 2864 14424 2916
rect 16212 2864 16264 2916
rect 18788 2864 18840 2916
rect 19524 2864 19576 2916
rect 13268 2796 13320 2848
rect 13728 2796 13780 2848
rect 16948 2796 17000 2848
rect 17316 2796 17368 2848
rect 17684 2796 17736 2848
rect 18972 2796 19024 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3056 2592 3108 2644
rect 5908 2592 5960 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 7840 2592 7892 2644
rect 9128 2592 9180 2644
rect 1952 2524 2004 2576
rect 4068 2456 4120 2508
rect 7196 2524 7248 2576
rect 11152 2524 11204 2576
rect 12808 2524 12860 2576
rect 13360 2592 13412 2644
rect 16672 2635 16724 2644
rect 13544 2524 13596 2576
rect 4528 2456 4580 2508
rect 7288 2456 7340 2508
rect 9588 2456 9640 2508
rect 10784 2499 10836 2508
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5080 2431 5132 2440
rect 5080 2397 5114 2431
rect 5114 2397 5132 2431
rect 5080 2388 5132 2397
rect 5908 2320 5960 2372
rect 8392 2388 8444 2440
rect 8484 2388 8536 2440
rect 9956 2388 10008 2440
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 10968 2388 11020 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13452 2456 13504 2508
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 17408 2592 17460 2644
rect 17776 2592 17828 2644
rect 18144 2592 18196 2644
rect 18512 2592 18564 2644
rect 15476 2524 15528 2576
rect 17040 2524 17092 2576
rect 15200 2456 15252 2508
rect 6644 2320 6696 2372
rect 3700 2252 3752 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 8484 2295 8536 2304
rect 7196 2252 7248 2261
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 8576 2252 8628 2304
rect 15568 2388 15620 2440
rect 16120 2388 16172 2440
rect 11244 2252 11296 2304
rect 12532 2252 12584 2304
rect 15108 2252 15160 2304
rect 15752 2252 15804 2304
rect 18420 2320 18472 2372
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 2228 2048 2280 2100
rect 3792 2048 3844 2100
rect 3976 2048 4028 2100
rect 7196 2048 7248 2100
rect 3332 1980 3384 2032
rect 5908 1980 5960 2032
rect 7104 1980 7156 2032
rect 13176 1980 13228 2032
rect 2596 1912 2648 1964
rect 8484 1912 8536 1964
rect 3792 1844 3844 1896
rect 8576 1844 8628 1896
rect 12348 1844 12400 1896
rect 8484 1504 8536 1556
rect 9220 1504 9272 1556
rect 5724 1368 5776 1420
rect 6276 1368 6328 1420
<< metal2 >>
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 6932 22222 7144 22250
rect 584 18426 612 22200
rect 952 20602 980 22200
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1320 20330 1348 22200
rect 1308 20324 1360 20330
rect 1308 20266 1360 20272
rect 572 18420 624 18426
rect 572 18362 624 18368
rect 1320 18358 1348 20266
rect 1688 20058 1716 22200
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1964 19417 1992 19450
rect 2056 19446 2084 22200
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2044 19440 2096 19446
rect 1950 19408 2006 19417
rect 2044 19382 2096 19388
rect 2240 19378 2268 19654
rect 2332 19514 2360 19751
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 1950 19343 2006 19352
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 1582 19000 1638 19009
rect 1582 18935 1584 18944
rect 1636 18935 1638 18944
rect 1584 18906 1636 18912
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1950 18592 2006 18601
rect 1950 18527 2006 18536
rect 1964 18426 1992 18527
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1308 18352 1360 18358
rect 1308 18294 1360 18300
rect 1766 18184 1822 18193
rect 1766 18119 1822 18128
rect 1780 17882 1808 18119
rect 2148 18086 2176 18702
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1780 17338 1808 17711
rect 1952 17672 2004 17678
rect 1950 17640 1952 17649
rect 2004 17640 2006 17649
rect 1950 17575 2006 17584
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1858 17368 1914 17377
rect 1768 17332 1820 17338
rect 1858 17303 1914 17312
rect 1768 17274 1820 17280
rect 1872 16794 1900 17303
rect 2056 17270 2084 17478
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2056 16726 2084 17206
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 1858 16552 1914 16561
rect 1858 16487 1914 16496
rect 1872 15706 1900 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1964 16153 1992 16186
rect 1950 16144 2006 16153
rect 1950 16079 2006 16088
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1766 15328 1822 15337
rect 1766 15263 1822 15272
rect 1780 15162 1808 15263
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 2148 15065 2176 18022
rect 2240 17241 2268 19314
rect 2424 19242 2452 22200
rect 2792 19718 2820 22200
rect 3160 19802 3188 22200
rect 3528 20346 3556 22200
rect 3698 22128 3754 22137
rect 3698 22063 3754 22072
rect 2976 19774 3188 19802
rect 3436 20318 3556 20346
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 2608 19378 2636 19654
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2884 19258 2912 19314
rect 2412 19236 2464 19242
rect 2412 19178 2464 19184
rect 2792 19230 2912 19258
rect 2792 19009 2820 19230
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2778 19000 2834 19009
rect 2778 18935 2834 18944
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18426 2360 18566
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2226 17232 2282 17241
rect 2226 17167 2282 17176
rect 2332 16590 2360 18226
rect 2792 17678 2820 18770
rect 2884 18766 2912 19110
rect 2976 18834 3004 19774
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3068 19378 3096 19654
rect 3160 19446 3188 19654
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 3068 18358 3096 19314
rect 3160 18902 3188 19382
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3148 18896 3200 18902
rect 3148 18838 3200 18844
rect 3146 18728 3202 18737
rect 3252 18698 3280 19178
rect 3344 18970 3372 19450
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3146 18663 3202 18672
rect 3240 18692 3292 18698
rect 3160 18408 3188 18663
rect 3240 18634 3292 18640
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3160 18380 3280 18408
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 17048 2820 17614
rect 2884 17338 2912 18158
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2792 17020 2912 17048
rect 2778 16960 2834 16969
rect 2778 16895 2834 16904
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2240 15502 2268 15846
rect 2318 15736 2374 15745
rect 2318 15671 2320 15680
rect 2372 15671 2374 15680
rect 2320 15642 2372 15648
rect 2608 15609 2636 16526
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2594 15600 2650 15609
rect 2594 15535 2650 15544
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2134 15056 2190 15065
rect 2134 14991 2190 15000
rect 1584 14544 1636 14550
rect 1582 14512 1584 14521
rect 1636 14512 1638 14521
rect 1582 14447 1638 14456
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 12986 1624 13631
rect 1688 13326 1716 14010
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13394 1992 13670
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1858 13288 1914 13297
rect 1858 13223 1914 13232
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1582 12472 1638 12481
rect 1872 12442 1900 13223
rect 1964 12918 1992 13330
rect 1952 12912 2004 12918
rect 1952 12854 2004 12860
rect 1582 12407 1584 12416
rect 1636 12407 1638 12416
rect 1860 12436 1912 12442
rect 1584 12378 1636 12384
rect 1860 12378 1912 12384
rect 2240 12322 2268 15438
rect 2608 14482 2636 15438
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 13530 2360 14350
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 14113 2544 14214
rect 2502 14104 2558 14113
rect 2502 14039 2558 14048
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2410 12880 2466 12889
rect 2410 12815 2466 12824
rect 2424 12442 2452 12815
rect 2608 12782 2636 13262
rect 2596 12776 2648 12782
rect 2700 12753 2728 15846
rect 2792 15706 2820 16895
rect 2884 16046 2912 17020
rect 3068 16454 3096 18158
rect 3160 16522 3188 18226
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2870 14920 2926 14929
rect 2870 14855 2926 14864
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14550 2820 14758
rect 2884 14618 2912 14855
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2596 12718 2648 12724
rect 2686 12744 2742 12753
rect 2686 12679 2742 12688
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2516 12374 2544 12582
rect 2976 12434 3004 15846
rect 3056 15088 3108 15094
rect 3056 15030 3108 15036
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3068 14226 3096 15030
rect 3160 14414 3188 15030
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3068 14198 3188 14226
rect 3160 14006 3188 14198
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3148 14000 3200 14006
rect 3252 13977 3280 18380
rect 3344 16590 3372 18566
rect 3436 18057 3464 20318
rect 3712 20262 3740 22063
rect 3896 21162 3924 22200
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 3974 21448 4030 21457
rect 3974 21383 4030 21392
rect 3804 21134 3924 21162
rect 3804 20346 3832 21134
rect 3882 21040 3938 21049
rect 3882 20975 3884 20984
rect 3936 20975 3938 20984
rect 3884 20946 3936 20952
rect 3988 20505 4016 21383
rect 4080 20806 4108 21791
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3974 20496 4030 20505
rect 3974 20431 4030 20440
rect 3804 20318 4108 20346
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3896 19514 3924 19722
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 3620 18630 3648 18838
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3620 18086 3648 18566
rect 3792 18216 3844 18222
rect 3896 18204 3924 19450
rect 3974 19408 4030 19417
rect 3974 19343 4030 19352
rect 3844 18176 3924 18204
rect 3792 18158 3844 18164
rect 3988 18154 4016 19343
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3608 18080 3660 18086
rect 3422 18048 3478 18057
rect 3608 18022 3660 18028
rect 4080 18034 4108 20318
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4172 19378 4200 19790
rect 4160 19372 4212 19378
rect 4160 19314 4212 19320
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4172 18902 4200 19110
rect 4160 18896 4212 18902
rect 4158 18864 4160 18873
rect 4212 18864 4214 18873
rect 4158 18799 4214 18808
rect 4080 18006 4200 18034
rect 3422 17983 3478 17992
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3528 17134 3556 17614
rect 4172 17354 4200 18006
rect 4264 17542 4292 22200
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4540 18737 4568 18770
rect 4526 18728 4582 18737
rect 4526 18663 4582 18672
rect 4528 18216 4580 18222
rect 4528 18158 4580 18164
rect 4540 17882 4568 18158
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4632 17678 4660 22200
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4724 19786 4752 20198
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4724 18834 4752 19450
rect 4802 19000 4858 19009
rect 4802 18935 4804 18944
rect 4856 18935 4858 18944
rect 4804 18906 4856 18912
rect 4896 18896 4948 18902
rect 4896 18838 4948 18844
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4252 17536 4304 17542
rect 4540 17524 4568 17614
rect 4540 17496 4660 17524
rect 4252 17478 4304 17484
rect 4172 17326 4476 17354
rect 3608 17264 3660 17270
rect 3884 17264 3936 17270
rect 3660 17224 3884 17252
rect 3608 17206 3660 17212
rect 3884 17206 3936 17212
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15570 3464 16050
rect 3712 15978 3740 16390
rect 3896 16250 3924 16390
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3896 14958 3924 16050
rect 4080 15162 4108 16458
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3344 14346 3372 14486
rect 3422 14376 3478 14385
rect 3332 14340 3384 14346
rect 3422 14311 3424 14320
rect 3332 14282 3384 14288
rect 3476 14311 3478 14320
rect 3424 14282 3476 14288
rect 3988 14278 4016 14962
rect 4066 14920 4122 14929
rect 4066 14855 4122 14864
rect 4080 14550 4108 14855
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3976 14272 4028 14278
rect 3974 14240 3976 14249
rect 4028 14240 4030 14249
rect 3974 14175 4030 14184
rect 4172 14006 4200 15642
rect 4160 14000 4212 14006
rect 3148 13942 3200 13948
rect 3238 13968 3294 13977
rect 3068 13190 3096 13942
rect 4160 13942 4212 13948
rect 3238 13903 3294 13912
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3148 13252 3200 13258
rect 3148 13194 3200 13200
rect 3332 13252 3384 13258
rect 3332 13194 3384 13200
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 3068 12986 3096 13126
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3160 12442 3188 13194
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3148 12436 3200 12442
rect 2976 12406 3096 12434
rect 2504 12368 2556 12374
rect 2240 12294 2360 12322
rect 2504 12310 2556 12316
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1216 8356 1268 8362
rect 1216 8298 1268 8304
rect 1228 7177 1256 8298
rect 1214 7168 1270 7177
rect 1214 7103 1270 7112
rect 1412 5914 1440 11999
rect 2240 11898 2268 12174
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10674 1532 11086
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 9450 1716 10610
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2056 9722 2084 9862
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1688 9042 1716 9386
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1504 6866 1532 7414
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1596 6458 1624 8842
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8634 1808 8774
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1504 5574 1532 6054
rect 1688 5794 1716 8366
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7206 1808 7686
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1596 5766 1716 5794
rect 1596 5642 1624 5766
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1504 3942 1532 5510
rect 1596 4486 1624 5578
rect 1688 5302 1716 5646
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1768 5296 1820 5302
rect 1768 5238 1820 5244
rect 1780 4826 1808 5238
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1490 2952 1546 2961
rect 1490 2887 1546 2896
rect 1504 800 1532 2887
rect 1596 2689 1624 4422
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3505 1808 3878
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1872 3097 1900 8502
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 6458 1992 7686
rect 2056 7546 2084 9522
rect 2148 8838 2176 9862
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 9178 2268 9454
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2136 8288 2188 8294
rect 2136 8230 2188 8236
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2148 7478 2176 8230
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2240 7002 2268 7890
rect 2332 7449 2360 12294
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 8634 2452 12038
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2516 8634 2544 11766
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2608 10470 2636 11018
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10130 2636 10406
rect 2700 10266 2728 11698
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2792 10266 2820 11630
rect 2976 11354 3004 11630
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2884 10146 2912 11222
rect 2976 10742 3004 11290
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 3068 10554 3096 12406
rect 3148 12378 3200 12384
rect 3252 12238 3280 13126
rect 3344 12306 3372 13194
rect 3988 12986 4016 13738
rect 4080 13462 4108 13806
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4172 13394 4200 13942
rect 4264 13530 4292 15982
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 14822 4384 15302
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4250 13424 4306 13433
rect 4160 13388 4212 13394
rect 4356 13394 4384 14758
rect 4250 13359 4306 13368
rect 4344 13388 4396 13394
rect 4160 13330 4212 13336
rect 4160 13252 4212 13258
rect 4264 13240 4292 13359
rect 4344 13330 4396 13336
rect 4212 13212 4292 13240
rect 4160 13194 4212 13200
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3896 12434 3924 12582
rect 3528 12406 3924 12434
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2792 10118 2912 10146
rect 2976 10526 3096 10554
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2608 8974 2636 9590
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2516 8430 2544 8570
rect 2608 8566 2636 8910
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2608 8430 2636 8502
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7478 2544 7686
rect 2504 7472 2556 7478
rect 2318 7440 2374 7449
rect 2504 7414 2556 7420
rect 2318 7375 2374 7384
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2148 5778 2176 6666
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5370 2084 5510
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 3738 1992 5170
rect 2148 4078 2176 5714
rect 2240 5166 2268 6598
rect 2424 6254 2452 7210
rect 2516 7188 2544 7414
rect 2608 7342 2636 8366
rect 2792 8362 2820 10118
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2884 8498 2912 8842
rect 2976 8809 3004 10526
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 2962 8800 3018 8809
rect 2962 8735 3018 8744
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2870 8120 2926 8129
rect 2870 8055 2872 8064
rect 2924 8055 2926 8064
rect 2872 8026 2924 8032
rect 3068 7970 3096 9862
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2884 7942 3096 7970
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7546 2820 7686
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2884 7410 2912 7942
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2596 7200 2648 7206
rect 2516 7160 2596 7188
rect 2596 7142 2648 7148
rect 2608 7018 2636 7142
rect 2608 6990 2728 7018
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2424 4282 2452 5170
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2516 3602 2544 4762
rect 2608 3602 2636 5238
rect 2700 4486 2728 6990
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2884 6322 2912 6938
rect 2976 6458 3004 7822
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 3068 7002 3096 7754
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3056 6656 3108 6662
rect 3054 6624 3056 6633
rect 3108 6624 3110 6633
rect 3054 6559 3110 6568
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2424 3194 2452 3334
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 1858 3088 1914 3097
rect 1914 3046 1992 3074
rect 1858 3023 1914 3032
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1872 800 1900 2926
rect 1964 2582 1992 3046
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 2228 2100 2280 2106
rect 2228 2042 2280 2048
rect 2240 800 2268 2042
rect 2596 1964 2648 1970
rect 2596 1906 2648 1912
rect 2608 800 2636 1906
rect 2700 1873 2728 4422
rect 2792 4214 2820 6190
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 4282 3004 4490
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2792 2281 2820 3470
rect 2976 3210 3004 4218
rect 3068 3913 3096 6559
rect 3160 5914 3188 8910
rect 3252 8906 3280 11766
rect 3344 9042 3372 12106
rect 3528 11642 3556 12406
rect 3988 12374 4016 12922
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3896 11665 3924 12310
rect 4080 11830 4108 12786
rect 4264 12782 4292 13212
rect 4356 13190 4384 13330
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 12306 4292 12582
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4252 12096 4304 12102
rect 4172 12056 4252 12084
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3436 11614 3556 11642
rect 3882 11656 3938 11665
rect 3436 9110 3464 11614
rect 3882 11591 3938 11600
rect 3976 11620 4028 11626
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3528 11150 3556 11290
rect 3896 11218 3924 11591
rect 3976 11562 4028 11568
rect 3988 11257 4016 11562
rect 3974 11248 4030 11257
rect 3884 11212 3936 11218
rect 3974 11183 4030 11192
rect 3884 11154 3936 11160
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 10674 3556 11086
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3436 8514 3464 9046
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3252 8498 3464 8514
rect 3240 8492 3464 8498
rect 3292 8486 3464 8492
rect 3240 8434 3292 8440
rect 3252 8022 3280 8434
rect 3528 8276 3556 8842
rect 3896 8401 3924 10202
rect 4080 10033 4108 10406
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9081 4016 9318
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3882 8392 3938 8401
rect 3882 8327 3938 8336
rect 3344 8248 3556 8276
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3252 6458 3280 7346
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3344 6202 3372 8248
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 7546 3648 7686
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3252 6174 3372 6202
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3252 5658 3280 6174
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5778 3372 6054
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3160 5630 3280 5658
rect 3054 3904 3110 3913
rect 3054 3839 3110 3848
rect 3160 3482 3188 5630
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5370 3280 5510
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3436 4706 3464 7210
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3792 6996 3844 7002
rect 3844 6956 3924 6984
rect 3792 6938 3844 6944
rect 3790 6896 3846 6905
rect 3516 6860 3568 6866
rect 3790 6831 3792 6840
rect 3516 6802 3568 6808
rect 3844 6831 3846 6840
rect 3792 6802 3844 6808
rect 3528 6254 3556 6802
rect 3790 6760 3846 6769
rect 3700 6724 3752 6730
rect 3790 6695 3846 6704
rect 3700 6666 3752 6672
rect 3606 6488 3662 6497
rect 3606 6423 3662 6432
rect 3620 6390 3648 6423
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3712 6254 3740 6666
rect 3804 6458 3832 6695
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3896 5273 3924 6956
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3344 4678 3464 4706
rect 3344 4146 3372 4678
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3602 3372 4082
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3160 3454 3280 3482
rect 3252 3398 3280 3454
rect 3884 3460 3936 3466
rect 3988 3448 4016 8910
rect 4080 8362 4108 9551
rect 4172 8498 4200 12056
rect 4252 12038 4304 12044
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4264 11354 4292 11766
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4264 11150 4292 11290
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10606 4292 11086
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4356 10146 4384 13126
rect 4448 11642 4476 17326
rect 4632 16998 4660 17496
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4632 16658 4660 16934
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4632 15706 4660 16594
rect 4724 16182 4752 18090
rect 4908 17746 4936 18838
rect 5000 18714 5028 22200
rect 5078 20632 5134 20641
rect 5078 20567 5134 20576
rect 5092 20534 5120 20567
rect 5080 20528 5132 20534
rect 5080 20470 5132 20476
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19854 5304 20198
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19378 5304 19790
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5000 18686 5120 18714
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4908 16046 4936 16730
rect 5000 16590 5028 17002
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4986 16144 5042 16153
rect 4986 16079 4988 16088
rect 5040 16079 5042 16088
rect 4988 16050 5040 16056
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4816 15366 4844 15914
rect 4908 15434 4936 15982
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14414 4568 14758
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12306 4568 13262
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4540 11830 4568 12242
rect 4632 12102 4660 13126
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4724 11898 4752 12854
rect 4816 12442 4844 15302
rect 4908 13852 4936 15370
rect 5000 15337 5028 16050
rect 4986 15328 5042 15337
rect 4986 15263 5042 15272
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 14278 5028 14418
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5000 14006 5028 14214
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4908 13824 5028 13852
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4908 12345 4936 12786
rect 4894 12336 4950 12345
rect 4894 12271 4950 12280
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4448 11614 4660 11642
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4540 10810 4568 11018
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4264 10118 4384 10146
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4160 7948 4212 7954
rect 4080 7002 4108 7919
rect 4160 7890 4212 7896
rect 4172 7206 4200 7890
rect 4264 7478 4292 10118
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9178 4384 9998
rect 4448 9722 4476 10542
rect 4540 10130 4568 10746
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9722 4568 9930
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4448 9602 4476 9658
rect 4448 9574 4568 9602
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4356 6610 4384 8978
rect 4448 8974 4476 9318
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4540 8634 4568 9574
rect 4632 8906 4660 11614
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4540 8430 4568 8570
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 8294 4568 8366
rect 4448 8266 4568 8294
rect 4448 7886 4476 8266
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4448 6798 4476 7414
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4264 6582 4384 6610
rect 4264 6372 4292 6582
rect 4436 6384 4488 6390
rect 4066 6352 4122 6361
rect 4264 6344 4384 6372
rect 4066 6287 4122 6296
rect 4080 6118 4108 6287
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5642 4108 5714
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4729 4108 5102
rect 4066 4720 4122 4729
rect 4066 4655 4122 4664
rect 4068 4480 4120 4486
rect 4172 4468 4200 5510
rect 4264 5370 4292 6122
rect 4356 5574 4384 6344
rect 4436 6326 4488 6332
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4448 5914 4476 6326
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4436 5772 4488 5778
rect 4540 5760 4568 6326
rect 4488 5732 4568 5760
rect 4436 5714 4488 5720
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4264 5234 4292 5306
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 4758 4292 5170
rect 4356 5030 4384 5510
rect 4448 5098 4476 5714
rect 4436 5092 4488 5098
rect 4436 5034 4488 5040
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4120 4440 4200 4468
rect 4252 4480 4304 4486
rect 4068 4422 4120 4428
rect 4252 4422 4304 4428
rect 4264 3738 4292 4422
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4160 3664 4212 3670
rect 3936 3420 4016 3448
rect 4080 3612 4160 3618
rect 4080 3606 4212 3612
rect 4080 3590 4200 3606
rect 3884 3402 3936 3408
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 2884 3182 3004 3210
rect 3160 3194 3188 3334
rect 3252 3194 3280 3334
rect 3148 3188 3200 3194
rect 2884 2922 2912 3182
rect 3148 3130 3200 3136
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2778 2272 2834 2281
rect 2778 2207 2834 2216
rect 2686 1864 2742 1873
rect 2686 1799 2742 1808
rect 2976 800 3004 3062
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3068 2650 3096 2994
rect 3528 2836 3556 3130
rect 3896 2854 3924 3402
rect 3436 2808 3556 2836
rect 3884 2848 3936 2854
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 3332 2032 3384 2038
rect 3332 1974 3384 1980
rect 3344 800 3372 1974
rect 3436 1465 3464 2808
rect 3884 2790 3936 2796
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 3712 800 3740 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3804 1902 3832 2042
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3896 649 3924 2790
rect 4080 2514 4108 3590
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4172 2446 4200 3470
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3988 898 4016 2042
rect 4356 1057 4384 4966
rect 4632 4826 4660 8434
rect 4724 8242 4752 11698
rect 4816 9042 4844 11834
rect 4908 11830 4936 12271
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 5000 11762 5028 13824
rect 5092 12889 5120 18686
rect 5184 18086 5212 19314
rect 5368 18850 5396 22200
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 20058 5488 20198
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5460 19378 5488 19994
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5552 19242 5580 20402
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5644 20058 5672 20334
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5632 19848 5684 19854
rect 5630 19816 5632 19825
rect 5684 19816 5686 19825
rect 5630 19751 5686 19760
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5736 18986 5764 22200
rect 6104 20788 6132 22200
rect 6472 20890 6500 22200
rect 6472 20862 6684 20890
rect 6012 20760 6132 20788
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5828 19514 5856 20538
rect 5906 20360 5962 20369
rect 5906 20295 5908 20304
rect 5960 20295 5962 20304
rect 5908 20266 5960 20272
rect 5816 19508 5868 19514
rect 6012 19496 6040 20760
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6460 19508 6512 19514
rect 6012 19468 6132 19496
rect 5816 19450 5868 19456
rect 5644 18958 5764 18986
rect 5368 18822 5488 18850
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17746 5212 18022
rect 5276 17882 5304 18226
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5184 16969 5212 17138
rect 5170 16960 5226 16969
rect 5170 16895 5226 16904
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5184 15502 5212 15982
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5078 12880 5134 12889
rect 5078 12815 5134 12824
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5092 11558 5120 12582
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 10742 5120 11494
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4896 9376 4948 9382
rect 4894 9344 4896 9353
rect 4948 9344 4950 9353
rect 4894 9279 4950 9288
rect 5000 9081 5028 9386
rect 5092 9382 5120 9658
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4986 9072 5042 9081
rect 4804 9036 4856 9042
rect 4986 9007 4988 9016
rect 4804 8978 4856 8984
rect 5040 9007 5042 9016
rect 5080 9036 5132 9042
rect 4988 8978 5040 8984
rect 5080 8978 5132 8984
rect 5092 8906 5120 8978
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4816 8634 4844 8774
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4804 8356 4856 8362
rect 4856 8316 4936 8344
rect 4804 8298 4856 8304
rect 4724 8214 4844 8242
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4724 7546 4752 7686
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4816 7324 4844 8214
rect 4908 7954 4936 8316
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7478 4936 7890
rect 5000 7886 5028 8774
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4896 7472 4948 7478
rect 4988 7472 5040 7478
rect 4896 7414 4948 7420
rect 4986 7440 4988 7449
rect 5040 7440 5042 7449
rect 5092 7410 5120 7686
rect 4986 7375 5042 7384
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4816 7296 4936 7324
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4724 5642 4752 6598
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4448 4078 4476 4762
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4448 3670 4476 4014
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4540 3602 4568 3878
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4342 1048 4398 1057
rect 4342 983 4398 992
rect 3988 870 4108 898
rect 4080 800 4108 870
rect 4448 800 4476 2994
rect 4540 2514 4568 3538
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4816 800 4844 7142
rect 4908 5166 4936 7296
rect 5092 6905 5120 7346
rect 5078 6896 5134 6905
rect 4988 6860 5040 6866
rect 5078 6831 5134 6840
rect 4988 6802 5040 6808
rect 5000 5574 5028 6802
rect 5184 6746 5212 14962
rect 5276 11778 5304 17478
rect 5368 17066 5396 18634
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5460 16969 5488 18822
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18358 5580 18770
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5552 17882 5580 18294
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5446 16960 5502 16969
rect 5446 16895 5502 16904
rect 5552 16250 5580 17478
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5540 15360 5592 15366
rect 5538 15328 5540 15337
rect 5592 15328 5594 15337
rect 5538 15263 5594 15272
rect 5644 15162 5672 18958
rect 5722 18864 5778 18873
rect 5722 18799 5724 18808
rect 5776 18799 5778 18808
rect 5724 18770 5776 18776
rect 5722 18728 5778 18737
rect 5722 18663 5778 18672
rect 5736 18630 5764 18663
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5828 17814 5856 19450
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5920 18834 5948 19246
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5920 18290 5948 18566
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 6012 17882 6040 19178
rect 6104 18737 6132 19468
rect 6460 19450 6512 19456
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6380 18834 6408 19178
rect 6472 19009 6500 19450
rect 6458 19000 6514 19009
rect 6458 18935 6514 18944
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6090 18728 6146 18737
rect 6472 18698 6500 18935
rect 6090 18663 6146 18672
rect 6460 18692 6512 18698
rect 6512 18652 6592 18680
rect 6460 18634 6512 18640
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6564 18408 6592 18652
rect 6472 18380 6592 18408
rect 6090 18320 6146 18329
rect 6090 18255 6146 18264
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 17354 5856 17478
rect 5736 17338 5856 17354
rect 5724 17332 5856 17338
rect 5776 17326 5856 17332
rect 5724 17274 5776 17280
rect 5920 17270 5948 17818
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5814 16960 5870 16969
rect 5814 16895 5870 16904
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5828 16674 5856 16895
rect 5920 16794 5948 17070
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 5736 16114 5764 16662
rect 5828 16646 5948 16674
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5828 16250 5856 16458
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15502 5764 16050
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5460 13530 5488 14894
rect 5552 14414 5580 14894
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14074 5580 14350
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5368 12850 5396 13330
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5460 12646 5488 13126
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5552 12288 5580 13126
rect 5644 12986 5672 14962
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 13530 5764 14554
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 13938 5856 14214
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 13394 5856 13874
rect 5816 13388 5868 13394
rect 5736 13348 5816 13376
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5630 12880 5686 12889
rect 5630 12815 5686 12824
rect 5460 12260 5580 12288
rect 5460 11898 5488 12260
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5276 11750 5488 11778
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 11082 5304 11290
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5262 9072 5318 9081
rect 5262 9007 5318 9016
rect 5276 6866 5304 9007
rect 5368 8906 5396 10678
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5354 8664 5410 8673
rect 5460 8650 5488 11750
rect 5552 11694 5580 12106
rect 5644 12073 5672 12815
rect 5736 12782 5764 13348
rect 5816 13330 5868 13336
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5630 12064 5686 12073
rect 5630 11999 5686 12008
rect 5828 11914 5856 13126
rect 5644 11886 5856 11914
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 11354 5580 11630
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5552 10198 5580 11290
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5552 8786 5580 9658
rect 5644 8922 5672 11886
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5828 11354 5856 11698
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5920 10690 5948 16646
rect 6012 15706 6040 17546
rect 6104 17524 6132 18255
rect 6472 17814 6500 18380
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6564 17882 6592 18226
rect 6656 18193 6684 20862
rect 6734 18864 6790 18873
rect 6734 18799 6790 18808
rect 6748 18290 6776 18799
rect 6840 18737 6868 22200
rect 6826 18728 6882 18737
rect 6826 18663 6882 18672
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18329 6868 18566
rect 6826 18320 6882 18329
rect 6736 18284 6788 18290
rect 6826 18255 6882 18264
rect 6736 18226 6788 18232
rect 6642 18184 6698 18193
rect 6642 18119 6698 18128
rect 6736 18148 6788 18154
rect 6788 18108 6868 18136
rect 6736 18090 6788 18096
rect 6642 18048 6698 18057
rect 6642 17983 6698 17992
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6460 17808 6512 17814
rect 6460 17750 6512 17756
rect 6564 17678 6592 17818
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6104 17496 6592 17524
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6092 17128 6144 17134
rect 6564 17082 6592 17496
rect 6092 17070 6144 17076
rect 6104 16726 6132 17070
rect 6472 17054 6592 17082
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6472 16522 6500 17054
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6380 15609 6408 15846
rect 6366 15600 6422 15609
rect 6366 15535 6422 15544
rect 6564 15434 6592 16934
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6380 14482 6408 14826
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6012 12918 6040 13806
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13394 6408 13670
rect 6564 13394 6592 14010
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6656 13190 6684 17983
rect 6840 17954 6868 18108
rect 6932 18057 6960 22222
rect 7116 22114 7144 22222
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8404 22222 8616 22250
rect 7208 22114 7236 22200
rect 7116 22086 7236 22114
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 20058 7144 20334
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7012 19984 7064 19990
rect 7012 19926 7064 19932
rect 7024 18766 7052 19926
rect 7116 19242 7144 19994
rect 7392 19922 7420 20198
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19514 7236 19654
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7104 19236 7156 19242
rect 7104 19178 7156 19184
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7116 18698 7144 19178
rect 7208 18970 7236 19314
rect 7300 18970 7328 19858
rect 7484 19825 7512 20198
rect 7470 19816 7526 19825
rect 7470 19751 7526 19760
rect 7484 19514 7512 19751
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 18222 7144 18634
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7012 18080 7064 18086
rect 6918 18048 6974 18057
rect 7208 18034 7236 18906
rect 7300 18222 7328 18906
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7064 18028 7236 18034
rect 7012 18022 7236 18028
rect 6918 17983 6974 17992
rect 7024 18006 7236 18022
rect 6748 17926 6868 17954
rect 6748 17882 6776 17926
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6734 17640 6790 17649
rect 6734 17575 6790 17584
rect 6748 14362 6776 17575
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 17105 6960 17138
rect 7024 17134 7052 18006
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7116 17270 7144 17682
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 7012 17128 7064 17134
rect 6918 17096 6974 17105
rect 7012 17070 7064 17076
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 6918 17031 6974 17040
rect 7024 16776 7052 17070
rect 6932 16748 7052 16776
rect 7104 16788 7156 16794
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16046 6868 16390
rect 6932 16182 6960 16748
rect 7104 16730 7156 16736
rect 7010 16688 7066 16697
rect 7010 16623 7012 16632
rect 7064 16623 7066 16632
rect 7012 16594 7064 16600
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15638 6868 15846
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6932 15570 6960 16118
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6826 15192 6882 15201
rect 6826 15127 6882 15136
rect 6920 15156 6972 15162
rect 6840 15026 6868 15127
rect 6920 15098 6972 15104
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6748 14334 6868 14362
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14074 6776 14214
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6840 13954 6868 14334
rect 6748 13926 6868 13954
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6748 13002 6776 13926
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 13394 6868 13806
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6826 13288 6882 13297
rect 6826 13223 6882 13232
rect 6564 12974 6776 13002
rect 6000 12912 6052 12918
rect 6000 12854 6052 12860
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12442 6040 12718
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6564 12238 6592 12974
rect 6840 12918 6868 13223
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6656 12374 6684 12786
rect 6736 12640 6788 12646
rect 6788 12600 6868 12628
rect 6736 12582 6788 12588
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6564 11218 6592 11630
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6012 10742 6040 10950
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6564 10810 6592 11154
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 5828 10662 5948 10690
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5736 9722 5764 10474
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5722 9480 5778 9489
rect 5722 9415 5778 9424
rect 5736 9042 5764 9415
rect 5828 9178 5856 10662
rect 6472 10606 6500 10678
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 5920 10062 5948 10542
rect 6564 10130 6592 10746
rect 6656 10266 6684 12038
rect 6748 11626 6776 12038
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6642 10160 6698 10169
rect 6552 10124 6604 10130
rect 6642 10095 6698 10104
rect 6552 10066 6604 10072
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6012 9654 6040 9998
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6550 9752 6606 9761
rect 6550 9687 6606 9696
rect 6564 9654 6592 9687
rect 6000 9648 6052 9654
rect 6552 9648 6604 9654
rect 6052 9608 6132 9636
rect 6000 9590 6052 9596
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5920 9353 5948 9454
rect 5906 9344 5962 9353
rect 5906 9279 5962 9288
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5644 8894 5764 8922
rect 5736 8838 5764 8894
rect 5724 8832 5776 8838
rect 5552 8758 5672 8786
rect 5724 8774 5776 8780
rect 5460 8622 5580 8650
rect 5354 8599 5356 8608
rect 5408 8599 5410 8608
rect 5356 8570 5408 8576
rect 5368 8430 5396 8570
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5460 7857 5488 8434
rect 5446 7848 5502 7857
rect 5356 7812 5408 7818
rect 5446 7783 5502 7792
rect 5356 7754 5408 7760
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5368 6798 5396 7754
rect 5552 7732 5580 8622
rect 5460 7704 5580 7732
rect 5356 6792 5408 6798
rect 5080 6724 5132 6730
rect 5184 6718 5304 6746
rect 5356 6734 5408 6740
rect 5080 6666 5132 6672
rect 5092 6633 5120 6666
rect 5276 6662 5304 6718
rect 5264 6656 5316 6662
rect 5078 6624 5134 6633
rect 5264 6598 5316 6604
rect 5078 6559 5134 6568
rect 5354 6488 5410 6497
rect 5354 6423 5410 6432
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 5234 5028 5510
rect 5078 5400 5134 5409
rect 5368 5370 5396 6423
rect 5078 5335 5134 5344
rect 5356 5364 5408 5370
rect 5092 5302 5120 5335
rect 5356 5306 5408 5312
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5172 5228 5224 5234
rect 5460 5216 5488 7704
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5552 5370 5580 5782
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5540 5228 5592 5234
rect 5460 5188 5540 5216
rect 5172 5170 5224 5176
rect 5540 5170 5592 5176
rect 4896 5160 4948 5166
rect 4894 5128 4896 5137
rect 4948 5128 4950 5137
rect 4950 5086 5028 5114
rect 4894 5063 4950 5072
rect 5000 4690 5028 5086
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4908 4214 4936 4626
rect 5078 4584 5134 4593
rect 5078 4519 5134 4528
rect 5092 4486 5120 4519
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4908 3602 4936 4150
rect 5092 4146 5120 4422
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5092 2446 5120 2790
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5184 800 5212 5170
rect 5552 4282 5580 5170
rect 5644 5012 5672 8758
rect 5736 8498 5764 8774
rect 5828 8634 5856 9114
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7721 5764 7754
rect 5722 7712 5778 7721
rect 5722 7647 5778 7656
rect 5816 7472 5868 7478
rect 5722 7440 5778 7449
rect 5816 7414 5868 7420
rect 5722 7375 5778 7384
rect 5736 6866 5764 7375
rect 5828 7313 5856 7414
rect 5920 7342 5948 8978
rect 6012 8566 6040 9454
rect 6104 9178 6132 9608
rect 6552 9590 6604 9596
rect 6564 9217 6592 9590
rect 6550 9208 6606 9217
rect 6092 9172 6144 9178
rect 6550 9143 6606 9152
rect 6092 9114 6144 9120
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6472 8838 6500 9046
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8616 6592 8978
rect 6380 8588 6592 8616
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6092 8424 6144 8430
rect 6090 8392 6092 8401
rect 6144 8392 6146 8401
rect 6090 8327 6146 8336
rect 6288 8022 6316 8434
rect 6380 8090 6408 8588
rect 6656 8548 6684 10095
rect 6840 10010 6868 12600
rect 6932 12170 6960 15098
rect 7024 14958 7052 16458
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14074 7052 14758
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7024 12918 7052 13738
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6932 10606 6960 11562
rect 7024 11121 7052 12038
rect 7010 11112 7066 11121
rect 7010 11047 7066 11056
rect 7024 11014 7052 11047
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7024 10198 7052 10542
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6472 8520 6684 8548
rect 6748 9982 6868 10010
rect 6920 9988 6972 9994
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6472 7732 6500 8520
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8090 6592 8298
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6748 7818 6776 9982
rect 6920 9930 6972 9936
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 8974 6868 9862
rect 6932 9382 6960 9930
rect 7010 9616 7066 9625
rect 7010 9551 7012 9560
rect 7064 9551 7066 9560
rect 7012 9522 7064 9528
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7024 9178 7052 9522
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6840 8514 6868 8774
rect 6840 8486 6960 8514
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6840 8090 6868 8327
rect 6932 8090 6960 8486
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6472 7704 6592 7732
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 5908 7336 5960 7342
rect 5814 7304 5870 7313
rect 5908 7278 5960 7284
rect 5814 7239 5870 7248
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5778 5764 6054
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5736 5166 5764 5714
rect 5828 5302 5856 6666
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5644 4984 5764 5012
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 3602 5672 4694
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5552 800 5580 3431
rect 5736 1426 5764 4984
rect 5920 4026 5948 6870
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6458 6760 6514 6769
rect 6458 6695 6514 6704
rect 6288 6662 6316 6695
rect 6472 6662 6500 6695
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 6322 6592 7704
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 6656 6730 6684 6831
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6656 6633 6684 6666
rect 6642 6624 6698 6633
rect 6642 6559 6698 6568
rect 6642 6488 6698 6497
rect 6642 6423 6698 6432
rect 6656 6390 6684 6423
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6182 6216 6238 6225
rect 6182 6151 6184 6160
rect 6236 6151 6238 6160
rect 6184 6122 6236 6128
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 5998 5808 6054 5817
rect 5998 5743 6000 5752
rect 6052 5743 6054 5752
rect 6000 5714 6052 5720
rect 6012 5114 6040 5714
rect 6380 5710 6408 6054
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6564 5642 6592 6258
rect 6748 5914 6776 7142
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6474 6868 6802
rect 6932 6644 6960 7890
rect 7024 7750 7052 8230
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7585 7052 7686
rect 7010 7576 7066 7585
rect 7010 7511 7066 7520
rect 7024 6798 7052 7511
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6932 6616 7052 6644
rect 6840 6446 6960 6474
rect 6932 6254 6960 6446
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6826 5944 6882 5953
rect 6736 5908 6788 5914
rect 6826 5879 6882 5888
rect 6736 5850 6788 5856
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6564 5370 6592 5578
rect 6840 5574 6868 5879
rect 6932 5778 6960 6190
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6642 5400 6698 5409
rect 6552 5364 6604 5370
rect 6642 5335 6698 5344
rect 6552 5306 6604 5312
rect 6552 5160 6604 5166
rect 6012 5086 6132 5114
rect 6656 5137 6684 5335
rect 6552 5102 6604 5108
rect 6642 5128 6698 5137
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4690 6040 4966
rect 6104 4826 6132 5086
rect 6564 5001 6592 5102
rect 6642 5063 6698 5072
rect 6550 4992 6606 5001
rect 6606 4950 6684 4978
rect 6550 4927 6606 4936
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6104 4468 6132 4626
rect 5828 3998 5948 4026
rect 6012 4440 6132 4468
rect 5828 2774 5856 3998
rect 6012 3942 6040 4440
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5908 3664 5960 3670
rect 5908 3606 5960 3612
rect 5920 3466 5948 3606
rect 6012 3602 6040 3878
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 6104 3505 6132 4014
rect 6196 3534 6224 4082
rect 6184 3528 6236 3534
rect 6090 3496 6146 3505
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 6012 3454 6090 3482
rect 5828 2746 5948 2774
rect 5920 2650 5948 2746
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5920 2038 5948 2314
rect 5908 2032 5960 2038
rect 5908 1974 5960 1980
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 6012 1034 6040 3454
rect 6184 3470 6236 3476
rect 6090 3431 6146 3440
rect 6104 3371 6132 3431
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6564 2922 6592 4218
rect 6656 4010 6684 4950
rect 6840 4128 6868 5510
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4282 6960 5102
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6920 4140 6972 4146
rect 6840 4100 6920 4128
rect 6920 4082 6972 4088
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6656 2378 6684 3062
rect 6920 2984 6972 2990
rect 6918 2952 6920 2961
rect 6972 2952 6974 2961
rect 6918 2887 6974 2896
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 6642 2272 6698 2281
rect 6148 2204 6456 2213
rect 6642 2207 6698 2216
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6276 1420 6328 1426
rect 6276 1362 6328 1368
rect 5920 1006 6040 1034
rect 5920 800 5948 1006
rect 6288 800 6316 1362
rect 6656 800 6684 2207
rect 7024 800 7052 6616
rect 7116 4826 7144 16730
rect 7208 12322 7236 17070
rect 7300 16590 7328 17274
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7300 16425 7328 16526
rect 7286 16416 7342 16425
rect 7286 16351 7342 16360
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7300 16017 7328 16186
rect 7286 16008 7342 16017
rect 7286 15943 7342 15952
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 14890 7328 15506
rect 7392 15502 7420 18566
rect 7484 18290 7512 18634
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16658 7512 17002
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7484 16046 7512 16594
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7392 14890 7420 15438
rect 7484 15162 7512 15642
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7300 14414 7328 14826
rect 7576 14770 7604 22200
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7668 17202 7696 19994
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7760 19446 7788 19790
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7838 18728 7894 18737
rect 7838 18663 7894 18672
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7656 16992 7708 16998
rect 7654 16960 7656 16969
rect 7708 16960 7710 16969
rect 7654 16895 7710 16904
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15706 7696 15846
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7852 15042 7880 18663
rect 7944 16794 7972 22200
rect 8312 22114 8340 22200
rect 8404 22114 8432 22222
rect 8312 22086 8432 22114
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8312 19174 8340 20402
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8036 18902 8064 19110
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 8036 18358 8064 18702
rect 8404 18426 8432 19654
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8496 18970 8524 19246
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8312 17746 8340 18158
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8036 16794 8064 17478
rect 8220 17338 8248 17478
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8114 17232 8170 17241
rect 8404 17218 8432 18022
rect 8496 17814 8524 18226
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8588 17649 8616 22222
rect 8666 22200 8722 23000
rect 8772 22222 8984 22250
rect 8680 22114 8708 22200
rect 8772 22114 8800 22222
rect 8680 22086 8800 22114
rect 8956 20346 8984 22222
rect 9034 22200 9090 23000
rect 9140 22222 9352 22250
rect 9048 22114 9076 22200
rect 9140 22114 9168 22222
rect 9048 22086 9168 22114
rect 8956 20318 9260 20346
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8680 19514 8708 19858
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8680 18834 8708 19450
rect 8772 19446 8800 19654
rect 8760 19440 8812 19446
rect 9048 19417 9076 19790
rect 8760 19382 8812 19388
rect 9034 19408 9090 19417
rect 9034 19343 9090 19352
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8574 17640 8630 17649
rect 8574 17575 8630 17584
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8114 17167 8170 17176
rect 8312 17190 8432 17218
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7576 14742 7696 14770
rect 7562 14648 7618 14657
rect 7562 14583 7618 14592
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 13938 7328 14350
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7300 12986 7328 13874
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7392 13258 7420 13466
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7392 13161 7420 13194
rect 7378 13152 7434 13161
rect 7378 13087 7434 13096
rect 7484 12986 7512 13262
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7300 12442 7328 12922
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7208 12294 7420 12322
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10810 7236 10950
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7300 10010 7328 12174
rect 7392 10418 7420 12294
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10538 7512 11018
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7392 10390 7512 10418
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7208 9982 7328 10010
rect 7208 7834 7236 9982
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7300 9178 7328 9862
rect 7392 9518 7420 10066
rect 7484 9874 7512 10390
rect 7576 9994 7604 14583
rect 7668 12442 7696 14742
rect 7760 14618 7788 15030
rect 7852 15014 7972 15042
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7852 14346 7880 14894
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7746 13424 7802 13433
rect 7746 13359 7748 13368
rect 7800 13359 7802 13368
rect 7748 13330 7800 13336
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7760 12434 7788 12786
rect 7852 12782 7880 14282
rect 7944 13190 7972 15014
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7930 12880 7986 12889
rect 7930 12815 7986 12824
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7760 12406 7880 12434
rect 7668 11898 7696 12378
rect 7760 12306 7788 12406
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 11694 7788 12106
rect 7748 11688 7800 11694
rect 7746 11656 7748 11665
rect 7800 11656 7802 11665
rect 7746 11591 7802 11600
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7484 9846 7604 9874
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 7954 7328 8978
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8294 7420 8910
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 8022 7420 8230
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7208 7806 7328 7834
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 7449 7236 7686
rect 7194 7440 7250 7449
rect 7194 7375 7250 7384
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7208 6730 7236 6870
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7300 5710 7328 7806
rect 7392 7478 7420 7958
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6254 7420 6802
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7116 4690 7144 4762
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 2990 7144 3878
rect 7208 3058 7236 5510
rect 7300 5370 7328 5646
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 4690 7328 5102
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7300 4282 7328 4626
rect 7392 4570 7420 6190
rect 7484 4758 7512 9454
rect 7576 7585 7604 9846
rect 7562 7576 7618 7585
rect 7562 7511 7618 7520
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7576 6934 7604 7346
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 5710 7604 6598
rect 7668 6322 7696 10406
rect 7746 9616 7802 9625
rect 7746 9551 7802 9560
rect 7760 9382 7788 9551
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 8022 7788 9318
rect 7852 9058 7880 12406
rect 7944 11558 7972 12815
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8036 11082 8064 16594
rect 8128 15722 8156 17167
rect 8312 16998 8340 17190
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16674 8340 16934
rect 8220 16658 8340 16674
rect 8208 16652 8340 16658
rect 8260 16646 8340 16652
rect 8208 16594 8260 16600
rect 8404 16590 8432 17070
rect 8588 16794 8616 17478
rect 8680 17338 8708 18158
rect 9048 18154 9076 18566
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9140 17814 9168 17845
rect 9128 17808 9180 17814
rect 9126 17776 9128 17785
rect 9180 17776 9182 17785
rect 9126 17711 9182 17720
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8772 17048 8800 17478
rect 9140 17338 9168 17711
rect 9232 17354 9260 20318
rect 9324 18737 9352 22222
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 21546 22200 21602 23000
rect 21652 22222 21864 22250
rect 9310 18728 9366 18737
rect 9310 18663 9366 18672
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 17882 9352 18566
rect 9416 18193 9444 22200
rect 9600 18970 9720 18986
rect 9588 18964 9720 18970
rect 9640 18958 9720 18964
rect 9588 18906 9640 18912
rect 9692 18630 9720 18958
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9588 18216 9640 18222
rect 9402 18184 9458 18193
rect 9588 18158 9640 18164
rect 9402 18119 9458 18128
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9128 17332 9180 17338
rect 9232 17326 9352 17354
rect 9128 17274 9180 17280
rect 8680 17020 8800 17048
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8128 15694 8340 15722
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8128 14414 8156 15098
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8114 14240 8170 14249
rect 8114 14175 8170 14184
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8036 10266 8064 10542
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7852 9030 8064 9058
rect 8036 8945 8064 9030
rect 8022 8936 8078 8945
rect 8022 8871 8078 8880
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7760 6798 7788 7686
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7746 6624 7802 6633
rect 7746 6559 7802 6568
rect 7760 6390 7788 6559
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 5778 7696 6054
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 7576 4690 7604 5238
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7392 4542 7512 4570
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7392 3194 7420 4422
rect 7484 3398 7512 4542
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7378 3088 7434 3097
rect 7196 3052 7248 3058
rect 7378 3023 7434 3032
rect 7196 2994 7248 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7208 2310 7236 2518
rect 7300 2514 7328 2926
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7116 2038 7144 2246
rect 7208 2106 7236 2246
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 7392 800 7420 3023
rect 7484 2990 7512 3334
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7576 2650 7604 4422
rect 7668 3126 7696 4966
rect 7852 4622 7880 5306
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7852 2650 7880 4422
rect 7944 4214 7972 4626
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 8036 3482 8064 8871
rect 8128 6458 8156 14175
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12306 8248 13262
rect 8312 12986 8340 15694
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8404 14958 8432 15574
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8496 14249 8524 16662
rect 8680 14929 8708 17020
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15162 9168 16050
rect 9232 15638 9260 16118
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8666 14920 8722 14929
rect 8666 14855 8722 14864
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14414 8708 14758
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9232 14482 9260 15370
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8482 14240 8538 14249
rect 8482 14175 8538 14184
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13433 8432 13670
rect 8390 13424 8446 13433
rect 8390 13359 8446 13368
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8312 12306 8340 12922
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8220 11354 8248 12242
rect 8312 11937 8340 12242
rect 8298 11928 8354 11937
rect 8298 11863 8354 11872
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8206 11112 8262 11121
rect 8206 11047 8262 11056
rect 8220 10198 8248 11047
rect 8312 11014 8340 11766
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8208 10192 8260 10198
rect 8206 10160 8208 10169
rect 8260 10160 8262 10169
rect 8206 10095 8262 10104
rect 8312 9722 8340 10610
rect 8404 10470 8432 13359
rect 8680 12434 8708 14350
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 14113 8984 14214
rect 8942 14104 8998 14113
rect 8942 14039 8998 14048
rect 9218 14104 9274 14113
rect 9218 14039 9274 14048
rect 9232 14006 9260 14039
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9128 13728 9180 13734
rect 9220 13728 9272 13734
rect 9128 13670 9180 13676
rect 9218 13696 9220 13705
rect 9272 13696 9274 13705
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12646 9076 13126
rect 9140 12986 9168 13670
rect 9218 13631 9274 13640
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12782 9260 13330
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8680 12406 9168 12434
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8574 11792 8630 11801
rect 8574 11727 8576 11736
rect 8628 11727 8630 11736
rect 8576 11698 8628 11704
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8588 10674 8616 11154
rect 8680 11150 8708 11834
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8588 10130 8616 10610
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 10124 8628 10130
rect 8576 10066 8628 10072
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8220 8673 8248 8842
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 7970 8248 8434
rect 8312 8090 8340 9454
rect 8404 9178 8432 9862
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8566 8432 8774
rect 8496 8634 8524 9862
rect 8588 9722 8616 10066
rect 8680 9897 8708 10406
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9048 9994 9076 10202
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8666 9888 8722 9897
rect 8666 9823 8722 9832
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8680 9110 8708 9590
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9140 9178 9168 12406
rect 9324 11778 9352 17326
rect 9416 16794 9444 17818
rect 9508 17746 9536 18090
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9508 17134 9536 17682
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9416 15162 9444 16730
rect 9600 16561 9628 18158
rect 9692 17134 9720 18566
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9586 16552 9642 16561
rect 9586 16487 9642 16496
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16250 9536 16390
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9588 16244 9640 16250
rect 9692 16232 9720 17070
rect 9640 16204 9720 16232
rect 9588 16186 9640 16192
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9416 14906 9444 15098
rect 9600 15065 9628 15098
rect 9586 15056 9642 15065
rect 9586 14991 9642 15000
rect 9588 14952 9640 14958
rect 9416 14878 9536 14906
rect 9588 14894 9640 14900
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14482 9444 14758
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9508 14362 9536 14878
rect 9600 14550 9628 14894
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9416 14334 9536 14362
rect 9588 14408 9640 14414
rect 9784 14396 9812 22200
rect 10152 19334 10180 22200
rect 10520 20618 10548 22200
rect 9968 19306 10180 19334
rect 10336 20590 10548 20618
rect 10888 20602 10916 22200
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10876 20596 10928 20602
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 14618 9904 16390
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9640 14368 9812 14396
rect 9588 14350 9640 14356
rect 9416 12102 9444 14334
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9494 13968 9550 13977
rect 9494 13903 9550 13912
rect 9508 13870 9536 13903
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9494 13696 9550 13705
rect 9600 13682 9628 13806
rect 9550 13654 9628 13682
rect 9494 13631 9550 13640
rect 9600 13326 9628 13654
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 12434 9536 12786
rect 9600 12782 9628 13262
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9508 12406 9628 12434
rect 9600 12102 9628 12406
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9416 11937 9444 12038
rect 9402 11928 9458 11937
rect 9402 11863 9458 11872
rect 9324 11750 9536 11778
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9232 11150 9260 11630
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9232 10810 9260 11086
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9218 10296 9274 10305
rect 9324 10266 9352 11494
rect 9416 11354 9444 11630
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9218 10231 9220 10240
rect 9272 10231 9274 10240
rect 9312 10260 9364 10266
rect 9220 10202 9272 10208
rect 9312 10202 9364 10208
rect 9416 10146 9444 10678
rect 9232 10118 9444 10146
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8673 8708 8842
rect 8666 8664 8722 8673
rect 8484 8628 8536 8634
rect 9140 8634 9168 9114
rect 8666 8599 8722 8608
rect 9128 8628 9180 8634
rect 8484 8570 8536 8576
rect 9128 8570 9180 8576
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8220 7942 8340 7970
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 6866 8248 7686
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8312 6848 8340 7942
rect 8404 7886 8432 8502
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7886 8524 8230
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 6860 8444 6866
rect 8312 6820 8392 6848
rect 8312 6662 8340 6820
rect 8392 6802 8444 6808
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8390 6624 8446 6633
rect 8390 6559 8446 6568
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8128 5778 8156 6190
rect 8404 5817 8432 6559
rect 8390 5808 8446 5817
rect 8116 5772 8168 5778
rect 8390 5743 8446 5752
rect 8116 5714 8168 5720
rect 8128 4690 8156 5714
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8206 5128 8262 5137
rect 8206 5063 8262 5072
rect 8220 4826 8248 5063
rect 8312 5030 8340 5646
rect 8404 5574 8432 5743
rect 8496 5710 8524 7822
rect 8588 7478 8616 7890
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5370 8524 5510
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8404 4826 8432 5170
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8116 4684 8168 4690
rect 8392 4684 8444 4690
rect 8168 4644 8248 4672
rect 8116 4626 8168 4632
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 7944 3454 8064 3482
rect 7944 2774 7972 3454
rect 8024 2984 8076 2990
rect 8022 2952 8024 2961
rect 8076 2952 8078 2961
rect 8022 2887 8078 2896
rect 7944 2746 8064 2774
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7760 870 7880 898
rect 7760 800 7788 870
rect 3882 640 3938 649
rect 3882 575 3938 584
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 7852 762 7880 870
rect 8036 762 8064 2746
rect 8128 800 8156 3975
rect 8220 3602 8248 4644
rect 8392 4626 8444 4632
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8312 3534 8340 3878
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8404 2446 8432 4626
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8496 2446 8524 4490
rect 8588 4282 8616 6054
rect 8680 5846 8708 7346
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9140 7002 9168 7210
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8956 6769 8984 6802
rect 8758 6760 8814 6769
rect 8942 6760 8998 6769
rect 8814 6718 8892 6746
rect 8758 6695 8814 6704
rect 8864 6662 8892 6718
rect 8942 6695 8998 6704
rect 9140 6662 9168 6802
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8852 6656 8904 6662
rect 9128 6656 9180 6662
rect 8852 6598 8904 6604
rect 8942 6624 8998 6633
rect 8772 6458 8800 6598
rect 9128 6598 9180 6604
rect 8942 6559 8998 6568
rect 8956 6458 8984 6559
rect 9126 6488 9182 6497
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8944 6452 8996 6458
rect 9126 6423 9128 6432
rect 8944 6394 8996 6400
rect 9180 6423 9182 6432
rect 9128 6394 9180 6400
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9126 5944 9182 5953
rect 9126 5879 9128 5888
rect 9180 5879 9182 5888
rect 9128 5850 9180 5856
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8680 5234 8708 5782
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8772 5166 8800 5646
rect 8864 5302 8892 5714
rect 9232 5681 9260 10118
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9310 9208 9366 9217
rect 9310 9143 9366 9152
rect 9218 5672 9274 5681
rect 9218 5607 9274 5616
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8944 5228 8996 5234
rect 8996 5188 9168 5216
rect 8944 5170 8996 5176
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8680 4282 8708 5034
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8760 4752 8812 4758
rect 8760 4694 8812 4700
rect 8772 4554 8800 4694
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8864 4185 8892 4490
rect 9140 4282 9168 5188
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8850 4176 8906 4185
rect 8668 4140 8720 4146
rect 8850 4111 8906 4120
rect 9036 4140 9088 4146
rect 8668 4082 8720 4088
rect 9036 4082 9088 4088
rect 8680 3738 8708 4082
rect 9048 4049 9076 4082
rect 9034 4040 9090 4049
rect 9034 3975 9090 3984
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 9036 3528 9088 3534
rect 9140 3516 9168 4218
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9088 3488 9168 3516
rect 9036 3470 9088 3476
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8588 3194 8616 3402
rect 9036 3392 9088 3398
rect 9088 3352 9168 3380
rect 9036 3334 9088 3340
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9140 2650 9168 3352
rect 9232 3194 9260 3946
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9324 3074 9352 9143
rect 9416 8294 9444 9318
rect 9508 8566 9536 11750
rect 9600 10742 9628 12038
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9588 10464 9640 10470
rect 9692 10452 9720 14214
rect 9784 13841 9812 14368
rect 9876 14074 9904 14418
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9864 13864 9916 13870
rect 9770 13832 9826 13841
rect 9864 13806 9916 13812
rect 9770 13767 9826 13776
rect 9876 13433 9904 13806
rect 9862 13424 9918 13433
rect 9862 13359 9918 13368
rect 9968 12986 9996 19306
rect 10046 18728 10102 18737
rect 10046 18663 10102 18672
rect 10060 18426 10088 18663
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10336 18057 10364 20590
rect 10876 20538 10928 20544
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10428 19514 10456 20402
rect 10520 19786 10548 20402
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 19961 10640 20266
rect 10980 19972 11008 20946
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11060 19984 11112 19990
rect 10598 19952 10654 19961
rect 10980 19944 11060 19972
rect 11060 19926 11112 19932
rect 11164 19922 11192 20198
rect 10598 19887 10654 19896
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 10508 19780 10560 19786
rect 10508 19722 10560 19728
rect 10600 19780 10652 19786
rect 10784 19780 10836 19786
rect 10652 19740 10732 19768
rect 10600 19722 10652 19728
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10612 18970 10640 19314
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10704 18630 10732 19740
rect 10784 19722 10836 19728
rect 10796 19310 10824 19722
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10888 18834 10916 19314
rect 10980 18970 11008 19382
rect 11072 19334 11100 19790
rect 11164 19394 11192 19858
rect 11256 19514 11284 22200
rect 11624 20890 11652 22200
rect 11624 20862 11744 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11532 19854 11560 20402
rect 11716 20330 11744 20862
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11992 20058 12020 22200
rect 12360 20602 12388 22200
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11716 19718 11744 19790
rect 11808 19718 11836 19994
rect 12084 19786 12112 20334
rect 12728 19990 12756 22200
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12716 19984 12768 19990
rect 12716 19926 12768 19932
rect 13004 19854 13032 20198
rect 13096 20058 13124 22200
rect 13084 20052 13136 20058
rect 13464 20040 13492 22200
rect 13544 20052 13596 20058
rect 13464 20012 13544 20040
rect 13084 19994 13136 20000
rect 13544 19994 13596 20000
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11164 19378 11284 19394
rect 11164 19372 11296 19378
rect 11164 19366 11244 19372
rect 11072 19306 11192 19334
rect 11244 19314 11296 19320
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18426 10916 18566
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10874 18320 10930 18329
rect 10874 18255 10930 18264
rect 10322 18048 10378 18057
rect 10322 17983 10378 17992
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 17338 10272 17682
rect 10692 17604 10744 17610
rect 10692 17546 10744 17552
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10060 16182 10088 16594
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10060 14482 10088 14826
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 10060 14006 10088 14039
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9876 12753 9904 12786
rect 9862 12744 9918 12753
rect 9862 12679 9918 12688
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 10810 9812 11698
rect 9968 11694 9996 12310
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9772 10464 9824 10470
rect 9692 10424 9772 10452
rect 9588 10406 9640 10412
rect 9772 10406 9824 10412
rect 9600 10130 9628 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9772 10124 9824 10130
rect 9876 10112 9904 11494
rect 9968 11082 9996 11630
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9824 10084 9904 10112
rect 9772 10066 9824 10072
rect 9968 10044 9996 10406
rect 10060 10062 10088 13942
rect 10152 12782 10180 16526
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10198 10180 10950
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 9876 10016 9996 10044
rect 10048 10056 10100 10062
rect 9876 9674 9904 10016
rect 10048 9998 10100 10004
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 9674 10088 9862
rect 9692 9646 9904 9674
rect 9968 9646 10088 9674
rect 9692 9110 9720 9646
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9600 8430 9628 8978
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9784 8634 9812 8842
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9402 7984 9458 7993
rect 9600 7954 9628 8366
rect 9784 7954 9812 8570
rect 9402 7919 9404 7928
rect 9456 7919 9458 7928
rect 9588 7948 9640 7954
rect 9404 7890 9456 7896
rect 9588 7890 9640 7896
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9862 7848 9918 7857
rect 9862 7783 9918 7792
rect 9876 7750 9904 7783
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9876 7478 9904 7686
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9416 6798 9444 7346
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 4758 9444 6598
rect 9508 6390 9536 7142
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9600 6254 9628 6870
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9692 6361 9720 6802
rect 9678 6352 9734 6361
rect 9678 6287 9734 6296
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5234 9536 5646
rect 9600 5642 9628 6054
rect 9678 5672 9734 5681
rect 9588 5636 9640 5642
rect 9678 5607 9734 5616
rect 9588 5578 9640 5584
rect 9600 5370 9628 5578
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9692 5250 9720 5607
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9600 5222 9720 5250
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9416 4622 9444 4694
rect 9508 4690 9536 5170
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9600 4468 9628 5222
rect 9784 4826 9812 6190
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4729 9904 5238
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9862 4584 9918 4593
rect 9862 4519 9918 4528
rect 9232 3046 9352 3074
rect 9416 4440 9628 4468
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8850 2544 8906 2553
rect 8850 2479 8906 2488
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8496 2310 8524 2382
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8496 1970 8524 2246
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8588 1902 8616 2246
rect 8576 1896 8628 1902
rect 8576 1838 8628 1844
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8496 800 8524 1498
rect 8864 800 8892 2479
rect 9232 1562 9260 3046
rect 9416 2774 9444 4440
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9508 3058 9536 3470
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9600 2938 9628 4082
rect 9692 3913 9720 4150
rect 9678 3904 9734 3913
rect 9678 3839 9734 3848
rect 9876 3641 9904 4519
rect 9862 3632 9918 3641
rect 9862 3567 9918 3576
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9324 2746 9444 2774
rect 9508 2910 9628 2938
rect 9784 2922 9812 3402
rect 9772 2916 9824 2922
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 9324 1442 9352 2746
rect 9232 1414 9352 1442
rect 9232 800 9260 1414
rect 9508 1034 9536 2910
rect 9772 2858 9824 2864
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 2514 9628 2790
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9876 1442 9904 3567
rect 9968 2446 9996 9646
rect 10138 9344 10194 9353
rect 10138 9279 10194 9288
rect 10046 8800 10102 8809
rect 10046 8735 10102 8744
rect 10060 6390 10088 8735
rect 10152 7721 10180 9279
rect 10244 7857 10272 17274
rect 10704 17202 10732 17546
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14074 10364 14418
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10322 13832 10378 13841
rect 10322 13767 10378 13776
rect 10336 13462 10364 13767
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10324 10736 10376 10742
rect 10322 10704 10324 10713
rect 10376 10704 10378 10713
rect 10322 10639 10378 10648
rect 10428 10577 10456 15030
rect 10520 14414 10548 15438
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10612 14958 10640 15370
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10612 13870 10640 14894
rect 10704 14346 10732 16118
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15502 10824 15846
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10888 15366 10916 18255
rect 10980 18222 11008 18906
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10980 17746 11008 18158
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 11072 16810 11100 17478
rect 10980 16782 11100 16810
rect 10980 16522 11008 16782
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 11072 15042 11100 16526
rect 11164 16114 11192 19306
rect 11716 18850 11744 19654
rect 12808 19168 12860 19174
rect 12806 19136 12808 19145
rect 12860 19136 12862 19145
rect 12806 19071 12862 19080
rect 12912 18970 12940 19790
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 11624 18822 11744 18850
rect 11624 18612 11652 18822
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11256 18584 11652 18612
rect 11256 17218 11284 18584
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11716 18358 11744 18634
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11612 18080 11664 18086
rect 11610 18048 11612 18057
rect 11664 18048 11666 18057
rect 11610 17983 11666 17992
rect 11716 17746 11744 18294
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11612 17332 11664 17338
rect 11716 17320 11744 17682
rect 11808 17338 11836 18906
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11900 17542 11928 18158
rect 11992 18154 12020 18634
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12254 18456 12310 18465
rect 12254 18391 12256 18400
rect 12308 18391 12310 18400
rect 12256 18362 12308 18368
rect 12162 18320 12218 18329
rect 12162 18255 12164 18264
rect 12216 18255 12218 18264
rect 12164 18226 12216 18232
rect 12348 18216 12400 18222
rect 12070 18184 12126 18193
rect 11980 18148 12032 18154
rect 12348 18158 12400 18164
rect 12070 18119 12126 18128
rect 11980 18090 12032 18096
rect 12084 17882 12112 18119
rect 12360 17882 12388 18158
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12544 17728 12572 18566
rect 12452 17700 12572 17728
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11664 17292 11744 17320
rect 11796 17332 11848 17338
rect 11612 17274 11664 17280
rect 11796 17274 11848 17280
rect 11256 17190 11376 17218
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11256 15162 11284 16662
rect 11348 16561 11376 17190
rect 11624 16658 11652 17274
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11334 16552 11390 16561
rect 11334 16487 11390 16496
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11072 15014 11284 15042
rect 11060 14952 11112 14958
rect 11058 14920 11060 14929
rect 11112 14920 11114 14929
rect 11058 14855 11114 14864
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13870 10916 14214
rect 10966 13968 11022 13977
rect 10966 13903 11022 13912
rect 10600 13864 10652 13870
rect 10876 13864 10928 13870
rect 10600 13806 10652 13812
rect 10874 13832 10876 13841
rect 10928 13832 10930 13841
rect 10874 13767 10930 13776
rect 10980 13734 11008 13903
rect 11072 13870 11100 14282
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11256 13802 11284 15014
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11244 13796 11296 13802
rect 11244 13738 11296 13744
rect 10968 13728 11020 13734
rect 11348 13682 11376 14010
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11532 13841 11560 13874
rect 11518 13832 11574 13841
rect 11518 13767 11574 13776
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 10968 13670 11020 13676
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12646 10640 13194
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12714 10732 13126
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12481 10640 12582
rect 10598 12472 10654 12481
rect 10598 12407 10654 12416
rect 10690 12336 10746 12345
rect 10690 12271 10746 12280
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10520 11014 10548 11698
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10810 10640 10950
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10600 10600 10652 10606
rect 10414 10568 10470 10577
rect 10600 10542 10652 10548
rect 10414 10503 10470 10512
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10130 10364 10406
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10428 9654 10456 10503
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10520 9897 10548 10066
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 10612 9722 10640 10542
rect 10704 9761 10732 12271
rect 10980 11132 11008 13670
rect 11256 13654 11376 13682
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11164 13190 11192 13262
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12850 11192 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12238 11192 12786
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11072 11626 11100 12038
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11060 11144 11112 11150
rect 10980 11104 11060 11132
rect 11060 11086 11112 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10796 10810 10824 11018
rect 11164 10962 11192 12038
rect 11256 11898 11284 13654
rect 11624 13546 11652 13738
rect 11716 13682 11744 16730
rect 11808 16454 11836 17070
rect 11900 16794 11928 17478
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12176 17082 12204 17206
rect 12084 17066 12204 17082
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12072 17060 12204 17066
rect 12124 17054 12204 17060
rect 12072 17002 12124 17008
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11978 16552 12034 16561
rect 11978 16487 12034 16496
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 13870 11836 16390
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11900 15162 11928 15302
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14618 11928 14962
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11716 13654 11836 13682
rect 11624 13518 11744 13546
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11072 10934 11192 10962
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 10470 10824 10746
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 10968 10668 11020 10674
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10690 9752 10746 9761
rect 10600 9716 10652 9722
rect 10796 9722 10824 10134
rect 10690 9687 10746 9696
rect 10784 9716 10836 9722
rect 10600 9658 10652 9664
rect 10784 9658 10836 9664
rect 10416 9648 10468 9654
rect 10322 9616 10378 9625
rect 10888 9602 10916 10639
rect 10968 10610 11020 10616
rect 10980 10198 11008 10610
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 11072 9674 11100 10934
rect 10416 9590 10468 9596
rect 10322 9551 10378 9560
rect 10704 9574 10916 9602
rect 10980 9646 11100 9674
rect 10230 7848 10286 7857
rect 10230 7783 10286 7792
rect 10138 7712 10194 7721
rect 10138 7647 10194 7656
rect 10152 7426 10180 7647
rect 10244 7546 10272 7783
rect 10336 7750 10364 9551
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 9178 10548 9454
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10520 8566 10548 9114
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10414 8256 10470 8265
rect 10414 8191 10470 8200
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10336 7478 10364 7686
rect 10324 7472 10376 7478
rect 10152 7398 10272 7426
rect 10324 7414 10376 7420
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10138 6080 10194 6089
rect 10060 4146 10088 6054
rect 10138 6015 10194 6024
rect 10152 5642 10180 6015
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4622 10180 4966
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10244 2774 10272 7398
rect 10428 7324 10456 8191
rect 10520 8129 10548 8502
rect 10506 8120 10562 8129
rect 10506 8055 10562 8064
rect 10612 7886 10640 9318
rect 10704 8022 10732 9574
rect 10980 8242 11008 9646
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10888 8214 11008 8242
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10336 7296 10456 7324
rect 10336 5914 10364 7296
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6186 10456 6666
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 5574 10456 6122
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10336 5166 10364 5306
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10428 4690 10456 5510
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10416 4480 10468 4486
rect 10322 4448 10378 4457
rect 10416 4422 10468 4428
rect 10322 4383 10378 4392
rect 10336 3942 10364 4383
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3641 10364 3878
rect 10428 3670 10456 4422
rect 10416 3664 10468 3670
rect 10322 3632 10378 3641
rect 10416 3606 10468 3612
rect 10322 3567 10378 3576
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10336 3126 10364 3334
rect 10520 3126 10548 7686
rect 10704 7546 10732 7958
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10888 6497 10916 8214
rect 10966 8120 11022 8129
rect 10966 8055 11022 8064
rect 10980 7954 11008 8055
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7206 11008 7346
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6866 11008 7142
rect 11072 6934 11100 8434
rect 11164 8294 11192 8910
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7478 11192 8230
rect 11256 7478 11284 11834
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 11348 11218 11376 11562
rect 11440 11354 11468 11834
rect 11520 11756 11572 11762
rect 11716 11744 11744 13518
rect 11572 11716 11744 11744
rect 11520 11698 11572 11704
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11348 10130 11376 10542
rect 11716 10470 11744 10950
rect 11808 10742 11836 13654
rect 11992 12434 12020 16487
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12084 13938 12112 15438
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12176 13734 12204 16934
rect 12360 16810 12388 17070
rect 12452 16946 12480 17700
rect 12636 17626 12664 18566
rect 12820 18290 12848 18770
rect 13004 18329 13032 19790
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 13188 19378 13216 19722
rect 13832 19514 13860 22200
rect 14200 20346 14228 22200
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14200 20318 14320 20346
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14292 20058 14320 20318
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19938 14412 20402
rect 14292 19910 14412 19938
rect 14292 19854 14320 19910
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13096 18902 13124 19246
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13096 18358 13124 18838
rect 13556 18834 13584 19178
rect 13636 19168 13688 19174
rect 13634 19136 13636 19145
rect 13688 19136 13690 19145
rect 13634 19071 13690 19080
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13084 18352 13136 18358
rect 12990 18320 13046 18329
rect 12808 18284 12860 18290
rect 13084 18294 13136 18300
rect 12990 18255 13046 18264
rect 12808 18226 12860 18232
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12728 17678 12756 18158
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12544 17610 12664 17626
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12532 17604 12664 17610
rect 12584 17598 12664 17604
rect 12532 17546 12584 17552
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17241 12756 17478
rect 12714 17232 12770 17241
rect 12714 17167 12770 17176
rect 12820 17134 12848 17682
rect 13096 17678 13124 18294
rect 13372 17814 13400 18566
rect 13556 18358 13584 18770
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17338 13032 17546
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 12808 17128 12860 17134
rect 12544 17066 12664 17082
rect 12808 17070 12860 17076
rect 12532 17060 12664 17066
rect 12584 17054 12664 17060
rect 12532 17002 12584 17008
rect 12452 16918 12572 16946
rect 12360 16782 12480 16810
rect 12348 16040 12400 16046
rect 12452 16028 12480 16782
rect 12544 16250 12572 16918
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12400 16000 12480 16028
rect 12348 15982 12400 15988
rect 12452 15706 12480 16000
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12636 15570 12664 17054
rect 13004 16998 13032 17274
rect 13096 17066 13124 17614
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13188 16590 13216 17070
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13280 16658 13308 17002
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 16250 13216 16526
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13464 15706 13492 16118
rect 13648 16114 13676 16458
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13530 12204 13670
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11992 12406 12112 12434
rect 12084 12209 12112 12406
rect 12070 12200 12126 12209
rect 12070 12135 12126 12144
rect 12164 12164 12216 12170
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11716 9722 11744 10202
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11716 8566 11744 9386
rect 11808 9217 11836 10503
rect 11900 10130 11928 11154
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10130 12020 10950
rect 12084 10577 12112 12135
rect 12164 12106 12216 12112
rect 12176 11898 12204 12106
rect 12268 12102 12296 15370
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 14822 12480 15302
rect 12544 14958 12572 15506
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14346 12480 14758
rect 12544 14618 12572 14894
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 14414 12572 14554
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12440 14340 12492 14346
rect 12360 14300 12440 14328
rect 12360 13190 12388 14300
rect 12440 14282 12492 14288
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12442 12388 12786
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 12360 11914 12388 12378
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12268 11886 12388 11914
rect 12268 11762 12296 11886
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12162 11656 12218 11665
rect 12162 11591 12218 11600
rect 12070 10568 12126 10577
rect 12176 10554 12204 11591
rect 12268 11286 12296 11698
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12360 11218 12388 11494
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12268 10849 12296 11018
rect 12254 10840 12310 10849
rect 12254 10775 12310 10784
rect 12268 10674 12296 10775
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12176 10526 12388 10554
rect 12070 10503 12126 10512
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11900 9110 11928 9522
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8673 11836 8774
rect 11794 8664 11850 8673
rect 11794 8599 11850 8608
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11992 8294 12020 9114
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11716 7698 11744 7958
rect 11808 7886 11836 8230
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11794 7712 11850 7721
rect 11716 7670 11794 7698
rect 11346 7644 11654 7653
rect 11794 7647 11850 7656
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11900 7206 11928 7346
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 10874 6488 10930 6497
rect 10874 6423 10930 6432
rect 10888 6338 10916 6423
rect 10704 6310 10916 6338
rect 10704 5302 10732 6310
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10796 5370 10824 6190
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5710 10916 5743
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10874 5536 10930 5545
rect 10874 5471 10930 5480
rect 10888 5370 10916 5471
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4865 10732 4966
rect 10690 4856 10746 4865
rect 10690 4791 10746 4800
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 4486 10640 4626
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10704 3398 10732 4694
rect 10796 4593 10824 5199
rect 10782 4584 10838 4593
rect 10782 4519 10838 4528
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10796 3210 10824 4519
rect 10888 4486 10916 5306
rect 10980 4826 11008 6802
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11072 4622 11100 6598
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11164 6186 11192 6423
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11152 5636 11204 5642
rect 11152 5578 11204 5584
rect 11164 5148 11192 5578
rect 11256 5574 11284 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11334 5944 11390 5953
rect 11334 5879 11390 5888
rect 11428 5908 11480 5914
rect 11348 5681 11376 5879
rect 11428 5850 11480 5856
rect 11334 5672 11390 5681
rect 11334 5607 11390 5616
rect 11440 5574 11468 5850
rect 11624 5710 11652 6122
rect 11716 6118 11744 6802
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11716 5624 11744 5850
rect 11716 5596 11775 5624
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11747 5234 11775 5596
rect 11704 5228 11775 5234
rect 11756 5188 11775 5228
rect 11704 5170 11756 5176
rect 11336 5160 11388 5166
rect 11164 5120 11336 5148
rect 11336 5102 11388 5108
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 10876 4480 10928 4486
rect 11060 4480 11112 4486
rect 10876 4422 10928 4428
rect 11058 4448 11060 4457
rect 11112 4448 11114 4457
rect 11058 4383 11114 4392
rect 10874 4176 10930 4185
rect 10874 4111 10876 4120
rect 10928 4111 10930 4120
rect 10876 4082 10928 4088
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10704 3182 10824 3210
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10244 2746 10364 2774
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9876 1414 9996 1442
rect 9508 1006 9628 1034
rect 9600 800 9628 1006
rect 9968 800 9996 1414
rect 10336 800 10364 2746
rect 10704 800 10732 3182
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10796 2514 10824 2994
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10980 2446 11008 3946
rect 11058 3768 11114 3777
rect 11058 3703 11114 3712
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11072 800 11100 3703
rect 11164 2582 11192 4966
rect 11808 4826 11836 6598
rect 11900 5030 11928 7142
rect 11992 7002 12020 7278
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11992 6458 12020 6559
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11992 5914 12020 6394
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11256 2310 11284 4762
rect 11624 4690 11652 4762
rect 11900 4690 11928 4966
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11336 4140 11388 4146
rect 11388 4100 11468 4128
rect 11336 4082 11388 4088
rect 11440 4010 11468 4100
rect 11624 4078 11652 4218
rect 11612 4072 11664 4078
rect 11716 4049 11744 4558
rect 11980 4480 12032 4486
rect 11794 4448 11850 4457
rect 12084 4468 12112 10406
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12176 9518 12204 9998
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12176 8906 12204 9454
rect 12360 9450 12388 10526
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 9178 12296 9318
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12176 8430 12204 8842
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12176 8090 12204 8366
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12176 7342 12204 8026
rect 12268 7546 12296 8434
rect 12346 7712 12402 7721
rect 12346 7647 12402 7656
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12254 7440 12310 7449
rect 12254 7375 12310 7384
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12164 7200 12216 7206
rect 12268 7177 12296 7375
rect 12164 7142 12216 7148
rect 12254 7168 12310 7177
rect 12176 6905 12204 7142
rect 12254 7103 12310 7112
rect 12162 6896 12218 6905
rect 12162 6831 12218 6840
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6390 12204 6734
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5710 12204 6122
rect 12254 6080 12310 6089
rect 12254 6015 12310 6024
rect 12268 5710 12296 6015
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12176 5098 12204 5646
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12032 4440 12112 4468
rect 11980 4422 12032 4428
rect 11794 4383 11850 4392
rect 11612 4014 11664 4020
rect 11702 4040 11758 4049
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11520 3936 11572 3942
rect 11518 3904 11520 3913
rect 11572 3904 11574 3913
rect 11518 3839 11574 3848
rect 11624 3738 11652 4014
rect 11702 3975 11758 3984
rect 11702 3904 11758 3913
rect 11702 3839 11758 3848
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 3839
rect 11808 800 11836 4383
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 3777 12020 4218
rect 12176 4146 12204 4694
rect 12256 4276 12308 4282
rect 12360 4264 12388 7647
rect 12452 4554 12480 13806
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12544 11762 12572 12922
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12636 11150 12664 12038
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12728 9058 12756 15574
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15366 12940 15506
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13394 12848 14214
rect 12912 14074 12940 14894
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13004 13394 13032 15302
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13372 13326 13400 14758
rect 13464 14074 13492 15302
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13004 12442 13032 12582
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12806 12336 12862 12345
rect 12806 12271 12862 12280
rect 12820 11830 12848 12271
rect 13004 12238 13032 12378
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12820 10810 12848 11766
rect 13188 11694 13216 12242
rect 13464 11830 13492 12582
rect 13452 11824 13504 11830
rect 13358 11792 13414 11801
rect 13452 11766 13504 11772
rect 13358 11727 13414 11736
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10130 12940 10950
rect 13082 10296 13138 10305
rect 13082 10231 13138 10240
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9178 12848 9522
rect 12990 9480 13046 9489
rect 12990 9415 13046 9424
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12636 9030 12756 9058
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12544 8401 12572 8842
rect 12636 8514 12664 9030
rect 12820 8945 12848 9114
rect 13004 9042 13032 9415
rect 13096 9042 13124 10231
rect 13188 10062 13216 11494
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10266 13308 10950
rect 13372 10606 13400 11727
rect 13452 11688 13504 11694
rect 13556 11642 13584 12650
rect 13504 11636 13584 11642
rect 13452 11630 13584 11636
rect 13464 11614 13584 11630
rect 13464 11218 13492 11614
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10742 13492 11154
rect 13648 10996 13676 16050
rect 13740 13530 13768 19382
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13832 17338 13860 19314
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 18426 14228 18770
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14292 18193 14320 19790
rect 14476 19446 14504 20402
rect 14568 20040 14596 22200
rect 14936 20346 14964 22200
rect 15304 20602 15332 22200
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 14936 20318 15240 20346
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 14648 20052 14700 20058
rect 14568 20012 14648 20040
rect 14648 19994 14700 20000
rect 14752 19854 14780 20198
rect 15120 19854 15148 20198
rect 15212 20058 15240 20318
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15488 19854 15516 20198
rect 15672 20058 15700 22200
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18834 14412 19110
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14278 18184 14334 18193
rect 14278 18119 14334 18128
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14476 17678 14504 18362
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14752 17610 14780 19790
rect 15120 19334 15148 19790
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15028 19306 15148 19334
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14292 16794 14320 17002
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14292 16182 14320 16730
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14476 16114 14504 16594
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14476 15706 14504 16050
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 13924 15473 13952 15574
rect 13910 15464 13966 15473
rect 13910 15399 13966 15408
rect 13924 15162 13952 15399
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14482 13860 14962
rect 14476 14958 14504 15642
rect 14752 15434 14780 16050
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 15570 14872 15982
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 15028 15502 15056 19306
rect 15212 16674 15240 19450
rect 15672 19446 15700 19790
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15660 19168 15712 19174
rect 15658 19136 15660 19145
rect 15712 19136 15714 19145
rect 15658 19071 15714 19080
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15580 18426 15608 18770
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15568 18420 15620 18426
rect 15620 18380 15700 18408
rect 15568 18362 15620 18368
rect 15672 17678 15700 18380
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15120 16646 15240 16674
rect 15120 16028 15148 16646
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15212 16182 15240 16458
rect 15304 16250 15332 17138
rect 15396 17134 15424 17478
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15396 16522 15424 17070
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15488 16046 15516 17614
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17338 15700 17478
rect 15764 17338 15792 18566
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15672 16794 15700 17138
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15764 16250 15792 16730
rect 15856 16250 15884 17138
rect 15948 16538 15976 19654
rect 16040 19514 16068 22200
rect 16408 19514 16436 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19854 16804 20266
rect 16960 20058 16988 20862
rect 17144 20602 17172 22200
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17236 20262 17264 20402
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16488 19304 16540 19310
rect 16960 19281 16988 19314
rect 16488 19246 16540 19252
rect 16946 19272 17002 19281
rect 16500 18737 16528 19246
rect 16946 19207 17002 19216
rect 16486 18728 16542 18737
rect 16486 18663 16542 18672
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 17052 18358 17080 19314
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16658 16068 16934
rect 16132 16658 16160 17002
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 15948 16510 16068 16538
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15476 16040 15528 16046
rect 15120 16000 15240 16028
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15106 15464 15162 15473
rect 14740 15428 14792 15434
rect 15106 15399 15162 15408
rect 14740 15370 14792 15376
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 14016 13870 14044 14554
rect 14292 13870 14320 14894
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14016 13716 14044 13806
rect 14016 13688 14412 13716
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13726 13424 13782 13433
rect 13726 13359 13728 13368
rect 13780 13359 13782 13368
rect 13728 13330 13780 13336
rect 13740 12986 13768 13330
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13740 12753 13768 12922
rect 13726 12744 13782 12753
rect 13726 12679 13782 12688
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11098 13768 12242
rect 13832 11830 13860 13194
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 14384 12434 14412 13688
rect 14292 12406 14412 12434
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13832 11354 13860 11766
rect 14200 11762 14228 12242
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13818 11248 13874 11257
rect 13818 11183 13820 11192
rect 13872 11183 13874 11192
rect 13820 11154 13872 11160
rect 13740 11070 13860 11098
rect 13648 10968 13768 10996
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 10266 13400 10542
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13648 10198 13676 10406
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12806 8936 12862 8945
rect 12806 8871 12862 8880
rect 13004 8634 13032 8978
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12636 8486 12756 8514
rect 12530 8392 12586 8401
rect 12530 8327 12586 8336
rect 12728 7324 12756 8486
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7546 12848 8230
rect 12912 8090 12940 8434
rect 13096 8378 13124 8774
rect 13004 8350 13124 8378
rect 13004 8294 13032 8350
rect 12992 8288 13044 8294
rect 13084 8288 13136 8294
rect 12992 8230 13044 8236
rect 13082 8256 13084 8265
rect 13136 8256 13138 8265
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7342 12940 7890
rect 13004 7750 13032 8230
rect 13082 8191 13138 8200
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7410 13032 7686
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 7336 12860 7342
rect 12728 7296 12808 7324
rect 12808 7278 12860 7284
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12544 7002 12572 7210
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12636 6866 12664 7210
rect 12820 7154 12848 7278
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 13004 7154 13032 7210
rect 13188 7206 13216 9046
rect 12820 7126 13032 7154
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12990 6896 13046 6905
rect 12624 6860 12676 6866
rect 12990 6831 12992 6840
rect 12624 6802 12676 6808
rect 13044 6831 13046 6840
rect 12992 6802 13044 6808
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12544 4826 12572 5170
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12308 4236 12388 4264
rect 12256 4218 12308 4224
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 11978 3768 12034 3777
rect 11978 3703 12034 3712
rect 12084 3466 12112 4014
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12176 3618 12204 3946
rect 12268 3738 12296 4014
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12176 3590 12296 3618
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 2854 12112 3402
rect 12176 3126 12204 3470
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12268 2774 12296 3590
rect 12360 3534 12388 4082
rect 12452 3942 12480 4082
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12348 3528 12400 3534
rect 12544 3482 12572 4422
rect 12348 3470 12400 3476
rect 12452 3454 12572 3482
rect 12452 2836 12480 3454
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3126 12572 3334
rect 12636 3194 12664 6802
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6474 12756 6598
rect 12898 6488 12954 6497
rect 12728 6446 12848 6474
rect 12820 5642 12848 6446
rect 12898 6423 12954 6432
rect 12912 6254 12940 6423
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 13096 6186 13124 6326
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5370 12756 5510
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12820 4706 12848 5578
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12728 4678 12848 4706
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12728 2961 12756 4678
rect 13004 4078 13032 4966
rect 13280 4622 13308 9862
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 8838 13400 9454
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13372 7750 13400 8502
rect 13464 8090 13492 9658
rect 13556 8634 13584 9998
rect 13648 9654 13676 10134
rect 13740 10033 13768 10968
rect 13832 10849 13860 11070
rect 13818 10840 13874 10849
rect 13818 10775 13820 10784
rect 13872 10775 13874 10784
rect 13820 10746 13872 10752
rect 13832 10715 13860 10746
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 13726 10024 13782 10033
rect 13726 9959 13782 9968
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13268 4616 13320 4622
rect 13188 4564 13268 4570
rect 13188 4558 13320 4564
rect 13188 4542 13308 4558
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12820 3194 12848 3470
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12714 2952 12770 2961
rect 12714 2887 12770 2896
rect 12176 2746 12296 2774
rect 12360 2808 12480 2836
rect 12176 800 12204 2746
rect 12360 1902 12388 2808
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12348 1896 12400 1902
rect 12348 1838 12400 1844
rect 12544 800 12572 2246
rect 12820 1170 12848 2518
rect 12912 2446 12940 3878
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13188 2038 13216 4542
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13176 2032 13228 2038
rect 13176 1974 13228 1980
rect 12820 1142 12940 1170
rect 12912 800 12940 1142
rect 13280 800 13308 2790
rect 13372 2650 13400 7686
rect 13556 5914 13584 8366
rect 13648 7800 13676 8774
rect 13740 8498 13768 9959
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13726 8392 13782 8401
rect 13726 8327 13728 8336
rect 13780 8327 13782 8336
rect 13728 8298 13780 8304
rect 13728 7812 13780 7818
rect 13648 7772 13728 7800
rect 13728 7754 13780 7760
rect 13740 7206 13768 7754
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13636 6928 13688 6934
rect 13634 6896 13636 6905
rect 13688 6896 13690 6905
rect 13634 6831 13690 6840
rect 13740 6168 13768 7142
rect 13832 6934 13860 9862
rect 14200 9722 14228 10066
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14292 8634 14320 12406
rect 14568 12238 14596 13806
rect 14660 13802 14688 14350
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13258 14688 13738
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14660 12918 14688 13194
rect 14752 13190 14780 15370
rect 14922 15056 14978 15065
rect 14922 14991 14924 15000
rect 14976 14991 14978 15000
rect 14924 14962 14976 14968
rect 14936 14278 14964 14962
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14660 12306 14688 12854
rect 14752 12850 14780 13126
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14384 10418 14412 10746
rect 14476 10538 14504 11698
rect 14568 11082 14596 12174
rect 14740 11892 14792 11898
rect 14844 11880 14872 12786
rect 14792 11852 14872 11880
rect 14740 11834 14792 11840
rect 14752 11218 14780 11834
rect 15120 11744 15148 15399
rect 15212 14618 15240 16000
rect 15476 15982 15528 15988
rect 15488 15570 15516 15982
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15384 15428 15436 15434
rect 15436 15388 15516 15416
rect 15384 15370 15436 15376
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 13530 15240 13806
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12646 15240 13194
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12306 15240 12582
rect 15292 12368 15344 12374
rect 15290 12336 15292 12345
rect 15344 12336 15346 12345
rect 15200 12300 15252 12306
rect 15290 12271 15346 12280
rect 15200 12242 15252 12248
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14844 11716 15148 11744
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14384 10390 14504 10418
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 9178 14412 9862
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14476 8838 14504 10390
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9042 14596 9522
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14292 8294 14320 8570
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6390 14320 6802
rect 14384 6798 14412 7142
rect 14476 7041 14504 7278
rect 14462 7032 14518 7041
rect 14462 6967 14518 6976
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6458 14412 6598
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 13820 6180 13872 6186
rect 13740 6140 13820 6168
rect 13820 6122 13872 6128
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13648 5302 13676 5714
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13648 4690 13676 5238
rect 13726 4856 13782 4865
rect 13726 4791 13728 4800
rect 13780 4791 13782 4800
rect 13728 4762 13780 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13728 4616 13780 4622
rect 13726 4584 13728 4593
rect 13780 4584 13782 4593
rect 13726 4519 13782 4528
rect 13832 4146 13860 6122
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14292 4758 14320 5510
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13452 3460 13504 3466
rect 13452 3402 13504 3408
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13464 2514 13492 3402
rect 13556 3126 13584 3878
rect 13740 3466 13768 4014
rect 13832 3942 13860 4082
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3720 13860 3878
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13832 3692 13952 3720
rect 13924 3534 13952 3692
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13556 2582 13584 2926
rect 13728 2848 13780 2854
rect 13648 2808 13728 2836
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13648 800 13676 2808
rect 13728 2790 13780 2796
rect 13832 1714 13860 3470
rect 13924 2990 13952 3470
rect 14384 3398 14412 4966
rect 14476 4214 14504 4966
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14568 4078 14596 8298
rect 14660 8294 14688 8910
rect 14648 8288 14700 8294
rect 14648 8230 14700 8236
rect 14646 8120 14702 8129
rect 14752 8090 14780 9862
rect 14844 8090 14872 11716
rect 15304 11354 15332 12038
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10810 14964 10950
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10266 15056 10542
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14936 9654 14964 9930
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 15120 9500 15148 11018
rect 15396 11014 15424 13874
rect 15488 11801 15516 15388
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15474 11792 15530 11801
rect 15580 11762 15608 12582
rect 15474 11727 15530 11736
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15580 11665 15608 11698
rect 15566 11656 15622 11665
rect 15566 11591 15622 11600
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11286 15608 11494
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15672 10826 15700 14214
rect 15764 12374 15792 16186
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15856 14482 15884 14758
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 13938 15976 14350
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13258 15884 13670
rect 15948 13462 15976 13874
rect 16040 13705 16068 16510
rect 16224 16250 16252 17546
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17338 16436 17478
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16776 16561 16804 16934
rect 16762 16552 16818 16561
rect 16762 16487 16764 16496
rect 16816 16487 16818 16496
rect 16764 16458 16816 16464
rect 16304 16448 16356 16454
rect 16776 16427 16804 16458
rect 17040 16448 17092 16454
rect 16304 16390 16356 16396
rect 17040 16390 17092 16396
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16316 16182 16344 16390
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15366 16160 16050
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16026 13696 16082 13705
rect 16026 13631 16082 13640
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15856 12986 15884 13194
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15948 12918 15976 13398
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15752 12368 15804 12374
rect 15804 12328 15884 12356
rect 15752 12310 15804 12316
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11898 15792 12174
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15856 11642 15884 12328
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15396 10798 15700 10826
rect 15764 11614 15884 11642
rect 14936 9472 15148 9500
rect 15200 9512 15252 9518
rect 14646 8055 14702 8064
rect 14740 8084 14792 8090
rect 14660 7585 14688 8055
rect 14740 8026 14792 8032
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14646 7576 14702 7585
rect 14646 7511 14702 7520
rect 14844 7342 14872 8026
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4622 14688 4966
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14660 4185 14688 4422
rect 14752 4298 14780 7210
rect 14844 7002 14872 7278
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6390 14872 6598
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14936 6202 14964 9472
rect 15200 9454 15252 9460
rect 15290 9480 15346 9489
rect 15212 9382 15240 9454
rect 15290 9415 15292 9424
rect 15344 9415 15346 9424
rect 15292 9386 15344 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15028 7818 15056 9318
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15120 8294 15148 8978
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 7342 15056 7754
rect 15304 7546 15332 8366
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 6866 15056 7278
rect 15120 6866 15148 7346
rect 15292 6928 15344 6934
rect 15396 6905 15424 10798
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15672 10130 15700 10678
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15764 9761 15792 11614
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11218 15884 11494
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15948 11014 15976 12038
rect 16040 11898 16068 12038
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16132 11257 16160 15302
rect 16316 15094 16344 15574
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16224 14822 16252 15030
rect 16408 15026 16436 15914
rect 16684 15502 16712 15982
rect 17052 15706 17080 16390
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15162 16988 15438
rect 17144 15162 17172 16050
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 14006 16344 14214
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16408 13802 16436 14962
rect 16592 14482 16620 15098
rect 17236 14906 17264 20198
rect 17512 19514 17540 22200
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 17604 19854 17632 20266
rect 17774 19952 17830 19961
rect 17774 19887 17776 19896
rect 17828 19887 17830 19896
rect 17776 19858 17828 19864
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17604 19446 17632 19790
rect 17880 19514 17908 22200
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 18248 19446 18276 22200
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18432 19922 18460 20334
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18524 19786 18552 20402
rect 18616 20058 18644 22200
rect 18984 20466 19012 22200
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19352 20330 19380 22200
rect 19430 20496 19486 20505
rect 19430 20431 19432 20440
rect 19484 20431 19486 20440
rect 19432 20402 19484 20408
rect 19720 20346 19748 22200
rect 20088 20466 20116 22200
rect 20350 22128 20406 22137
rect 20350 22063 20406 22072
rect 20258 21856 20314 21865
rect 20258 21791 20314 21800
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 19720 20330 19840 20346
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19708 20324 19840 20330
rect 19760 20318 19840 20324
rect 19708 20266 19760 20272
rect 19706 20224 19762 20233
rect 19143 20156 19451 20165
rect 19706 20159 19762 20168
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18616 19854 18644 19994
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18512 19780 18564 19786
rect 18512 19722 18564 19728
rect 18524 19514 18552 19722
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18616 19310 18644 19790
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17144 14878 17264 14906
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 12714 16252 13670
rect 16408 13530 16436 13738
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16868 13462 16896 13874
rect 16960 13530 16988 14214
rect 17052 14074 17080 14282
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 16316 12442 16344 13330
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16960 12918 16988 13330
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12986 17080 13262
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12918 17172 14878
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 12918 17264 14758
rect 17328 14482 17356 14962
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16670 12336 16726 12345
rect 16670 12271 16726 12280
rect 16684 12238 16712 12271
rect 16672 12232 16724 12238
rect 16868 12209 16896 12582
rect 16960 12306 16988 12854
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16854 12200 16910 12209
rect 16672 12174 16724 12180
rect 16776 12170 16854 12186
rect 16764 12164 16854 12170
rect 16816 12158 16854 12164
rect 16854 12135 16910 12144
rect 16764 12106 16816 12112
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16118 11248 16174 11257
rect 16118 11183 16174 11192
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15750 9752 15806 9761
rect 15750 9687 15806 9696
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 8906 15516 9318
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15488 8566 15516 8842
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15672 8294 15700 9454
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 7954 15700 8230
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15856 7750 15884 10950
rect 16132 10266 16160 11086
rect 16224 10810 16252 11698
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16316 11354 16344 11630
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16868 11218 16896 11562
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 17052 11150 17080 12786
rect 17144 11694 17172 12854
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12481 17264 12582
rect 17222 12472 17278 12481
rect 17222 12407 17278 12416
rect 17236 12170 17264 12407
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17132 11688 17184 11694
rect 17130 11656 17132 11665
rect 17184 11656 17186 11665
rect 17130 11591 17186 11600
rect 17328 11558 17356 14282
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17040 11144 17092 11150
rect 16302 11112 16358 11121
rect 17040 11086 17092 11092
rect 16302 11047 16358 11056
rect 16948 11076 17000 11082
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16224 10130 16252 10474
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16316 9722 16344 11047
rect 16948 11018 17000 11024
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10810 16436 10950
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16486 10432 16542 10441
rect 16486 10367 16542 10376
rect 16500 10062 16528 10367
rect 16684 10266 16712 10746
rect 16762 10568 16818 10577
rect 16960 10538 16988 11018
rect 17328 10674 17356 11222
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 16762 10503 16818 10512
rect 16948 10532 17000 10538
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16684 9926 16712 10202
rect 16776 10198 16804 10503
rect 16948 10474 17000 10480
rect 17052 10305 17080 10610
rect 17316 10532 17368 10538
rect 17316 10474 17368 10480
rect 17038 10296 17094 10305
rect 17038 10231 17094 10240
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 17328 10062 17356 10474
rect 16764 10056 16816 10062
rect 17132 10056 17184 10062
rect 16816 10004 17080 10010
rect 16764 9998 17080 10004
rect 17316 10056 17368 10062
rect 17184 10016 17264 10044
rect 17132 9998 17184 10004
rect 16776 9982 17080 9998
rect 16672 9920 16724 9926
rect 16948 9920 17000 9926
rect 16672 9862 16724 9868
rect 16946 9888 16948 9897
rect 17000 9888 17002 9897
rect 16544 9820 16852 9829
rect 16946 9823 17002 9832
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16394 9752 16450 9761
rect 16544 9755 16852 9764
rect 16304 9716 16356 9722
rect 16946 9752 17002 9761
rect 16394 9687 16450 9696
rect 16856 9716 16908 9722
rect 16304 9658 16356 9664
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 8430 15976 8774
rect 16040 8634 16068 9318
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 16132 8090 16160 8434
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16028 7948 16080 7954
rect 16080 7908 16160 7936
rect 16028 7890 16080 7896
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15488 7342 15516 7686
rect 15580 7546 15608 7686
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15292 6870 15344 6876
rect 15382 6896 15438 6905
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15028 6322 15056 6802
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 14936 6174 15056 6202
rect 14830 5400 14886 5409
rect 14830 5335 14886 5344
rect 14844 5234 14872 5335
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4486 14872 5170
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14752 4270 14872 4298
rect 14646 4176 14702 4185
rect 14646 4111 14702 4120
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14476 3534 14504 4014
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3602 14596 3878
rect 14752 3738 14780 4014
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14660 3058 14688 3538
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14292 2514 14320 2926
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 13832 1686 14044 1714
rect 14016 800 14044 1686
rect 14384 800 14412 2858
rect 14844 2774 14872 4270
rect 14936 4214 14964 4966
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14936 3602 14964 4014
rect 15028 3942 15056 6174
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15120 3641 15148 6258
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4282 15240 4422
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15106 3632 15162 3641
rect 14924 3596 14976 3602
rect 15106 3567 15162 3576
rect 14924 3538 14976 3544
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3194 14964 3334
rect 15120 3194 15148 3567
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15120 3058 15148 3130
rect 15304 3058 15332 6870
rect 15382 6831 15438 6840
rect 15396 6338 15424 6831
rect 15488 6798 15516 7278
rect 15580 7002 15608 7346
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15672 6662 15700 7482
rect 15856 7177 15884 7686
rect 15936 7200 15988 7206
rect 15842 7168 15898 7177
rect 15936 7142 15988 7148
rect 15842 7103 15898 7112
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15948 6458 15976 7142
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15396 6310 15700 6338
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15396 5710 15424 6122
rect 15566 5808 15622 5817
rect 15566 5743 15622 5752
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15580 5574 15608 5743
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15396 5166 15424 5510
rect 15580 5370 15608 5510
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15488 4729 15516 5170
rect 15672 4978 15700 6310
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15764 5710 15792 6122
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15750 5264 15806 5273
rect 15750 5199 15806 5208
rect 15580 4950 15700 4978
rect 15474 4720 15530 4729
rect 15474 4655 15530 4664
rect 15382 3904 15438 3913
rect 15382 3839 15438 3848
rect 15396 3534 15424 3839
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15580 3074 15608 4950
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15672 4690 15700 4762
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4214 15700 4626
rect 15764 4622 15792 5199
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15764 4282 15792 4558
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15488 3046 15608 3074
rect 15856 3058 15884 6054
rect 15948 5778 15976 6190
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16040 5302 16068 6598
rect 16132 5896 16160 7908
rect 16224 7546 16252 8230
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 6656 16264 6662
rect 16210 6624 16212 6633
rect 16264 6624 16266 6633
rect 16210 6559 16266 6568
rect 16316 6497 16344 9318
rect 16408 7954 16436 9687
rect 16488 9686 16540 9692
rect 16946 9687 17002 9696
rect 16856 9658 16908 9664
rect 16488 9628 16540 9634
rect 16580 9648 16632 9654
rect 16500 9518 16528 9628
rect 16580 9590 16632 9596
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16592 8838 16620 9590
rect 16672 9376 16724 9382
rect 16670 9344 16672 9353
rect 16764 9376 16816 9382
rect 16724 9344 16726 9353
rect 16764 9318 16816 9324
rect 16670 9279 16726 9288
rect 16776 8974 16804 9318
rect 16764 8968 16816 8974
rect 16868 8945 16896 9658
rect 16764 8910 16816 8916
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8498 16988 9687
rect 17052 9654 17080 9982
rect 17236 9908 17264 10016
rect 17316 9998 17368 10004
rect 17130 9888 17186 9897
rect 17236 9880 17356 9908
rect 17130 9823 17186 9832
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17144 8362 17172 9823
rect 17222 9752 17278 9761
rect 17222 9687 17278 9696
rect 17236 9654 17264 9687
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17236 8430 17264 8774
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 17236 7834 17264 8366
rect 17328 8362 17356 9880
rect 17420 8634 17448 16526
rect 17604 16522 17632 19110
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17880 16250 17908 16662
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15706 17816 15982
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17512 11830 17540 15370
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 15094 17816 15302
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17788 14770 17816 15030
rect 17696 14742 17816 14770
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 13394 17632 14418
rect 17696 13870 17724 14742
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 14074 17816 14214
rect 17880 14074 17908 15846
rect 18248 15502 18276 16118
rect 18340 15502 18368 18294
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18432 15570 18460 15982
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18328 15496 18380 15502
rect 18524 15473 18552 16118
rect 18800 16046 18828 19110
rect 18984 18970 19012 19790
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19076 18970 19104 19246
rect 19352 19174 19380 19314
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18984 18766 19012 18906
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19536 18086 19564 18226
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16794 19564 18022
rect 19628 17542 19656 19858
rect 19720 19446 19748 20159
rect 19812 19854 19840 20318
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19708 19440 19760 19446
rect 19708 19382 19760 19388
rect 19798 19408 19854 19417
rect 19798 19343 19854 19352
rect 19812 18426 19840 19343
rect 19904 19310 19932 20198
rect 20088 19802 20116 20402
rect 20180 20262 20208 20402
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20088 19786 20208 19802
rect 20088 19780 20220 19786
rect 20088 19774 20168 19780
rect 20168 19722 20220 19728
rect 20272 19446 20300 21791
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19628 16674 19656 17478
rect 19352 16646 19656 16674
rect 19352 16574 19380 16646
rect 18892 16546 19380 16574
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18328 15438 18380 15444
rect 18510 15464 18566 15473
rect 18510 15399 18566 15408
rect 18892 15366 18920 16546
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18892 15026 18920 15302
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18236 14816 18288 14822
rect 18156 14776 18236 14804
rect 18156 14346 18184 14776
rect 18236 14758 18288 14764
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17592 13388 17644 13394
rect 17592 13330 17644 13336
rect 17788 13258 17816 13806
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17498 11112 17554 11121
rect 17498 11047 17554 11056
rect 17512 9994 17540 11047
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17052 7806 17264 7834
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16948 7336 17000 7342
rect 17052 7324 17080 7806
rect 17224 7744 17276 7750
rect 17328 7732 17356 7822
rect 17276 7704 17356 7732
rect 17224 7686 17276 7692
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17052 7296 17172 7324
rect 17236 7313 17264 7482
rect 16948 7278 17000 7284
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16302 6488 16358 6497
rect 16544 6491 16852 6500
rect 16960 6458 16988 7278
rect 17144 6798 17172 7296
rect 17222 7304 17278 7313
rect 17222 7239 17278 7248
rect 17328 7206 17356 7704
rect 17512 7528 17540 9522
rect 17420 7500 17540 7528
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17328 6798 17356 7142
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17040 6656 17092 6662
rect 17038 6624 17040 6633
rect 17092 6624 17094 6633
rect 17038 6559 17094 6568
rect 16302 6423 16358 6432
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16394 6216 16450 6225
rect 16394 6151 16450 6160
rect 16132 5868 16344 5896
rect 16118 5808 16174 5817
rect 16118 5743 16174 5752
rect 16132 5710 16160 5743
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 5302 16160 5646
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15948 4826 15976 5102
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16040 4690 16068 5238
rect 16120 5160 16172 5166
rect 16118 5128 16120 5137
rect 16172 5128 16174 5137
rect 16118 5063 16174 5072
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16040 3602 16068 4626
rect 16132 4146 16160 4626
rect 16224 4486 16252 5034
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 3738 16160 4082
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16224 3398 16252 4422
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16224 3126 16252 3334
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16316 3058 16344 5868
rect 16408 5658 16436 6151
rect 17328 6118 17356 6734
rect 17420 6338 17448 7500
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17512 6458 17540 7346
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17420 6322 17540 6338
rect 17420 6316 17552 6322
rect 17420 6310 17500 6316
rect 17500 6258 17552 6264
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16762 5808 16818 5817
rect 16818 5752 16988 5760
rect 16762 5743 16764 5752
rect 16816 5732 16988 5752
rect 16764 5714 16816 5720
rect 16408 5642 16620 5658
rect 16408 5636 16632 5642
rect 16408 5630 16580 5636
rect 16408 5370 16436 5630
rect 16580 5578 16632 5584
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16960 5250 16988 5732
rect 17052 5545 17080 5850
rect 17420 5710 17448 6190
rect 17512 6118 17540 6258
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17408 5704 17460 5710
rect 17406 5672 17408 5681
rect 17460 5672 17462 5681
rect 17512 5642 17540 6054
rect 17406 5607 17462 5616
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17316 5568 17368 5574
rect 17038 5536 17094 5545
rect 17316 5510 17368 5516
rect 17038 5471 17094 5480
rect 17328 5370 17356 5510
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 16684 5222 16988 5250
rect 17040 5228 17092 5234
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16408 4622 16436 5102
rect 16684 4690 16712 5222
rect 17040 5170 17092 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16408 3534 16436 4558
rect 16776 4486 16804 5102
rect 16868 4826 16896 5102
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16856 4684 16908 4690
rect 17052 4672 17080 5170
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 16908 4644 17080 4672
rect 16856 4626 16908 4632
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16856 4004 16908 4010
rect 16960 3992 16988 4422
rect 17052 4146 17080 4644
rect 17144 4282 17172 4762
rect 17222 4720 17278 4729
rect 17222 4655 17278 4664
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17144 4078 17172 4218
rect 17236 4214 17264 4655
rect 17420 4282 17448 4966
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16908 3964 16988 3992
rect 16856 3946 16908 3952
rect 17604 3670 17632 12582
rect 17788 12434 17816 13194
rect 17696 12406 17816 12434
rect 17696 11098 17724 12406
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 11898 17816 12038
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17788 11354 17816 11630
rect 17880 11626 17908 13194
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17972 12646 18000 12922
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18064 12442 18092 12718
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18156 12306 18184 14282
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17972 11626 18000 11766
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17960 11144 18012 11150
rect 17696 11070 17908 11098
rect 17960 11086 18012 11092
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10470 17724 10950
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 9081 17724 10406
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17682 9072 17738 9081
rect 17788 9042 17816 9930
rect 17880 9654 17908 11070
rect 17972 11014 18000 11086
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 18064 10418 18092 11494
rect 18156 11218 18184 12242
rect 18248 11558 18276 12786
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18234 10568 18290 10577
rect 18234 10503 18290 10512
rect 17972 10390 18092 10418
rect 17972 9722 18000 10390
rect 18050 10296 18106 10305
rect 18050 10231 18106 10240
rect 18144 10260 18196 10266
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17682 9007 17738 9016
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17880 8634 17908 9454
rect 18064 9382 18092 10231
rect 18144 10202 18196 10208
rect 18156 9674 18184 10202
rect 18248 10062 18276 10503
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18156 9646 18276 9674
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17972 9081 18000 9114
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17958 8936 18014 8945
rect 17958 8871 18014 8880
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17684 8424 17736 8430
rect 17972 8378 18000 8871
rect 17684 8366 17736 8372
rect 17696 8022 17724 8366
rect 17880 8350 18000 8378
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17788 6798 17816 7278
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17788 6458 17816 6734
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 5710 17816 6190
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17696 3738 17724 4082
rect 17788 4049 17816 5646
rect 17880 4826 17908 8350
rect 17960 7472 18012 7478
rect 17958 7440 17960 7449
rect 18012 7440 18014 7449
rect 17958 7375 18014 7384
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 17972 6730 18000 6831
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 18064 5778 18092 9318
rect 18142 7848 18198 7857
rect 18142 7783 18198 7792
rect 18156 7750 18184 7783
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 5846 18184 7278
rect 18144 5840 18196 5846
rect 18144 5782 18196 5788
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18248 5522 18276 9646
rect 18340 6066 18368 12582
rect 18432 9761 18460 14350
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18524 12186 18552 13670
rect 18708 12646 18736 14282
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 13326 18828 14214
rect 19628 14006 19656 15438
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 13530 18920 13806
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18984 13462 19012 13874
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 18788 13320 18840 13326
rect 19076 13274 19104 13738
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 18788 13262 18840 13268
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18800 12306 18828 13262
rect 18984 13246 19104 13274
rect 18984 13190 19012 13246
rect 18972 13184 19024 13190
rect 19536 13138 19564 13874
rect 19720 13870 19748 14962
rect 19812 14890 19840 18090
rect 19904 17814 19932 19246
rect 20364 18766 20392 22063
rect 20456 20602 20484 22200
rect 20626 21448 20682 21457
rect 20626 21383 20682 21392
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20456 19854 20484 20538
rect 20548 19922 20576 20742
rect 20640 19922 20668 21383
rect 20824 20058 20852 22200
rect 20996 20528 21048 20534
rect 20994 20496 20996 20505
rect 21048 20496 21050 20505
rect 20994 20431 21050 20440
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20456 19378 20484 19790
rect 21192 19446 21220 22200
rect 21454 21040 21510 21049
rect 21454 20975 21510 20984
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20456 18766 20484 19314
rect 20352 18760 20404 18766
rect 20166 18728 20222 18737
rect 20352 18702 20404 18708
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20166 18663 20222 18672
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 18972 13126 19024 13132
rect 18984 12918 19012 13126
rect 19444 13110 19564 13138
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19444 12986 19472 13110
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18524 12158 18736 12186
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11354 18644 12038
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18616 10266 18644 10610
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18708 10146 18736 12158
rect 19076 12102 19104 12582
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 18786 11792 18842 11801
rect 18786 11727 18842 11736
rect 18616 10118 18736 10146
rect 18418 9752 18474 9761
rect 18418 9687 18474 9696
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 8974 18552 9318
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8900 18472 8906
rect 18420 8842 18472 8848
rect 18432 8634 18460 8842
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18524 8498 18552 8910
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18524 7585 18552 7822
rect 18510 7576 18566 7585
rect 18616 7546 18644 10118
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18708 9450 18736 9658
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18708 8974 18736 9386
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8634 18736 8774
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18694 8528 18750 8537
rect 18694 8463 18750 8472
rect 18510 7511 18566 7520
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6866 18644 7142
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18340 6038 18552 6066
rect 18156 5494 18276 5522
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17880 4486 17908 4626
rect 18064 4622 18092 5102
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17774 4040 17830 4049
rect 17774 3975 17830 3984
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16500 3398 16528 3606
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17420 3058 17448 3470
rect 17604 3126 17632 3606
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17788 3058 17816 3975
rect 17880 3602 17908 4422
rect 18050 4176 18106 4185
rect 18050 4111 18106 4120
rect 17958 4040 18014 4049
rect 17958 3975 17960 3984
rect 18012 3975 18014 3984
rect 17960 3946 18012 3952
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17972 3466 18000 3674
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 15844 3052 15896 3058
rect 15488 2774 15516 3046
rect 15844 2994 15896 3000
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 14752 2746 14872 2774
rect 15212 2746 15516 2774
rect 14752 800 14780 2746
rect 15212 2514 15240 2746
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 800 15148 2246
rect 15488 800 15516 2518
rect 15580 2446 15608 2926
rect 16132 2446 16160 2926
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15752 2304 15804 2310
rect 15804 2264 15884 2292
rect 15752 2246 15804 2252
rect 15856 800 15884 2264
rect 16224 800 16252 2858
rect 16684 2650 16712 2994
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1170 16988 2790
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 16868 1142 16988 1170
rect 16592 870 16712 898
rect 16592 800 16620 870
rect 11532 734 11744 762
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16684 762 16712 870
rect 16868 762 16896 1142
rect 17052 898 17080 2518
rect 16960 870 17080 898
rect 16960 800 16988 870
rect 17328 800 17356 2790
rect 17420 2650 17448 2994
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17696 800 17724 2790
rect 17788 2650 17816 2994
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18064 800 18092 4111
rect 18156 3058 18184 5494
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18248 4826 18276 5170
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18248 4078 18276 4762
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4282 18368 4422
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18418 3496 18474 3505
rect 18418 3431 18420 3440
rect 18472 3431 18474 3440
rect 18420 3402 18472 3408
rect 18524 3058 18552 6038
rect 18708 4185 18736 8463
rect 18800 8294 18828 11727
rect 18984 11558 19012 11834
rect 19076 11762 19104 12038
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 19076 11200 19104 11698
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19076 11172 19196 11200
rect 19168 11082 19196 11172
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 18972 11008 19024 11014
rect 18892 10968 18972 10996
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18892 8106 18920 10968
rect 18972 10950 19024 10956
rect 18972 10532 19024 10538
rect 18972 10474 19024 10480
rect 18984 10266 19012 10474
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18984 9722 19012 10202
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18800 8078 18920 8106
rect 18694 4176 18750 4185
rect 18694 4111 18750 4120
rect 18800 3058 18828 8078
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18892 7002 18920 7754
rect 19076 7562 19104 11018
rect 19168 10742 19196 11018
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19168 10538 19196 10678
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19536 9654 19564 12922
rect 19720 12442 19748 13126
rect 19812 12986 19840 13738
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19708 12436 19760 12442
rect 19904 12434 19932 16934
rect 19996 16658 20024 17138
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19996 15094 20024 16050
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19996 13258 20024 14554
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19708 12378 19760 12384
rect 19812 12406 19932 12434
rect 20088 12434 20116 18158
rect 20180 17338 20208 18663
rect 20456 18290 20484 18702
rect 20548 18426 20576 19314
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20456 17882 20484 18226
rect 20732 18034 20760 18838
rect 21284 18766 21312 20198
rect 21362 19816 21418 19825
rect 21362 19751 21418 19760
rect 21376 18970 21404 19751
rect 21468 19446 21496 20975
rect 21560 20398 21588 22200
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 21454 19000 21510 19009
rect 21364 18964 21416 18970
rect 21454 18935 21510 18944
rect 21364 18906 21416 18912
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20640 18006 20760 18034
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 13190 20208 16458
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20088 12406 20300 12434
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19628 10810 19656 11698
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19628 10130 19656 10746
rect 19720 10606 19748 11018
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 9722 19748 9862
rect 19708 9716 19760 9722
rect 19708 9658 19760 9664
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8378 19288 8910
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19260 8350 19472 8378
rect 19444 8294 19472 8350
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19536 8090 19564 8434
rect 19628 8294 19656 8325
rect 19616 8288 19668 8294
rect 19720 8242 19748 8434
rect 19668 8236 19748 8242
rect 19616 8230 19748 8236
rect 19628 8214 19748 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 18984 7534 19196 7562
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 5574 18920 6598
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 5302 18920 5510
rect 18984 5302 19012 7534
rect 19168 7410 19196 7534
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19076 7002 19104 7346
rect 19352 7324 19380 7686
rect 19444 7546 19472 7822
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19536 7478 19564 8026
rect 19628 7750 19656 8214
rect 19812 7993 19840 12406
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19904 8974 19932 11290
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19904 8362 19932 8910
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19798 7984 19854 7993
rect 19798 7919 19854 7928
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19904 7528 19932 8298
rect 19812 7500 19932 7528
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19352 7296 19564 7324
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6633 19472 6734
rect 19536 6662 19564 7296
rect 19524 6656 19576 6662
rect 19430 6624 19486 6633
rect 19524 6598 19576 6604
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19430 6559 19486 6568
rect 19720 6254 19748 6598
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19524 5636 19576 5642
rect 19524 5578 19576 5584
rect 19536 5370 19564 5578
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4486 18920 4966
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18984 4026 19012 5238
rect 19536 5166 19564 5306
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 4282 19288 4422
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19524 4072 19576 4078
rect 18984 3998 19104 4026
rect 19524 4014 19576 4020
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18984 3670 19012 3878
rect 19076 3738 19104 3998
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 19076 3534 19104 3674
rect 19536 3602 19564 4014
rect 19628 4010 19656 5170
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19720 4486 19748 4762
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 19076 3097 19104 3470
rect 19720 3398 19748 4422
rect 19812 4146 19840 7500
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 6458 19932 7346
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19904 6186 19932 6258
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19904 5914 19932 6122
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19904 4214 19932 5102
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19062 3088 19118 3097
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18788 3052 18840 3058
rect 19062 3023 19118 3032
rect 18788 2994 18840 3000
rect 18156 2650 18184 2994
rect 18524 2650 18552 2994
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 18432 800 18460 2314
rect 18800 800 18828 2858
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18984 1442 19012 2790
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 18984 1414 19196 1442
rect 19168 800 19196 1414
rect 19536 800 19564 2858
rect 19996 2774 20024 12242
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 10810 20208 12174
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 10266 20116 10610
rect 20272 10418 20300 12406
rect 20180 10390 20300 10418
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20088 8362 20116 8570
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20088 6934 20116 7278
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20088 4758 20116 5510
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20088 3942 20116 4218
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19904 2746 20024 2774
rect 19904 800 19932 2746
rect 20088 2417 20116 3878
rect 20180 2774 20208 10390
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 8090 20300 9522
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20364 7562 20392 17478
rect 20640 17082 20668 18006
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20548 17054 20668 17082
rect 20548 13433 20576 17054
rect 20824 16998 20852 17138
rect 20812 16992 20864 16998
rect 20626 16960 20682 16969
rect 20812 16934 20864 16940
rect 20626 16895 20682 16904
rect 20640 16250 20668 16895
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20534 13424 20590 13433
rect 20534 13359 20590 13368
rect 20548 13326 20576 13359
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 12986 20484 13126
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20548 12918 20576 13262
rect 20640 13002 20668 15982
rect 20916 14618 20944 16050
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20640 12974 20760 13002
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20626 12880 20682 12889
rect 20444 12844 20496 12850
rect 20626 12815 20682 12824
rect 20444 12786 20496 12792
rect 20456 12374 20484 12786
rect 20534 12472 20590 12481
rect 20640 12442 20668 12815
rect 20534 12407 20590 12416
rect 20628 12436 20680 12442
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20456 11082 20484 11494
rect 20548 11354 20576 12407
rect 20628 12378 20680 12384
rect 20732 12306 20760 12974
rect 20916 12646 20944 13262
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20456 9518 20484 10134
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 9042 20484 9454
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20548 8634 20576 9862
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20640 9489 20668 9522
rect 20626 9480 20682 9489
rect 20626 9415 20682 9424
rect 20732 9178 20760 10610
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20824 10266 20852 10542
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9722 20852 9930
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 9110 20852 9454
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20824 8430 20852 9046
rect 20812 8424 20864 8430
rect 20732 8384 20812 8412
rect 20442 7984 20498 7993
rect 20732 7954 20760 8384
rect 20812 8366 20864 8372
rect 20442 7919 20444 7928
rect 20496 7919 20498 7928
rect 20720 7948 20772 7954
rect 20444 7890 20496 7896
rect 20720 7890 20772 7896
rect 20456 7698 20484 7890
rect 20456 7670 20576 7698
rect 20364 7534 20484 7562
rect 20548 7546 20576 7670
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20364 6390 20392 6802
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 5914 20300 6190
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20180 2746 20300 2774
rect 20074 2408 20130 2417
rect 20074 2343 20130 2352
rect 20272 800 20300 2746
rect 20364 1465 20392 3946
rect 20456 2774 20484 7534
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20732 7342 20760 7890
rect 20916 7886 20944 9862
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7410 20944 7686
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20548 6390 20576 6734
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20824 5817 20852 6258
rect 20810 5808 20866 5817
rect 20810 5743 20866 5752
rect 20824 5370 20852 5743
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20916 5302 20944 6734
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 20456 2746 20668 2774
rect 20350 1456 20406 1465
rect 20350 1391 20406 1400
rect 20640 800 20668 2746
rect 21008 800 21036 18634
rect 21468 18426 21496 18935
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21362 18184 21418 18193
rect 21362 18119 21418 18128
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 21100 17338 21128 17711
rect 21376 17338 21404 18119
rect 21560 17882 21588 19994
rect 21652 18358 21680 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22296 18630 22324 22200
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21086 17232 21142 17241
rect 21086 17167 21142 17176
rect 21100 16794 21128 17167
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21086 16552 21142 16561
rect 21086 16487 21142 16496
rect 21100 16250 21128 16487
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21192 16114 21220 16390
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21376 16153 21404 16186
rect 21362 16144 21418 16153
rect 21180 16108 21232 16114
rect 21362 16079 21418 16088
rect 21180 16050 21232 16056
rect 21362 15736 21418 15745
rect 21362 15671 21364 15680
rect 21416 15671 21418 15680
rect 21364 15642 21416 15648
rect 21086 15464 21142 15473
rect 21086 15399 21142 15408
rect 21100 15366 21128 15399
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21362 14920 21418 14929
rect 21362 14855 21418 14864
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21088 14544 21140 14550
rect 21086 14512 21088 14521
rect 21140 14512 21142 14521
rect 21086 14447 21142 14456
rect 21192 14414 21220 14758
rect 21376 14618 21404 14855
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13977 21128 14010
rect 21086 13968 21142 13977
rect 21086 13903 21142 13912
rect 21086 13288 21142 13297
rect 21086 13223 21142 13232
rect 21100 13190 21128 13223
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21192 11830 21220 14350
rect 21454 13696 21510 13705
rect 21454 13631 21510 13640
rect 21468 13530 21496 13631
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12918 21312 13262
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 21560 12434 21588 17546
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 21468 12406 21588 12434
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21376 11762 21404 12038
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21100 7818 21128 11086
rect 21192 9654 21220 11562
rect 21284 11082 21312 11562
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21284 10810 21312 11018
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21192 7546 21220 9454
rect 21284 7886 21312 9862
rect 21376 8974 21404 11494
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21376 7954 21404 8502
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21100 6322 21128 7346
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21100 5574 21128 5850
rect 21284 5574 21312 7686
rect 21376 7274 21404 7754
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21376 6118 21404 7210
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5642 21404 6054
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21100 4468 21128 5510
rect 21180 4480 21232 4486
rect 21100 4440 21180 4468
rect 21180 4422 21232 4428
rect 21192 2689 21220 4422
rect 21468 2774 21496 12406
rect 21546 12200 21602 12209
rect 21546 12135 21602 12144
rect 21560 6662 21588 12135
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21652 11082 21680 11630
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21652 10538 21680 11018
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21640 10532 21692 10538
rect 21640 10474 21692 10480
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21652 8362 21680 9862
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21640 8356 21692 8362
rect 21640 8298 21692 8304
rect 21652 7750 21680 8298
rect 21744 7818 21772 8570
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21560 5030 21588 6258
rect 22112 5914 22140 11698
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22204 5794 22232 11018
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22112 5766 22232 5794
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21560 4486 21588 4966
rect 21652 4554 21680 5510
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 3505 21588 4422
rect 21546 3496 21602 3505
rect 21546 3431 21602 3440
rect 21376 2746 21496 2774
rect 21178 2680 21234 2689
rect 21178 2615 21234 2624
rect 21376 800 21404 2746
rect 21652 1873 21680 4490
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 22112 4282 22140 5766
rect 22296 5710 22324 8366
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21638 1864 21694 1873
rect 21638 1799 21694 1808
rect 22006 1048 22062 1057
rect 22204 1034 22232 5578
rect 22062 1006 22232 1034
rect 22006 983 22062 992
rect 16684 734 16896 762
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 22006 640 22062 649
rect 22296 626 22324 5646
rect 22388 4622 22416 12582
rect 22480 6390 22508 16934
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22572 4826 22600 16458
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22062 598 22324 626
rect 22006 575 22062 584
<< via2 >>
rect 2318 19760 2374 19816
rect 1950 19352 2006 19408
rect 1582 18964 1638 19000
rect 1582 18944 1584 18964
rect 1584 18944 1636 18964
rect 1636 18944 1638 18964
rect 1950 18536 2006 18592
rect 1766 18128 1822 18184
rect 1766 17720 1822 17776
rect 1950 17620 1952 17640
rect 1952 17620 2004 17640
rect 2004 17620 2006 17640
rect 1950 17584 2006 17620
rect 1858 17312 1914 17368
rect 1858 16496 1914 16552
rect 1950 16088 2006 16144
rect 1766 15272 1822 15328
rect 3698 22072 3754 22128
rect 2778 18944 2834 19000
rect 2226 17176 2282 17232
rect 3146 18672 3202 18728
rect 2778 16904 2834 16960
rect 2318 15700 2374 15736
rect 2318 15680 2320 15700
rect 2320 15680 2372 15700
rect 2372 15680 2374 15700
rect 2594 15544 2650 15600
rect 2134 15000 2190 15056
rect 1582 14492 1584 14512
rect 1584 14492 1636 14512
rect 1636 14492 1638 14512
rect 1582 14456 1638 14492
rect 1582 13640 1638 13696
rect 1858 13232 1914 13288
rect 1582 12436 1638 12472
rect 1582 12416 1584 12436
rect 1584 12416 1636 12436
rect 1636 12416 1638 12436
rect 2502 14048 2558 14104
rect 2410 12824 2466 12880
rect 2870 14864 2926 14920
rect 2686 12688 2742 12744
rect 4066 21800 4122 21856
rect 3974 21392 4030 21448
rect 3882 21004 3938 21040
rect 3882 20984 3884 21004
rect 3884 20984 3936 21004
rect 3936 20984 3938 21004
rect 3974 20440 4030 20496
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3974 19352 4030 19408
rect 3422 17992 3478 18048
rect 4158 18844 4160 18864
rect 4160 18844 4212 18864
rect 4212 18844 4214 18864
rect 4158 18808 4214 18844
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 4526 18672 4582 18728
rect 4802 18964 4858 19000
rect 4802 18944 4804 18964
rect 4804 18944 4856 18964
rect 4856 18944 4858 18964
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3422 14340 3478 14376
rect 3422 14320 3424 14340
rect 3424 14320 3476 14340
rect 3476 14320 3478 14340
rect 4066 14864 4122 14920
rect 3974 14220 3976 14240
rect 3976 14220 4028 14240
rect 4028 14220 4030 14240
rect 3974 14184 4030 14220
rect 3238 13912 3294 13968
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 1398 12008 1454 12064
rect 1214 7112 1270 7168
rect 1490 2896 1546 2952
rect 1766 3440 1822 3496
rect 4250 13368 4306 13424
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 2318 7384 2374 7440
rect 2962 8744 3018 8800
rect 2870 8084 2926 8120
rect 2870 8064 2872 8084
rect 2872 8064 2924 8084
rect 2924 8064 2926 8084
rect 3054 6604 3056 6624
rect 3056 6604 3108 6624
rect 3108 6604 3110 6624
rect 3054 6568 3110 6604
rect 1858 3032 1914 3088
rect 1582 2624 1638 2680
rect 3882 11600 3938 11656
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3974 11192 4030 11248
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 4066 9968 4122 10024
rect 4066 9560 4122 9616
rect 3974 9016 4030 9072
rect 3882 8336 3938 8392
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3054 3848 3110 3904
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3790 6860 3846 6896
rect 3790 6840 3792 6860
rect 3792 6840 3844 6860
rect 3844 6840 3846 6860
rect 3790 6704 3846 6760
rect 3606 6432 3662 6488
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3882 5208 3938 5264
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 5078 20576 5134 20632
rect 4986 16108 5042 16144
rect 4986 16088 4988 16108
rect 4988 16088 5040 16108
rect 5040 16088 5042 16108
rect 4986 15272 5042 15328
rect 4894 12280 4950 12336
rect 4066 7928 4122 7984
rect 4066 6296 4122 6352
rect 4066 4664 4122 4720
rect 2778 2216 2834 2272
rect 2686 1808 2742 1864
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 1400 3478 1456
rect 5630 19796 5632 19816
rect 5632 19796 5684 19816
rect 5684 19796 5686 19816
rect 5630 19760 5686 19796
rect 5906 20324 5962 20360
rect 5906 20304 5908 20324
rect 5908 20304 5960 20324
rect 5960 20304 5962 20324
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5170 16904 5226 16960
rect 5078 12824 5134 12880
rect 4894 9324 4896 9344
rect 4896 9324 4948 9344
rect 4948 9324 4950 9344
rect 4894 9288 4950 9324
rect 4986 9036 5042 9072
rect 4986 9016 4988 9036
rect 4988 9016 5040 9036
rect 5040 9016 5042 9036
rect 4986 7420 4988 7440
rect 4988 7420 5040 7440
rect 5040 7420 5042 7440
rect 4986 7384 5042 7420
rect 4342 992 4398 1048
rect 5078 6840 5134 6896
rect 5446 16904 5502 16960
rect 5538 15308 5540 15328
rect 5540 15308 5592 15328
rect 5592 15308 5594 15328
rect 5538 15272 5594 15308
rect 5722 18828 5778 18864
rect 5722 18808 5724 18828
rect 5724 18808 5776 18828
rect 5776 18808 5778 18828
rect 5722 18672 5778 18728
rect 6458 18944 6514 19000
rect 6090 18672 6146 18728
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6090 18264 6146 18320
rect 5814 16904 5870 16960
rect 5630 12824 5686 12880
rect 5262 9016 5318 9072
rect 5354 8628 5410 8664
rect 5354 8608 5356 8628
rect 5356 8608 5408 8628
rect 5408 8608 5410 8628
rect 5630 12008 5686 12064
rect 6734 18808 6790 18864
rect 6826 18672 6882 18728
rect 6826 18264 6882 18320
rect 6642 18128 6698 18184
rect 6642 17992 6698 18048
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6366 15544 6422 15600
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 7470 19760 7526 19816
rect 6918 17992 6974 18048
rect 6734 17584 6790 17640
rect 6918 17040 6974 17096
rect 7010 16652 7066 16688
rect 7010 16632 7012 16652
rect 7012 16632 7064 16652
rect 7064 16632 7066 16652
rect 6826 15136 6882 15192
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6826 13232 6882 13288
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5722 9424 5778 9480
rect 6642 10104 6698 10160
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6550 9696 6606 9752
rect 5906 9288 5962 9344
rect 5446 7792 5502 7848
rect 5078 6568 5134 6624
rect 5354 6432 5410 6488
rect 5078 5344 5134 5400
rect 4894 5108 4896 5128
rect 4896 5108 4948 5128
rect 4948 5108 4950 5128
rect 4894 5072 4950 5108
rect 5078 4528 5134 4584
rect 5722 7656 5778 7712
rect 5722 7384 5778 7440
rect 6550 9152 6606 9208
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6090 8372 6092 8392
rect 6092 8372 6144 8392
rect 6144 8372 6146 8392
rect 6090 8336 6146 8372
rect 7010 11056 7066 11112
rect 7010 9580 7066 9616
rect 7010 9560 7012 9580
rect 7012 9560 7064 9580
rect 7064 9560 7066 9580
rect 6826 8336 6882 8392
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5814 7248 5870 7304
rect 5538 3440 5594 3496
rect 6274 6704 6330 6760
rect 6458 6704 6514 6760
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6642 6840 6698 6896
rect 6642 6568 6698 6624
rect 6642 6432 6698 6488
rect 6182 6180 6238 6216
rect 6182 6160 6184 6180
rect 6184 6160 6236 6180
rect 6236 6160 6238 6180
rect 5998 5772 6054 5808
rect 5998 5752 6000 5772
rect 6000 5752 6052 5772
rect 6052 5752 6054 5772
rect 7010 7520 7066 7576
rect 6826 5888 6882 5944
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6642 5344 6698 5400
rect 6642 5072 6698 5128
rect 6550 4936 6606 4992
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6090 3440 6146 3496
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6918 2932 6920 2952
rect 6920 2932 6972 2952
rect 6972 2932 6974 2952
rect 6918 2896 6974 2932
rect 6642 2216 6698 2272
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7286 16360 7342 16416
rect 7286 15952 7342 16008
rect 7838 18672 7894 18728
rect 7654 16940 7656 16960
rect 7656 16940 7708 16960
rect 7708 16940 7710 16960
rect 7654 16904 7710 16940
rect 8114 17176 8170 17232
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 9034 19352 9090 19408
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8574 17584 8630 17640
rect 7562 14592 7618 14648
rect 7378 13096 7434 13152
rect 7746 13388 7802 13424
rect 7746 13368 7748 13388
rect 7748 13368 7800 13388
rect 7800 13368 7802 13388
rect 7930 12824 7986 12880
rect 7746 11636 7748 11656
rect 7748 11636 7800 11656
rect 7800 11636 7802 11656
rect 7746 11600 7802 11636
rect 7194 7384 7250 7440
rect 7562 7520 7618 7576
rect 7746 9560 7802 9616
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 9126 17756 9128 17776
rect 9128 17756 9180 17776
rect 9180 17756 9182 17776
rect 9126 17720 9182 17756
rect 9310 18672 9366 18728
rect 9402 18128 9458 18184
rect 8114 14184 8170 14240
rect 8022 8880 8078 8936
rect 7746 6568 7802 6624
rect 7378 3032 7434 3088
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8666 14864 8722 14920
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8482 14184 8538 14240
rect 8390 13368 8446 13424
rect 8298 11872 8354 11928
rect 8206 11056 8262 11112
rect 8206 10140 8208 10160
rect 8208 10140 8260 10160
rect 8260 10140 8262 10160
rect 8206 10104 8262 10140
rect 8942 14048 8998 14104
rect 9218 14048 9274 14104
rect 9218 13676 9220 13696
rect 9220 13676 9272 13696
rect 9272 13676 9274 13696
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9218 13640 9274 13676
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8574 11756 8630 11792
rect 8574 11736 8576 11756
rect 8576 11736 8628 11756
rect 8628 11736 8630 11756
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8206 8608 8262 8664
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8666 9832 8722 9888
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9586 16496 9642 16552
rect 9586 15000 9642 15056
rect 9494 13912 9550 13968
rect 9494 13640 9550 13696
rect 9402 11872 9458 11928
rect 9218 10260 9274 10296
rect 9218 10240 9220 10260
rect 9220 10240 9272 10260
rect 9272 10240 9274 10260
rect 8666 8608 8722 8664
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8390 6568 8446 6624
rect 8390 5752 8446 5808
rect 8206 5072 8262 5128
rect 8114 3984 8170 4040
rect 8022 2932 8024 2952
rect 8024 2932 8076 2952
rect 8076 2932 8078 2952
rect 8022 2896 8078 2932
rect 3882 584 3938 640
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8758 6704 8814 6760
rect 8942 6704 8998 6760
rect 8942 6568 8998 6624
rect 9126 6452 9182 6488
rect 9126 6432 9128 6452
rect 9128 6432 9180 6452
rect 9180 6432 9182 6452
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9126 5908 9182 5944
rect 9126 5888 9128 5908
rect 9128 5888 9180 5908
rect 9180 5888 9182 5908
rect 9310 9152 9366 9208
rect 9218 5616 9274 5672
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8850 4120 8906 4176
rect 9034 3984 9090 4040
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9770 13776 9826 13832
rect 9862 13368 9918 13424
rect 10046 18672 10102 18728
rect 10598 19896 10654 19952
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10874 18264 10930 18320
rect 10322 17992 10378 18048
rect 10046 14048 10102 14104
rect 9862 12688 9918 12744
rect 9402 7948 9458 7984
rect 9402 7928 9404 7948
rect 9404 7928 9456 7948
rect 9456 7928 9458 7948
rect 9862 7792 9918 7848
rect 9678 6296 9734 6352
rect 9678 5616 9734 5672
rect 9862 4664 9918 4720
rect 9862 4528 9918 4584
rect 8850 2488 8906 2544
rect 9678 3848 9734 3904
rect 9862 3576 9918 3632
rect 10138 9288 10194 9344
rect 10046 8744 10102 8800
rect 10322 13776 10378 13832
rect 10322 10684 10324 10704
rect 10324 10684 10376 10704
rect 10376 10684 10378 10704
rect 10322 10648 10378 10684
rect 12806 19116 12808 19136
rect 12808 19116 12860 19136
rect 12860 19116 12862 19136
rect 12806 19080 12862 19116
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11610 18028 11612 18048
rect 11612 18028 11664 18048
rect 11664 18028 11666 18048
rect 11610 17992 11666 18028
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 12254 18420 12310 18456
rect 12254 18400 12256 18420
rect 12256 18400 12308 18420
rect 12308 18400 12310 18420
rect 12162 18284 12218 18320
rect 12162 18264 12164 18284
rect 12164 18264 12216 18284
rect 12216 18264 12218 18284
rect 12070 18128 12126 18184
rect 11334 16496 11390 16552
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11058 14900 11060 14920
rect 11060 14900 11112 14920
rect 11112 14900 11114 14920
rect 11058 14864 11114 14900
rect 10966 13912 11022 13968
rect 10874 13812 10876 13832
rect 10876 13812 10928 13832
rect 10928 13812 10930 13832
rect 10874 13776 10930 13812
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11518 13776 11574 13832
rect 10598 12416 10654 12472
rect 10690 12280 10746 12336
rect 10414 10512 10470 10568
rect 10506 9832 10562 9888
rect 11978 16496 12034 16552
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10874 10648 10930 10704
rect 10690 9696 10746 9752
rect 10322 9560 10378 9616
rect 10230 7792 10286 7848
rect 10138 7656 10194 7712
rect 10414 8200 10470 8256
rect 10138 6024 10194 6080
rect 10506 8064 10562 8120
rect 10322 4392 10378 4448
rect 10322 3576 10378 3632
rect 10966 8064 11022 8120
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13634 19116 13636 19136
rect 13636 19116 13688 19136
rect 13688 19116 13690 19136
rect 13634 19080 13690 19116
rect 12990 18264 13046 18320
rect 12714 17176 12770 17232
rect 12070 12144 12126 12200
rect 11794 10512 11850 10568
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 12162 11600 12218 11656
rect 12070 10512 12126 10568
rect 12254 10784 12310 10840
rect 11794 9152 11850 9208
rect 11794 8608 11850 8664
rect 11794 7656 11850 7712
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10874 6432 10930 6488
rect 10874 5752 10930 5808
rect 10874 5480 10930 5536
rect 10782 5208 10838 5264
rect 10690 4800 10746 4856
rect 10782 4528 10838 4584
rect 11150 6432 11206 6488
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11334 5888 11390 5944
rect 11334 5616 11390 5672
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11058 4428 11060 4448
rect 11060 4428 11112 4448
rect 11112 4428 11114 4448
rect 11058 4392 11114 4428
rect 10874 4140 10930 4176
rect 10874 4120 10876 4140
rect 10876 4120 10928 4140
rect 10928 4120 10930 4140
rect 11058 3712 11114 3768
rect 11978 6568 12034 6624
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11794 4392 11850 4448
rect 12346 7656 12402 7712
rect 12254 7384 12310 7440
rect 12254 7112 12310 7168
rect 12162 6840 12218 6896
rect 12254 6024 12310 6080
rect 11518 3884 11520 3904
rect 11520 3884 11572 3904
rect 11572 3884 11574 3904
rect 11518 3848 11574 3884
rect 11702 3984 11758 4040
rect 11702 3848 11758 3904
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12806 12280 12862 12336
rect 13358 11736 13414 11792
rect 13082 10240 13138 10296
rect 12990 9424 13046 9480
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 14278 18128 14334 18184
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13910 15408 13966 15464
rect 15658 19116 15660 19136
rect 15660 19116 15712 19136
rect 15712 19116 15714 19136
rect 15658 19080 15714 19116
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16946 19216 17002 19272
rect 16486 18672 16542 18728
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 15106 15408 15162 15464
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13726 13388 13782 13424
rect 13726 13368 13728 13388
rect 13728 13368 13780 13388
rect 13780 13368 13782 13388
rect 13726 12688 13782 12744
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13818 11212 13874 11248
rect 13818 11192 13820 11212
rect 13820 11192 13872 11212
rect 13872 11192 13874 11212
rect 12806 8880 12862 8936
rect 12530 8336 12586 8392
rect 13082 8236 13084 8256
rect 13084 8236 13136 8256
rect 13136 8236 13138 8256
rect 13082 8200 13138 8236
rect 12990 6860 13046 6896
rect 12990 6840 12992 6860
rect 12992 6840 13044 6860
rect 13044 6840 13046 6860
rect 11978 3712 12034 3768
rect 12898 6432 12954 6488
rect 13818 10804 13874 10840
rect 13818 10784 13820 10804
rect 13820 10784 13872 10804
rect 13872 10784 13874 10804
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13726 9968 13782 10024
rect 12714 2896 12770 2952
rect 13726 8356 13782 8392
rect 13726 8336 13728 8356
rect 13728 8336 13780 8356
rect 13780 8336 13782 8356
rect 13634 6876 13636 6896
rect 13636 6876 13688 6896
rect 13688 6876 13690 6896
rect 13634 6840 13690 6876
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14922 15020 14978 15056
rect 14922 15000 14924 15020
rect 14924 15000 14976 15020
rect 14976 15000 14978 15020
rect 15290 12316 15292 12336
rect 15292 12316 15344 12336
rect 15344 12316 15346 12336
rect 15290 12280 15346 12316
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 14462 6976 14518 7032
rect 13726 4820 13782 4856
rect 13726 4800 13728 4820
rect 13728 4800 13780 4820
rect 13780 4800 13782 4820
rect 13726 4564 13728 4584
rect 13728 4564 13780 4584
rect 13780 4564 13782 4584
rect 13726 4528 13782 4564
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14646 8064 14702 8120
rect 15474 11736 15530 11792
rect 15566 11600 15622 11656
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16762 16516 16818 16552
rect 16762 16496 16764 16516
rect 16764 16496 16816 16516
rect 16816 16496 16818 16516
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16026 13640 16082 13696
rect 14646 7520 14702 7576
rect 15290 9444 15346 9480
rect 15290 9424 15292 9444
rect 15292 9424 15344 9444
rect 15344 9424 15346 9444
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 17774 19916 17830 19952
rect 17774 19896 17776 19916
rect 17776 19896 17828 19916
rect 17828 19896 17830 19916
rect 19430 20460 19486 20496
rect 19430 20440 19432 20460
rect 19432 20440 19484 20460
rect 19484 20440 19486 20460
rect 20350 22072 20406 22128
rect 20258 21800 20314 21856
rect 19706 20168 19762 20224
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16670 12280 16726 12336
rect 16854 12144 16910 12200
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16118 11192 16174 11248
rect 15750 9696 15806 9752
rect 17222 12416 17278 12472
rect 17130 11636 17132 11656
rect 17132 11636 17184 11656
rect 17184 11636 17186 11656
rect 17130 11600 17186 11636
rect 16302 11056 16358 11112
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16486 10376 16542 10432
rect 16762 10512 16818 10568
rect 17038 10240 17094 10296
rect 16946 9868 16948 9888
rect 16948 9868 17000 9888
rect 17000 9868 17002 9888
rect 16946 9832 17002 9868
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16394 9696 16450 9752
rect 14830 5344 14886 5400
rect 14646 4120 14702 4176
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15106 3576 15162 3632
rect 15382 6840 15438 6896
rect 15842 7112 15898 7168
rect 15566 5752 15622 5808
rect 15750 5208 15806 5264
rect 15474 4664 15530 4720
rect 15382 3848 15438 3904
rect 16210 6604 16212 6624
rect 16212 6604 16264 6624
rect 16264 6604 16266 6624
rect 16210 6568 16266 6604
rect 16946 9696 17002 9752
rect 16670 9324 16672 9344
rect 16672 9324 16724 9344
rect 16724 9324 16726 9344
rect 16670 9288 16726 9324
rect 16854 8880 16910 8936
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 17130 9832 17186 9888
rect 17222 9696 17278 9752
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19798 19352 19854 19408
rect 18510 15408 18566 15464
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 17498 11056 17554 11112
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16302 6432 16358 6488
rect 17222 7248 17278 7304
rect 17038 6604 17040 6624
rect 17040 6604 17092 6624
rect 17092 6604 17094 6624
rect 17038 6568 17094 6604
rect 16394 6160 16450 6216
rect 16118 5752 16174 5808
rect 16118 5108 16120 5128
rect 16120 5108 16172 5128
rect 16172 5108 16174 5128
rect 16118 5072 16174 5108
rect 16762 5772 16818 5808
rect 16762 5752 16764 5772
rect 16764 5752 16816 5772
rect 16816 5752 16818 5772
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17406 5652 17408 5672
rect 17408 5652 17460 5672
rect 17460 5652 17462 5672
rect 17406 5616 17462 5652
rect 17038 5480 17094 5536
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17222 4664 17278 4720
rect 17682 9016 17738 9072
rect 18234 10512 18290 10568
rect 18050 10240 18106 10296
rect 17958 9016 18014 9072
rect 17958 8880 18014 8936
rect 17958 7420 17960 7440
rect 17960 7420 18012 7440
rect 18012 7420 18014 7440
rect 17958 7384 18014 7420
rect 17958 6840 18014 6896
rect 18142 7792 18198 7848
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 20626 21392 20682 21448
rect 20994 20476 20996 20496
rect 20996 20476 21048 20496
rect 21048 20476 21050 20496
rect 20994 20440 21050 20476
rect 21454 20984 21510 21040
rect 20166 18672 20222 18728
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18786 11736 18842 11792
rect 18418 9696 18474 9752
rect 18510 7520 18566 7576
rect 18694 8472 18750 8528
rect 17774 3984 17830 4040
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 18050 4120 18106 4176
rect 17958 4004 18014 4040
rect 17958 3984 17960 4004
rect 17960 3984 18012 4004
rect 18012 3984 18014 4004
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 18418 3460 18474 3496
rect 18418 3440 18420 3460
rect 18420 3440 18472 3460
rect 18472 3440 18474 3460
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 18694 4120 18750 4176
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 21362 19760 21418 19816
rect 21454 18944 21510 19000
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19798 7928 19854 7984
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19430 6568 19486 6624
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19062 3032 19118 3088
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20626 16904 20682 16960
rect 20534 13368 20590 13424
rect 20626 12824 20682 12880
rect 20534 12416 20590 12472
rect 20626 9424 20682 9480
rect 20442 7948 20498 7984
rect 20442 7928 20444 7948
rect 20444 7928 20496 7948
rect 20496 7928 20498 7948
rect 20074 2352 20130 2408
rect 20810 5752 20866 5808
rect 20350 1400 20406 1456
rect 21362 18128 21418 18184
rect 21086 17720 21142 17776
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21086 17176 21142 17232
rect 21086 16496 21142 16552
rect 21362 16088 21418 16144
rect 21362 15700 21418 15736
rect 21362 15680 21364 15700
rect 21364 15680 21416 15700
rect 21416 15680 21418 15700
rect 21086 15408 21142 15464
rect 21362 14864 21418 14920
rect 21086 14492 21088 14512
rect 21088 14492 21140 14512
rect 21140 14492 21142 14512
rect 21086 14456 21142 14492
rect 21086 13912 21142 13968
rect 21086 13232 21142 13288
rect 21454 13640 21510 13696
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21546 12144 21602 12200
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21546 3440 21602 3496
rect 21178 2624 21234 2680
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21638 1808 21694 1864
rect 22006 992 22062 1048
rect 22006 584 22062 640
<< metal3 >>
rect 0 22266 800 22296
rect 22200 22266 23000 22296
rect 0 22206 2790 22266
rect 0 22176 800 22206
rect 2730 22130 2790 22206
rect 20486 22206 23000 22266
rect 3693 22130 3759 22133
rect 2730 22128 3759 22130
rect 2730 22072 3698 22128
rect 3754 22072 3759 22128
rect 2730 22070 3759 22072
rect 3693 22067 3759 22070
rect 20345 22130 20411 22133
rect 20486 22130 20546 22206
rect 22200 22176 23000 22206
rect 20345 22128 20546 22130
rect 20345 22072 20350 22128
rect 20406 22072 20546 22128
rect 20345 22070 20546 22072
rect 20345 22067 20411 22070
rect 0 21858 800 21888
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 800 21798
rect 4061 21795 4127 21798
rect 20253 21858 20319 21861
rect 22200 21858 23000 21888
rect 20253 21856 23000 21858
rect 20253 21800 20258 21856
rect 20314 21800 23000 21856
rect 20253 21798 23000 21800
rect 20253 21795 20319 21798
rect 22200 21768 23000 21798
rect 0 21450 800 21480
rect 3969 21450 4035 21453
rect 0 21448 4035 21450
rect 0 21392 3974 21448
rect 4030 21392 4035 21448
rect 0 21390 4035 21392
rect 0 21360 800 21390
rect 3969 21387 4035 21390
rect 20621 21450 20687 21453
rect 22200 21450 23000 21480
rect 20621 21448 23000 21450
rect 20621 21392 20626 21448
rect 20682 21392 23000 21448
rect 20621 21390 23000 21392
rect 20621 21387 20687 21390
rect 22200 21360 23000 21390
rect 0 21042 800 21072
rect 3877 21042 3943 21045
rect 0 21040 3943 21042
rect 0 20984 3882 21040
rect 3938 20984 3943 21040
rect 0 20982 3943 20984
rect 0 20952 800 20982
rect 3877 20979 3943 20982
rect 21449 21042 21515 21045
rect 22200 21042 23000 21072
rect 21449 21040 23000 21042
rect 21449 20984 21454 21040
rect 21510 20984 23000 21040
rect 21449 20982 23000 20984
rect 21449 20979 21515 20982
rect 22200 20952 23000 20982
rect 6144 20704 6460 20705
rect 0 20634 800 20664
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 5073 20634 5139 20637
rect 22200 20634 23000 20664
rect 0 20632 5139 20634
rect 0 20576 5078 20632
rect 5134 20576 5139 20632
rect 0 20574 5139 20576
rect 0 20544 800 20574
rect 5073 20571 5139 20574
rect 22142 20544 23000 20634
rect 3969 20498 4035 20501
rect 19425 20498 19491 20501
rect 3969 20496 19491 20498
rect 3969 20440 3974 20496
rect 4030 20440 19430 20496
rect 19486 20440 19491 20496
rect 3969 20438 19491 20440
rect 3969 20435 4035 20438
rect 19425 20435 19491 20438
rect 20989 20498 21055 20501
rect 22142 20498 22202 20544
rect 20989 20496 22202 20498
rect 20989 20440 20994 20496
rect 21050 20440 22202 20496
rect 20989 20438 22202 20440
rect 20989 20435 21055 20438
rect 5901 20362 5967 20365
rect 3374 20360 5967 20362
rect 3374 20304 5906 20360
rect 5962 20304 5967 20360
rect 3374 20302 5967 20304
rect 0 20226 800 20256
rect 3374 20226 3434 20302
rect 5901 20299 5967 20302
rect 0 20166 3434 20226
rect 19701 20226 19767 20229
rect 22200 20226 23000 20256
rect 19701 20224 23000 20226
rect 19701 20168 19706 20224
rect 19762 20168 23000 20224
rect 19701 20166 23000 20168
rect 0 20136 800 20166
rect 19701 20163 19767 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22200 20136 23000 20166
rect 19139 20095 19455 20096
rect 10593 19954 10659 19957
rect 17769 19954 17835 19957
rect 10593 19952 17835 19954
rect 10593 19896 10598 19952
rect 10654 19896 17774 19952
rect 17830 19896 17835 19952
rect 10593 19894 17835 19896
rect 10593 19891 10659 19894
rect 17769 19891 17835 19894
rect 0 19818 800 19848
rect 2313 19818 2379 19821
rect 0 19816 2379 19818
rect 0 19760 2318 19816
rect 2374 19760 2379 19816
rect 0 19758 2379 19760
rect 0 19728 800 19758
rect 2313 19755 2379 19758
rect 5625 19818 5691 19821
rect 7465 19818 7531 19821
rect 5625 19816 7531 19818
rect 5625 19760 5630 19816
rect 5686 19760 7470 19816
rect 7526 19760 7531 19816
rect 5625 19758 7531 19760
rect 5625 19755 5691 19758
rect 7465 19755 7531 19758
rect 21357 19818 21423 19821
rect 22200 19818 23000 19848
rect 21357 19816 23000 19818
rect 21357 19760 21362 19816
rect 21418 19760 23000 19816
rect 21357 19758 23000 19760
rect 21357 19755 21423 19758
rect 22200 19728 23000 19758
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 0 19410 800 19440
rect 1945 19410 2011 19413
rect 0 19408 2011 19410
rect 0 19352 1950 19408
rect 2006 19352 2011 19408
rect 0 19350 2011 19352
rect 0 19320 800 19350
rect 1945 19347 2011 19350
rect 3969 19410 4035 19413
rect 9029 19410 9095 19413
rect 3969 19408 9095 19410
rect 3969 19352 3974 19408
rect 4030 19352 9034 19408
rect 9090 19352 9095 19408
rect 3969 19350 9095 19352
rect 3969 19347 4035 19350
rect 9029 19347 9095 19350
rect 19793 19410 19859 19413
rect 22200 19410 23000 19440
rect 19793 19408 23000 19410
rect 19793 19352 19798 19408
rect 19854 19352 23000 19408
rect 19793 19350 23000 19352
rect 19793 19347 19859 19350
rect 22200 19320 23000 19350
rect 16941 19276 17007 19277
rect 16941 19274 16988 19276
rect 16896 19272 16988 19274
rect 16896 19216 16946 19272
rect 16896 19214 16988 19216
rect 16941 19212 16988 19214
rect 17052 19212 17058 19276
rect 16941 19211 17007 19212
rect 12801 19138 12867 19141
rect 13629 19138 13695 19141
rect 15653 19140 15719 19141
rect 15653 19138 15700 19140
rect 12801 19136 13695 19138
rect 12801 19080 12806 19136
rect 12862 19080 13634 19136
rect 13690 19080 13695 19136
rect 12801 19078 13695 19080
rect 15608 19136 15700 19138
rect 15608 19080 15658 19136
rect 15608 19078 15700 19080
rect 12801 19075 12867 19078
rect 13629 19075 13695 19078
rect 15653 19076 15700 19078
rect 15764 19076 15770 19140
rect 15653 19075 15719 19076
rect 3545 19072 3861 19073
rect 0 19002 800 19032
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 1577 19002 1643 19005
rect 0 19000 1643 19002
rect 0 18944 1582 19000
rect 1638 18944 1643 19000
rect 0 18942 1643 18944
rect 0 18912 800 18942
rect 1577 18939 1643 18942
rect 2773 19002 2839 19005
rect 4797 19002 4863 19005
rect 6453 19002 6519 19005
rect 2773 19000 2882 19002
rect 2773 18944 2778 19000
rect 2834 18944 2882 19000
rect 2773 18939 2882 18944
rect 4797 19000 6519 19002
rect 4797 18944 4802 19000
rect 4858 18944 6458 19000
rect 6514 18944 6519 19000
rect 4797 18942 6519 18944
rect 4797 18939 4863 18942
rect 6453 18939 6519 18942
rect 21449 19002 21515 19005
rect 22200 19002 23000 19032
rect 21449 19000 23000 19002
rect 21449 18944 21454 19000
rect 21510 18944 23000 19000
rect 21449 18942 23000 18944
rect 21449 18939 21515 18942
rect 2822 18730 2882 18939
rect 22200 18912 23000 18942
rect 4153 18866 4219 18869
rect 5717 18866 5783 18869
rect 6729 18866 6795 18869
rect 4153 18864 6795 18866
rect 4153 18808 4158 18864
rect 4214 18808 5722 18864
rect 5778 18808 6734 18864
rect 6790 18808 6795 18864
rect 4153 18806 6795 18808
rect 4153 18803 4219 18806
rect 5717 18803 5783 18806
rect 6729 18803 6795 18806
rect 3141 18730 3207 18733
rect 2822 18728 3207 18730
rect 2822 18672 3146 18728
rect 3202 18672 3207 18728
rect 2822 18670 3207 18672
rect 3141 18667 3207 18670
rect 4521 18730 4587 18733
rect 5717 18730 5783 18733
rect 6085 18730 6151 18733
rect 4521 18728 5783 18730
rect 4521 18672 4526 18728
rect 4582 18672 5722 18728
rect 5778 18672 5783 18728
rect 4521 18670 5783 18672
rect 4521 18667 4587 18670
rect 5717 18667 5783 18670
rect 5950 18728 6151 18730
rect 5950 18672 6090 18728
rect 6146 18672 6151 18728
rect 5950 18670 6151 18672
rect 0 18594 800 18624
rect 1945 18594 2011 18597
rect 0 18592 2011 18594
rect 0 18536 1950 18592
rect 2006 18536 2011 18592
rect 0 18534 2011 18536
rect 0 18504 800 18534
rect 1945 18531 2011 18534
rect 5950 18322 6010 18670
rect 6085 18667 6151 18670
rect 6821 18730 6887 18733
rect 7833 18730 7899 18733
rect 6821 18728 7899 18730
rect 6821 18672 6826 18728
rect 6882 18672 7838 18728
rect 7894 18672 7899 18728
rect 6821 18670 7899 18672
rect 6821 18667 6887 18670
rect 7833 18667 7899 18670
rect 8334 18668 8340 18732
rect 8404 18730 8410 18732
rect 9305 18730 9371 18733
rect 8404 18728 9371 18730
rect 8404 18672 9310 18728
rect 9366 18672 9371 18728
rect 8404 18670 9371 18672
rect 8404 18668 8410 18670
rect 9305 18667 9371 18670
rect 10041 18730 10107 18733
rect 16481 18730 16547 18733
rect 10041 18728 16547 18730
rect 10041 18672 10046 18728
rect 10102 18672 16486 18728
rect 16542 18672 16547 18728
rect 10041 18670 16547 18672
rect 10041 18667 10107 18670
rect 16481 18667 16547 18670
rect 20161 18730 20227 18733
rect 20161 18728 22202 18730
rect 20161 18672 20166 18728
rect 20222 18672 22202 18728
rect 20161 18670 22202 18672
rect 20161 18667 20227 18670
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 11830 18396 11836 18460
rect 11900 18458 11906 18460
rect 12249 18458 12315 18461
rect 11900 18456 12315 18458
rect 11900 18400 12254 18456
rect 12310 18400 12315 18456
rect 11900 18398 12315 18400
rect 11900 18396 11906 18398
rect 12249 18395 12315 18398
rect 6085 18322 6151 18325
rect 5950 18320 6151 18322
rect 5950 18264 6090 18320
rect 6146 18264 6151 18320
rect 5950 18262 6151 18264
rect 6085 18259 6151 18262
rect 6821 18322 6887 18325
rect 10869 18322 10935 18325
rect 6821 18320 10935 18322
rect 6821 18264 6826 18320
rect 6882 18264 10874 18320
rect 10930 18264 10935 18320
rect 6821 18262 10935 18264
rect 6821 18259 6887 18262
rect 10869 18259 10935 18262
rect 12157 18322 12223 18325
rect 12985 18322 13051 18325
rect 12157 18320 13051 18322
rect 12157 18264 12162 18320
rect 12218 18264 12990 18320
rect 13046 18264 13051 18320
rect 12157 18262 13051 18264
rect 12157 18259 12223 18262
rect 12985 18259 13051 18262
rect 0 18186 800 18216
rect 1761 18186 1827 18189
rect 0 18184 1827 18186
rect 0 18128 1766 18184
rect 1822 18128 1827 18184
rect 0 18126 1827 18128
rect 0 18096 800 18126
rect 1761 18123 1827 18126
rect 6637 18188 6703 18189
rect 6637 18184 6684 18188
rect 6748 18186 6754 18188
rect 6637 18128 6642 18184
rect 6637 18124 6684 18128
rect 6748 18126 6794 18186
rect 6748 18124 6754 18126
rect 8518 18124 8524 18188
rect 8588 18186 8594 18188
rect 9397 18186 9463 18189
rect 8588 18184 9463 18186
rect 8588 18128 9402 18184
rect 9458 18128 9463 18184
rect 8588 18126 9463 18128
rect 8588 18124 8594 18126
rect 6637 18123 6703 18124
rect 9397 18123 9463 18126
rect 12065 18186 12131 18189
rect 14273 18186 14339 18189
rect 12065 18184 14339 18186
rect 12065 18128 12070 18184
rect 12126 18128 14278 18184
rect 14334 18128 14339 18184
rect 12065 18126 14339 18128
rect 12065 18123 12131 18126
rect 14273 18123 14339 18126
rect 21357 18186 21423 18189
rect 22200 18186 23000 18216
rect 21357 18184 23000 18186
rect 21357 18128 21362 18184
rect 21418 18128 23000 18184
rect 21357 18126 23000 18128
rect 21357 18123 21423 18126
rect 22200 18096 23000 18126
rect 3182 17988 3188 18052
rect 3252 18050 3258 18052
rect 3417 18050 3483 18053
rect 3252 18048 3483 18050
rect 3252 17992 3422 18048
rect 3478 17992 3483 18048
rect 3252 17990 3483 17992
rect 3252 17988 3258 17990
rect 3417 17987 3483 17990
rect 6637 18050 6703 18053
rect 6913 18050 6979 18053
rect 6637 18048 6979 18050
rect 6637 17992 6642 18048
rect 6698 17992 6918 18048
rect 6974 17992 6979 18048
rect 6637 17990 6979 17992
rect 6637 17987 6703 17990
rect 6913 17987 6979 17990
rect 9254 17988 9260 18052
rect 9324 18050 9330 18052
rect 10317 18050 10383 18053
rect 9324 18048 10383 18050
rect 9324 17992 10322 18048
rect 10378 17992 10383 18048
rect 9324 17990 10383 17992
rect 9324 17988 9330 17990
rect 10317 17987 10383 17990
rect 11605 18050 11671 18053
rect 11830 18050 11836 18052
rect 11605 18048 11836 18050
rect 11605 17992 11610 18048
rect 11666 17992 11836 18048
rect 11605 17990 11836 17992
rect 11605 17987 11671 17990
rect 11830 17988 11836 17990
rect 11900 17988 11906 18052
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 0 17778 800 17808
rect 1761 17778 1827 17781
rect 9121 17778 9187 17781
rect 9990 17778 9996 17780
rect 0 17776 1827 17778
rect 0 17720 1766 17776
rect 1822 17720 1827 17776
rect 0 17718 1827 17720
rect 0 17688 800 17718
rect 1761 17715 1827 17718
rect 2730 17776 9996 17778
rect 2730 17720 9126 17776
rect 9182 17720 9996 17776
rect 2730 17718 9996 17720
rect 1945 17642 2011 17645
rect 2730 17642 2790 17718
rect 9121 17715 9187 17718
rect 9990 17716 9996 17718
rect 10060 17716 10066 17780
rect 21081 17778 21147 17781
rect 22200 17778 23000 17808
rect 21081 17776 23000 17778
rect 21081 17720 21086 17776
rect 21142 17720 23000 17776
rect 21081 17718 23000 17720
rect 21081 17715 21147 17718
rect 22200 17688 23000 17718
rect 1945 17640 2790 17642
rect 1945 17584 1950 17640
rect 2006 17584 2790 17640
rect 1945 17582 2790 17584
rect 6729 17642 6795 17645
rect 8569 17642 8635 17645
rect 6729 17640 8635 17642
rect 6729 17584 6734 17640
rect 6790 17584 8574 17640
rect 8630 17584 8635 17640
rect 6729 17582 8635 17584
rect 1945 17579 2011 17582
rect 6729 17579 6795 17582
rect 8569 17579 8635 17582
rect 6144 17440 6460 17441
rect 0 17370 800 17400
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 1853 17370 1919 17373
rect 22200 17370 23000 17400
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 800 17310
rect 1853 17307 1919 17310
rect 22142 17280 23000 17370
rect 2221 17234 2287 17237
rect 8109 17234 8175 17237
rect 12709 17234 12775 17237
rect 2221 17232 12775 17234
rect 2221 17176 2226 17232
rect 2282 17176 8114 17232
rect 8170 17176 12714 17232
rect 12770 17176 12775 17232
rect 2221 17174 12775 17176
rect 2221 17171 2287 17174
rect 8109 17171 8175 17174
rect 12709 17171 12775 17174
rect 21081 17234 21147 17237
rect 22142 17234 22202 17280
rect 21081 17232 22202 17234
rect 21081 17176 21086 17232
rect 21142 17176 22202 17232
rect 21081 17174 22202 17176
rect 21081 17171 21147 17174
rect 5758 17036 5764 17100
rect 5828 17098 5834 17100
rect 6913 17098 6979 17101
rect 5828 17096 6979 17098
rect 5828 17040 6918 17096
rect 6974 17040 6979 17096
rect 5828 17038 6979 17040
rect 5828 17036 5834 17038
rect 6913 17035 6979 17038
rect 0 16962 800 16992
rect 2773 16962 2839 16965
rect 0 16960 2839 16962
rect 0 16904 2778 16960
rect 2834 16904 2839 16960
rect 0 16902 2839 16904
rect 0 16872 800 16902
rect 2773 16899 2839 16902
rect 5022 16900 5028 16964
rect 5092 16962 5098 16964
rect 5165 16962 5231 16965
rect 5092 16960 5231 16962
rect 5092 16904 5170 16960
rect 5226 16904 5231 16960
rect 5092 16902 5231 16904
rect 5092 16900 5098 16902
rect 5165 16899 5231 16902
rect 5441 16962 5507 16965
rect 5809 16962 5875 16965
rect 7649 16964 7715 16965
rect 5441 16960 5875 16962
rect 5441 16904 5446 16960
rect 5502 16904 5814 16960
rect 5870 16904 5875 16960
rect 5441 16902 5875 16904
rect 5441 16899 5507 16902
rect 5809 16899 5875 16902
rect 7598 16900 7604 16964
rect 7668 16962 7715 16964
rect 20621 16962 20687 16965
rect 22200 16962 23000 16992
rect 7668 16960 7760 16962
rect 7710 16904 7760 16960
rect 7668 16902 7760 16904
rect 20621 16960 23000 16962
rect 20621 16904 20626 16960
rect 20682 16904 23000 16960
rect 20621 16902 23000 16904
rect 7668 16900 7715 16902
rect 7649 16899 7715 16900
rect 20621 16899 20687 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 5574 16628 5580 16692
rect 5644 16690 5650 16692
rect 7005 16690 7071 16693
rect 5644 16688 7071 16690
rect 5644 16632 7010 16688
rect 7066 16632 7071 16688
rect 5644 16630 7071 16632
rect 5644 16628 5650 16630
rect 7005 16627 7071 16630
rect 0 16554 800 16584
rect 1853 16554 1919 16557
rect 0 16552 1919 16554
rect 0 16496 1858 16552
rect 1914 16496 1919 16552
rect 0 16494 1919 16496
rect 0 16464 800 16494
rect 1853 16491 1919 16494
rect 6862 16492 6868 16556
rect 6932 16554 6938 16556
rect 9581 16554 9647 16557
rect 11329 16554 11395 16557
rect 6932 16552 9647 16554
rect 6932 16496 9586 16552
rect 9642 16496 9647 16552
rect 6932 16494 9647 16496
rect 6932 16492 6938 16494
rect 9581 16491 9647 16494
rect 11102 16552 11395 16554
rect 11102 16496 11334 16552
rect 11390 16496 11395 16552
rect 11102 16494 11395 16496
rect 7281 16418 7347 16421
rect 9438 16418 9444 16420
rect 7281 16416 9444 16418
rect 7281 16360 7286 16416
rect 7342 16360 9444 16416
rect 7281 16358 9444 16360
rect 7281 16355 7347 16358
rect 9438 16356 9444 16358
rect 9508 16356 9514 16420
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 0 16146 800 16176
rect 1945 16146 2011 16149
rect 0 16144 2011 16146
rect 0 16088 1950 16144
rect 2006 16088 2011 16144
rect 0 16086 2011 16088
rect 0 16056 800 16086
rect 1945 16083 2011 16086
rect 4981 16146 5047 16149
rect 11102 16146 11162 16494
rect 11329 16491 11395 16494
rect 11973 16554 12039 16557
rect 16757 16554 16823 16557
rect 11973 16552 16823 16554
rect 11973 16496 11978 16552
rect 12034 16496 16762 16552
rect 16818 16496 16823 16552
rect 11973 16494 16823 16496
rect 11973 16491 12039 16494
rect 16757 16491 16823 16494
rect 21081 16554 21147 16557
rect 22200 16554 23000 16584
rect 21081 16552 23000 16554
rect 21081 16496 21086 16552
rect 21142 16496 23000 16552
rect 21081 16494 23000 16496
rect 21081 16491 21147 16494
rect 22200 16464 23000 16494
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 4981 16144 11162 16146
rect 4981 16088 4986 16144
rect 5042 16088 11162 16144
rect 4981 16086 11162 16088
rect 21357 16146 21423 16149
rect 22200 16146 23000 16176
rect 21357 16144 23000 16146
rect 21357 16088 21362 16144
rect 21418 16088 23000 16144
rect 21357 16086 23000 16088
rect 4981 16083 5047 16086
rect 21357 16083 21423 16086
rect 22200 16056 23000 16086
rect 7046 15948 7052 16012
rect 7116 16010 7122 16012
rect 7281 16010 7347 16013
rect 7116 16008 7347 16010
rect 7116 15952 7286 16008
rect 7342 15952 7347 16008
rect 7116 15950 7347 15952
rect 7116 15948 7122 15950
rect 7281 15947 7347 15950
rect 3545 15808 3861 15809
rect 0 15738 800 15768
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 2313 15738 2379 15741
rect 0 15736 2379 15738
rect 0 15680 2318 15736
rect 2374 15680 2379 15736
rect 0 15678 2379 15680
rect 0 15648 800 15678
rect 2313 15675 2379 15678
rect 21357 15738 21423 15741
rect 22200 15738 23000 15768
rect 21357 15736 23000 15738
rect 21357 15680 21362 15736
rect 21418 15680 23000 15736
rect 21357 15678 23000 15680
rect 21357 15675 21423 15678
rect 22200 15648 23000 15678
rect 2589 15604 2655 15605
rect 2589 15600 2636 15604
rect 2700 15602 2706 15604
rect 2589 15544 2594 15600
rect 2589 15540 2636 15544
rect 2700 15542 2746 15602
rect 2700 15540 2706 15542
rect 3366 15540 3372 15604
rect 3436 15602 3442 15604
rect 6361 15602 6427 15605
rect 3436 15600 6427 15602
rect 3436 15544 6366 15600
rect 6422 15544 6427 15600
rect 3436 15542 6427 15544
rect 3436 15540 3442 15542
rect 2589 15539 2655 15540
rect 6361 15539 6427 15542
rect 13905 15466 13971 15469
rect 15101 15466 15167 15469
rect 18505 15466 18571 15469
rect 13905 15464 18571 15466
rect 13905 15408 13910 15464
rect 13966 15408 15106 15464
rect 15162 15408 18510 15464
rect 18566 15408 18571 15464
rect 13905 15406 18571 15408
rect 13905 15403 13971 15406
rect 15101 15403 15167 15406
rect 18505 15403 18571 15406
rect 21081 15466 21147 15469
rect 21081 15464 22202 15466
rect 21081 15408 21086 15464
rect 21142 15408 22202 15464
rect 21081 15406 22202 15408
rect 21081 15403 21147 15406
rect 22142 15360 22202 15406
rect 0 15330 800 15360
rect 1761 15330 1827 15333
rect 0 15328 1827 15330
rect 0 15272 1766 15328
rect 1822 15272 1827 15328
rect 0 15270 1827 15272
rect 0 15240 800 15270
rect 1761 15267 1827 15270
rect 4981 15330 5047 15333
rect 5206 15330 5212 15332
rect 4981 15328 5212 15330
rect 4981 15272 4986 15328
rect 5042 15272 5212 15328
rect 4981 15270 5212 15272
rect 4981 15267 5047 15270
rect 5206 15268 5212 15270
rect 5276 15330 5282 15332
rect 5533 15330 5599 15333
rect 5276 15328 5599 15330
rect 5276 15272 5538 15328
rect 5594 15272 5599 15328
rect 5276 15270 5599 15272
rect 22142 15270 23000 15360
rect 5276 15268 5282 15270
rect 5533 15267 5599 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 6678 15132 6684 15196
rect 6748 15194 6754 15196
rect 6821 15194 6887 15197
rect 6748 15192 9874 15194
rect 6748 15136 6826 15192
rect 6882 15136 9874 15192
rect 6748 15134 9874 15136
rect 6748 15132 6754 15134
rect 6821 15131 6887 15134
rect 2129 15058 2195 15061
rect 7966 15058 7972 15060
rect 2129 15056 7972 15058
rect 2129 15000 2134 15056
rect 2190 15000 7972 15056
rect 2129 14998 7972 15000
rect 2129 14995 2195 14998
rect 7966 14996 7972 14998
rect 8036 15058 8042 15060
rect 9581 15058 9647 15061
rect 9814 15058 9874 15134
rect 14917 15058 14983 15061
rect 8036 15056 9690 15058
rect 8036 15000 9586 15056
rect 9642 15000 9690 15056
rect 8036 14998 9690 15000
rect 9814 15056 14983 15058
rect 9814 15000 14922 15056
rect 14978 15000 14983 15056
rect 9814 14998 14983 15000
rect 8036 14996 8042 14998
rect 9581 14995 9690 14998
rect 14917 14995 14983 14998
rect 0 14922 800 14952
rect 2865 14922 2931 14925
rect 0 14920 2931 14922
rect 0 14864 2870 14920
rect 2926 14864 2931 14920
rect 0 14862 2931 14864
rect 0 14832 800 14862
rect 2865 14859 2931 14862
rect 4061 14922 4127 14925
rect 5390 14922 5396 14924
rect 4061 14920 5396 14922
rect 4061 14864 4066 14920
rect 4122 14864 5396 14920
rect 4061 14862 5396 14864
rect 4061 14859 4127 14862
rect 5390 14860 5396 14862
rect 5460 14922 5466 14924
rect 8661 14922 8727 14925
rect 5460 14920 8727 14922
rect 5460 14864 8666 14920
rect 8722 14864 8727 14920
rect 5460 14862 8727 14864
rect 9630 14922 9690 14995
rect 11053 14922 11119 14925
rect 9630 14920 11119 14922
rect 9630 14864 11058 14920
rect 11114 14864 11119 14920
rect 9630 14862 11119 14864
rect 5460 14860 5466 14862
rect 8661 14859 8727 14862
rect 11053 14859 11119 14862
rect 21357 14922 21423 14925
rect 22200 14922 23000 14952
rect 21357 14920 23000 14922
rect 21357 14864 21362 14920
rect 21418 14864 23000 14920
rect 21357 14862 23000 14864
rect 21357 14859 21423 14862
rect 22200 14832 23000 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 7557 14650 7623 14653
rect 8334 14650 8340 14652
rect 7557 14648 8340 14650
rect 7557 14592 7562 14648
rect 7618 14592 8340 14648
rect 7557 14590 8340 14592
rect 7557 14587 7623 14590
rect 8334 14588 8340 14590
rect 8404 14588 8410 14652
rect 0 14514 800 14544
rect 1577 14514 1643 14517
rect 0 14512 1643 14514
rect 0 14456 1582 14512
rect 1638 14456 1643 14512
rect 0 14454 1643 14456
rect 0 14424 800 14454
rect 1577 14451 1643 14454
rect 21081 14514 21147 14517
rect 22200 14514 23000 14544
rect 21081 14512 23000 14514
rect 21081 14456 21086 14512
rect 21142 14456 23000 14512
rect 21081 14454 23000 14456
rect 21081 14451 21147 14454
rect 22200 14424 23000 14454
rect 3417 14378 3483 14381
rect 7046 14378 7052 14380
rect 3417 14376 7052 14378
rect 3417 14320 3422 14376
rect 3478 14320 7052 14376
rect 3417 14318 7052 14320
rect 3417 14315 3483 14318
rect 7046 14316 7052 14318
rect 7116 14316 7122 14380
rect 3969 14244 4035 14245
rect 3918 14180 3924 14244
rect 3988 14242 4035 14244
rect 8109 14242 8175 14245
rect 8477 14242 8543 14245
rect 3988 14240 4080 14242
rect 4030 14184 4080 14240
rect 3988 14182 4080 14184
rect 8109 14240 8543 14242
rect 8109 14184 8114 14240
rect 8170 14184 8482 14240
rect 8538 14184 8543 14240
rect 8109 14182 8543 14184
rect 3988 14180 4035 14182
rect 3969 14179 4035 14180
rect 8109 14179 8175 14182
rect 8477 14179 8543 14182
rect 6144 14176 6460 14177
rect 0 14106 800 14136
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 2497 14106 2563 14109
rect 0 14104 2563 14106
rect 0 14048 2502 14104
rect 2558 14048 2563 14104
rect 0 14046 2563 14048
rect 0 14016 800 14046
rect 2497 14043 2563 14046
rect 8150 14044 8156 14108
rect 8220 14106 8226 14108
rect 8937 14106 9003 14109
rect 8220 14104 9003 14106
rect 8220 14048 8942 14104
rect 8998 14048 9003 14104
rect 8220 14046 9003 14048
rect 8220 14044 8226 14046
rect 8937 14043 9003 14046
rect 9213 14106 9279 14109
rect 10041 14106 10107 14109
rect 22200 14106 23000 14136
rect 9213 14104 10107 14106
rect 9213 14048 9218 14104
rect 9274 14048 10046 14104
rect 10102 14048 10107 14104
rect 9213 14046 10107 14048
rect 9213 14043 9279 14046
rect 10041 14043 10107 14046
rect 22142 14016 23000 14106
rect 3233 13970 3299 13973
rect 9489 13970 9555 13973
rect 10961 13970 11027 13973
rect 3233 13968 11027 13970
rect 3233 13912 3238 13968
rect 3294 13912 9494 13968
rect 9550 13912 10966 13968
rect 11022 13912 11027 13968
rect 3233 13910 11027 13912
rect 3233 13907 3299 13910
rect 9489 13907 9555 13910
rect 10961 13907 11027 13910
rect 21081 13970 21147 13973
rect 22142 13970 22202 14016
rect 21081 13968 22202 13970
rect 21081 13912 21086 13968
rect 21142 13912 22202 13968
rect 21081 13910 22202 13912
rect 21081 13907 21147 13910
rect 9765 13834 9831 13837
rect 10317 13834 10383 13837
rect 10869 13836 10935 13837
rect 10869 13834 10916 13836
rect 9765 13832 10383 13834
rect 9765 13776 9770 13832
rect 9826 13776 10322 13832
rect 10378 13776 10383 13832
rect 9765 13774 10383 13776
rect 10824 13832 10916 13834
rect 10824 13776 10874 13832
rect 10824 13774 10916 13776
rect 9765 13771 9831 13774
rect 10317 13771 10383 13774
rect 10869 13772 10916 13774
rect 10980 13772 10986 13836
rect 11094 13772 11100 13836
rect 11164 13834 11170 13836
rect 11513 13834 11579 13837
rect 11164 13832 11579 13834
rect 11164 13776 11518 13832
rect 11574 13776 11579 13832
rect 11164 13774 11579 13776
rect 11164 13772 11170 13774
rect 10869 13771 10935 13772
rect 11513 13771 11579 13774
rect 0 13698 800 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 800 13638
rect 1577 13635 1643 13638
rect 9213 13698 9279 13701
rect 9489 13698 9555 13701
rect 9213 13696 9555 13698
rect 9213 13640 9218 13696
rect 9274 13640 9494 13696
rect 9550 13640 9555 13696
rect 9213 13638 9555 13640
rect 9213 13635 9279 13638
rect 9489 13635 9555 13638
rect 14774 13636 14780 13700
rect 14844 13698 14850 13700
rect 16021 13698 16087 13701
rect 14844 13696 16087 13698
rect 14844 13640 16026 13696
rect 16082 13640 16087 13696
rect 14844 13638 16087 13640
rect 14844 13636 14850 13638
rect 16021 13635 16087 13638
rect 21449 13698 21515 13701
rect 22200 13698 23000 13728
rect 21449 13696 23000 13698
rect 21449 13640 21454 13696
rect 21510 13640 23000 13696
rect 21449 13638 23000 13640
rect 21449 13635 21515 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 4245 13426 4311 13429
rect 7741 13426 7807 13429
rect 4245 13424 7807 13426
rect 4245 13368 4250 13424
rect 4306 13368 7746 13424
rect 7802 13368 7807 13424
rect 4245 13366 7807 13368
rect 4245 13363 4311 13366
rect 7741 13363 7807 13366
rect 8385 13426 8451 13429
rect 9857 13426 9923 13429
rect 8385 13424 9923 13426
rect 8385 13368 8390 13424
rect 8446 13368 9862 13424
rect 9918 13368 9923 13424
rect 8385 13366 9923 13368
rect 8385 13363 8451 13366
rect 9857 13363 9923 13366
rect 13721 13426 13787 13429
rect 20529 13426 20595 13429
rect 13721 13424 20595 13426
rect 13721 13368 13726 13424
rect 13782 13368 20534 13424
rect 20590 13368 20595 13424
rect 13721 13366 20595 13368
rect 13721 13363 13787 13366
rect 20529 13363 20595 13366
rect 0 13290 800 13320
rect 1853 13290 1919 13293
rect 0 13288 1919 13290
rect 0 13232 1858 13288
rect 1914 13232 1919 13288
rect 0 13230 1919 13232
rect 0 13200 800 13230
rect 1853 13227 1919 13230
rect 6821 13290 6887 13293
rect 11830 13290 11836 13292
rect 6821 13288 11836 13290
rect 6821 13232 6826 13288
rect 6882 13232 11836 13288
rect 6821 13230 11836 13232
rect 6821 13227 6887 13230
rect 11830 13228 11836 13230
rect 11900 13228 11906 13292
rect 21081 13290 21147 13293
rect 22200 13290 23000 13320
rect 21081 13288 23000 13290
rect 21081 13232 21086 13288
rect 21142 13232 23000 13288
rect 21081 13230 23000 13232
rect 21081 13227 21147 13230
rect 22200 13200 23000 13230
rect 7373 13156 7439 13157
rect 7373 13152 7420 13156
rect 7484 13154 7490 13156
rect 7373 13096 7378 13152
rect 7373 13092 7420 13096
rect 7484 13094 7530 13154
rect 7484 13092 7490 13094
rect 7373 13091 7439 13092
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 0 12882 800 12912
rect 2405 12882 2471 12885
rect 0 12880 2471 12882
rect 0 12824 2410 12880
rect 2466 12824 2471 12880
rect 0 12822 2471 12824
rect 0 12792 800 12822
rect 2405 12819 2471 12822
rect 5073 12882 5139 12885
rect 5625 12882 5691 12885
rect 5073 12880 5691 12882
rect 5073 12824 5078 12880
rect 5134 12824 5630 12880
rect 5686 12824 5691 12880
rect 5073 12822 5691 12824
rect 5073 12819 5139 12822
rect 5625 12819 5691 12822
rect 7925 12882 7991 12885
rect 20621 12882 20687 12885
rect 22200 12882 23000 12912
rect 7925 12880 12450 12882
rect 7925 12824 7930 12880
rect 7986 12824 12450 12880
rect 7925 12822 12450 12824
rect 7925 12819 7991 12822
rect 2681 12746 2747 12749
rect 9857 12746 9923 12749
rect 2681 12744 9923 12746
rect 2681 12688 2686 12744
rect 2742 12688 9862 12744
rect 9918 12688 9923 12744
rect 2681 12686 9923 12688
rect 12390 12746 12450 12822
rect 20621 12880 23000 12882
rect 20621 12824 20626 12880
rect 20682 12824 23000 12880
rect 20621 12822 23000 12824
rect 20621 12819 20687 12822
rect 22200 12792 23000 12822
rect 13721 12746 13787 12749
rect 12390 12744 13787 12746
rect 12390 12688 13726 12744
rect 13782 12688 13787 12744
rect 12390 12686 13787 12688
rect 2681 12683 2747 12686
rect 9857 12683 9923 12686
rect 13721 12683 13787 12686
rect 3545 12544 3861 12545
rect 0 12474 800 12504
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 1577 12474 1643 12477
rect 0 12472 1643 12474
rect 0 12416 1582 12472
rect 1638 12416 1643 12472
rect 0 12414 1643 12416
rect 0 12384 800 12414
rect 1577 12411 1643 12414
rect 10593 12474 10659 12477
rect 17217 12474 17283 12477
rect 10593 12472 12634 12474
rect 10593 12416 10598 12472
rect 10654 12416 12634 12472
rect 10593 12414 12634 12416
rect 10593 12411 10659 12414
rect 4889 12338 4955 12341
rect 10685 12338 10751 12341
rect 12574 12338 12634 12414
rect 14414 12472 17283 12474
rect 14414 12416 17222 12472
rect 17278 12416 17283 12472
rect 14414 12414 17283 12416
rect 12801 12338 12867 12341
rect 14414 12338 14474 12414
rect 17217 12411 17283 12414
rect 20529 12474 20595 12477
rect 22200 12474 23000 12504
rect 20529 12472 23000 12474
rect 20529 12416 20534 12472
rect 20590 12416 23000 12472
rect 20529 12414 23000 12416
rect 20529 12411 20595 12414
rect 22200 12384 23000 12414
rect 4889 12336 6930 12338
rect 4889 12280 4894 12336
rect 4950 12280 6930 12336
rect 4889 12278 6930 12280
rect 4889 12275 4955 12278
rect 5574 12140 5580 12204
rect 5644 12202 5650 12204
rect 5942 12202 5948 12204
rect 5644 12142 5948 12202
rect 5644 12140 5650 12142
rect 5942 12140 5948 12142
rect 6012 12140 6018 12204
rect 6870 12202 6930 12278
rect 10685 12336 12450 12338
rect 10685 12280 10690 12336
rect 10746 12280 12450 12336
rect 10685 12278 12450 12280
rect 12574 12336 14474 12338
rect 12574 12280 12806 12336
rect 12862 12280 14474 12336
rect 12574 12278 14474 12280
rect 15285 12338 15351 12341
rect 16665 12338 16731 12341
rect 15285 12336 16731 12338
rect 15285 12280 15290 12336
rect 15346 12280 16670 12336
rect 16726 12280 16731 12336
rect 15285 12278 16731 12280
rect 10685 12275 10751 12278
rect 12065 12202 12131 12205
rect 6870 12200 12131 12202
rect 6870 12144 12070 12200
rect 12126 12144 12131 12200
rect 6870 12142 12131 12144
rect 12390 12202 12450 12278
rect 12801 12275 12867 12278
rect 15285 12275 15351 12278
rect 16665 12275 16731 12278
rect 16849 12202 16915 12205
rect 12390 12200 16915 12202
rect 12390 12144 16854 12200
rect 16910 12144 16915 12200
rect 12390 12142 16915 12144
rect 12065 12139 12131 12142
rect 16849 12139 16915 12142
rect 21541 12202 21607 12205
rect 21541 12200 22202 12202
rect 21541 12144 21546 12200
rect 21602 12144 22202 12200
rect 21541 12142 22202 12144
rect 21541 12139 21607 12142
rect 22142 12096 22202 12142
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 5625 12068 5691 12069
rect 5574 12066 5580 12068
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 5534 12006 5580 12066
rect 5644 12064 5691 12068
rect 5686 12008 5691 12064
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 5574 12004 5580 12006
rect 5644 12004 5691 12008
rect 22142 12006 23000 12096
rect 5625 12003 5691 12004
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 8293 11932 8359 11933
rect 8293 11928 8340 11932
rect 8404 11930 8410 11932
rect 9397 11930 9463 11933
rect 8293 11872 8298 11928
rect 8293 11868 8340 11872
rect 8404 11870 8450 11930
rect 9397 11928 9690 11930
rect 9397 11872 9402 11928
rect 9458 11872 9690 11928
rect 9397 11870 9690 11872
rect 8404 11868 8410 11870
rect 8293 11867 8359 11868
rect 9397 11867 9463 11870
rect 8569 11796 8635 11797
rect 8518 11794 8524 11796
rect 8478 11734 8524 11794
rect 8588 11792 8635 11796
rect 8630 11736 8635 11792
rect 8518 11732 8524 11734
rect 8588 11732 8635 11736
rect 9630 11794 9690 11870
rect 13353 11794 13419 11797
rect 9630 11792 13419 11794
rect 9630 11736 13358 11792
rect 13414 11736 13419 11792
rect 9630 11734 13419 11736
rect 8569 11731 8635 11732
rect 13353 11731 13419 11734
rect 15469 11794 15535 11797
rect 18781 11794 18847 11797
rect 15469 11792 19350 11794
rect 15469 11736 15474 11792
rect 15530 11736 18786 11792
rect 18842 11736 19350 11792
rect 15469 11734 19350 11736
rect 15469 11731 15535 11734
rect 18781 11731 18847 11734
rect 0 11658 800 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 800 11598
rect 3877 11595 3943 11598
rect 7741 11658 7807 11661
rect 12157 11658 12223 11661
rect 15561 11658 15627 11661
rect 7741 11656 15627 11658
rect 7741 11600 7746 11656
rect 7802 11600 12162 11656
rect 12218 11600 15566 11656
rect 15622 11600 15627 11656
rect 7741 11598 15627 11600
rect 7741 11595 7807 11598
rect 12157 11595 12223 11598
rect 15561 11595 15627 11598
rect 17125 11660 17191 11661
rect 17125 11656 17172 11660
rect 17236 11658 17242 11660
rect 19290 11658 19350 11734
rect 22200 11658 23000 11688
rect 17125 11600 17130 11656
rect 17125 11596 17172 11600
rect 17236 11598 17282 11658
rect 19290 11598 23000 11658
rect 17236 11596 17242 11598
rect 17125 11595 17191 11596
rect 22200 11568 23000 11598
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 0 11250 800 11280
rect 3969 11250 4035 11253
rect 0 11248 4035 11250
rect 0 11192 3974 11248
rect 4030 11192 4035 11248
rect 0 11190 4035 11192
rect 0 11160 800 11190
rect 3969 11187 4035 11190
rect 13813 11250 13879 11253
rect 16113 11250 16179 11253
rect 22200 11250 23000 11280
rect 13813 11248 23000 11250
rect 13813 11192 13818 11248
rect 13874 11192 16118 11248
rect 16174 11192 23000 11248
rect 13813 11190 23000 11192
rect 13813 11187 13879 11190
rect 16113 11187 16179 11190
rect 22200 11160 23000 11190
rect 7005 11114 7071 11117
rect 7230 11114 7236 11116
rect 7005 11112 7236 11114
rect 7005 11056 7010 11112
rect 7066 11056 7236 11112
rect 7005 11054 7236 11056
rect 7005 11051 7071 11054
rect 7230 11052 7236 11054
rect 7300 11052 7306 11116
rect 7966 11052 7972 11116
rect 8036 11114 8042 11116
rect 8201 11114 8267 11117
rect 8036 11112 8267 11114
rect 8036 11056 8206 11112
rect 8262 11056 8267 11112
rect 8036 11054 8267 11056
rect 8036 11052 8042 11054
rect 8201 11051 8267 11054
rect 16297 11114 16363 11117
rect 17493 11114 17559 11117
rect 16297 11112 17559 11114
rect 16297 11056 16302 11112
rect 16358 11056 17498 11112
rect 17554 11056 17559 11112
rect 16297 11054 17559 11056
rect 16297 11051 16363 11054
rect 17493 11051 17559 11054
rect 6144 10912 6460 10913
rect 0 10842 800 10872
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 12249 10842 12315 10845
rect 13813 10842 13879 10845
rect 22200 10842 23000 10872
rect 0 10782 2790 10842
rect 0 10752 800 10782
rect 2730 10706 2790 10782
rect 12249 10840 13879 10842
rect 12249 10784 12254 10840
rect 12310 10784 13818 10840
rect 13874 10784 13879 10840
rect 12249 10782 13879 10784
rect 12249 10779 12315 10782
rect 13813 10779 13879 10782
rect 22142 10752 23000 10842
rect 10317 10706 10383 10709
rect 2730 10704 10383 10706
rect 2730 10648 10322 10704
rect 10378 10648 10383 10704
rect 2730 10646 10383 10648
rect 10317 10643 10383 10646
rect 10869 10706 10935 10709
rect 22142 10706 22202 10752
rect 10869 10704 22202 10706
rect 10869 10648 10874 10704
rect 10930 10648 22202 10704
rect 10869 10646 22202 10648
rect 10869 10643 10935 10646
rect 10409 10570 10475 10573
rect 2270 10568 10475 10570
rect 2270 10512 10414 10568
rect 10470 10512 10475 10568
rect 2270 10510 10475 10512
rect 0 10434 800 10464
rect 2270 10434 2330 10510
rect 10409 10507 10475 10510
rect 11789 10570 11855 10573
rect 12065 10570 12131 10573
rect 11789 10568 12131 10570
rect 11789 10512 11794 10568
rect 11850 10512 12070 10568
rect 12126 10512 12131 10568
rect 11789 10510 12131 10512
rect 11789 10507 11855 10510
rect 12065 10507 12131 10510
rect 16757 10570 16823 10573
rect 18229 10570 18295 10573
rect 16757 10568 18295 10570
rect 16757 10512 16762 10568
rect 16818 10512 18234 10568
rect 18290 10512 18295 10568
rect 16757 10510 18295 10512
rect 16757 10507 16823 10510
rect 18229 10507 18295 10510
rect 0 10374 2330 10434
rect 16481 10434 16547 10437
rect 17350 10434 17356 10436
rect 16481 10432 17356 10434
rect 16481 10376 16486 10432
rect 16542 10376 17356 10432
rect 16481 10374 17356 10376
rect 0 10344 800 10374
rect 16481 10371 16547 10374
rect 17350 10372 17356 10374
rect 17420 10372 17426 10436
rect 22200 10434 23000 10464
rect 19566 10374 23000 10434
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 9213 10298 9279 10301
rect 13077 10298 13143 10301
rect 9213 10296 13143 10298
rect 9213 10240 9218 10296
rect 9274 10240 13082 10296
rect 13138 10240 13143 10296
rect 9213 10238 13143 10240
rect 9213 10235 9279 10238
rect 13077 10235 13143 10238
rect 17033 10298 17099 10301
rect 18045 10298 18111 10301
rect 17033 10296 18111 10298
rect 17033 10240 17038 10296
rect 17094 10240 18050 10296
rect 18106 10240 18111 10296
rect 17033 10238 18111 10240
rect 17033 10235 17099 10238
rect 18045 10235 18111 10238
rect 6637 10162 6703 10165
rect 7046 10162 7052 10164
rect 6637 10160 7052 10162
rect 6637 10104 6642 10160
rect 6698 10104 7052 10160
rect 6637 10102 7052 10104
rect 6637 10099 6703 10102
rect 7046 10100 7052 10102
rect 7116 10100 7122 10164
rect 8201 10162 8267 10165
rect 12934 10162 12940 10164
rect 8201 10160 12940 10162
rect 8201 10104 8206 10160
rect 8262 10104 12940 10160
rect 8201 10102 12940 10104
rect 8201 10099 8267 10102
rect 12934 10100 12940 10102
rect 13004 10162 13010 10164
rect 19566 10162 19626 10374
rect 22200 10344 23000 10374
rect 13004 10102 19626 10162
rect 13004 10100 13010 10102
rect 0 10026 800 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 800 9966
rect 4061 9963 4127 9966
rect 5942 9964 5948 10028
rect 6012 10026 6018 10028
rect 7046 10026 7052 10028
rect 6012 9966 7052 10026
rect 6012 9964 6018 9966
rect 7046 9964 7052 9966
rect 7116 9964 7122 10028
rect 13721 10026 13787 10029
rect 22200 10026 23000 10056
rect 13721 10024 23000 10026
rect 13721 9968 13726 10024
rect 13782 9968 23000 10024
rect 13721 9966 23000 9968
rect 13721 9963 13787 9966
rect 22200 9936 23000 9966
rect 8661 9890 8727 9893
rect 10501 9890 10567 9893
rect 8661 9888 10567 9890
rect 8661 9832 8666 9888
rect 8722 9832 10506 9888
rect 10562 9832 10567 9888
rect 8661 9830 10567 9832
rect 8661 9827 8727 9830
rect 10501 9827 10567 9830
rect 16941 9888 17007 9893
rect 16941 9832 16946 9888
rect 17002 9832 17007 9888
rect 16941 9827 17007 9832
rect 17125 9890 17191 9893
rect 17350 9890 17356 9892
rect 17125 9888 17356 9890
rect 17125 9832 17130 9888
rect 17186 9832 17356 9888
rect 17125 9830 17356 9832
rect 17125 9827 17191 9830
rect 17350 9828 17356 9830
rect 17420 9828 17426 9892
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 16944 9757 17004 9827
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 6545 9754 6611 9757
rect 10685 9754 10751 9757
rect 6545 9752 10751 9754
rect 6545 9696 6550 9752
rect 6606 9696 10690 9752
rect 10746 9696 10751 9752
rect 6545 9694 10751 9696
rect 6545 9691 6611 9694
rect 10685 9691 10751 9694
rect 15745 9754 15811 9757
rect 16389 9754 16455 9757
rect 15745 9752 16455 9754
rect 15745 9696 15750 9752
rect 15806 9696 16394 9752
rect 16450 9696 16455 9752
rect 15745 9694 16455 9696
rect 15745 9691 15811 9694
rect 16389 9691 16455 9694
rect 16941 9752 17007 9757
rect 16941 9696 16946 9752
rect 17002 9696 17007 9752
rect 16941 9691 17007 9696
rect 17217 9754 17283 9757
rect 18413 9754 18479 9757
rect 17217 9752 18479 9754
rect 17217 9696 17222 9752
rect 17278 9696 18418 9752
rect 18474 9696 18479 9752
rect 17217 9694 18479 9696
rect 17217 9691 17283 9694
rect 18413 9691 18479 9694
rect 0 9618 800 9648
rect 4061 9618 4127 9621
rect 0 9616 4127 9618
rect 0 9560 4066 9616
rect 4122 9560 4127 9616
rect 0 9558 4127 9560
rect 0 9528 800 9558
rect 4061 9555 4127 9558
rect 6862 9556 6868 9620
rect 6932 9618 6938 9620
rect 7005 9618 7071 9621
rect 6932 9616 7071 9618
rect 6932 9560 7010 9616
rect 7066 9560 7071 9616
rect 6932 9558 7071 9560
rect 6932 9556 6938 9558
rect 7005 9555 7071 9558
rect 7741 9618 7807 9621
rect 8150 9618 8156 9620
rect 7741 9616 8156 9618
rect 7741 9560 7746 9616
rect 7802 9560 8156 9616
rect 7741 9558 8156 9560
rect 7741 9555 7807 9558
rect 8150 9556 8156 9558
rect 8220 9556 8226 9620
rect 9990 9556 9996 9620
rect 10060 9618 10066 9620
rect 10317 9618 10383 9621
rect 22200 9618 23000 9648
rect 10060 9616 23000 9618
rect 10060 9560 10322 9616
rect 10378 9560 23000 9616
rect 10060 9558 23000 9560
rect 10060 9556 10066 9558
rect 10317 9555 10383 9558
rect 22200 9528 23000 9558
rect 5717 9482 5783 9485
rect 12985 9482 13051 9485
rect 15285 9482 15351 9485
rect 20621 9482 20687 9485
rect 5717 9480 13051 9482
rect 5717 9424 5722 9480
rect 5778 9424 12990 9480
rect 13046 9424 13051 9480
rect 5717 9422 13051 9424
rect 5717 9419 5783 9422
rect 12985 9419 13051 9422
rect 13724 9422 15210 9482
rect 4889 9346 4955 9349
rect 5901 9346 5967 9349
rect 6678 9346 6684 9348
rect 4889 9344 6684 9346
rect 4889 9288 4894 9344
rect 4950 9288 5906 9344
rect 5962 9288 6684 9344
rect 4889 9286 6684 9288
rect 4889 9283 4955 9286
rect 5901 9283 5967 9286
rect 6678 9284 6684 9286
rect 6748 9284 6754 9348
rect 10133 9346 10199 9349
rect 13724 9346 13784 9422
rect 10133 9344 13784 9346
rect 10133 9288 10138 9344
rect 10194 9288 13784 9344
rect 10133 9286 13784 9288
rect 15150 9346 15210 9422
rect 15285 9480 20687 9482
rect 15285 9424 15290 9480
rect 15346 9424 20626 9480
rect 20682 9424 20687 9480
rect 15285 9422 20687 9424
rect 15285 9419 15351 9422
rect 20621 9419 20687 9422
rect 16665 9346 16731 9349
rect 16982 9346 16988 9348
rect 15150 9344 16988 9346
rect 15150 9288 16670 9344
rect 16726 9288 16988 9344
rect 15150 9286 16988 9288
rect 10133 9283 10199 9286
rect 16665 9283 16731 9286
rect 16982 9284 16988 9286
rect 17052 9284 17058 9348
rect 3545 9280 3861 9281
rect 0 9210 800 9240
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9150 3480 9210
rect 0 9120 800 9150
rect 3420 8938 3480 9150
rect 5942 9148 5948 9212
rect 6012 9210 6018 9212
rect 6545 9210 6611 9213
rect 6012 9208 6611 9210
rect 6012 9152 6550 9208
rect 6606 9152 6611 9208
rect 6012 9150 6611 9152
rect 6012 9148 6018 9150
rect 6545 9147 6611 9150
rect 9305 9210 9371 9213
rect 11094 9210 11100 9212
rect 9305 9208 11100 9210
rect 9305 9152 9310 9208
rect 9366 9152 11100 9208
rect 9305 9150 11100 9152
rect 9305 9147 9371 9150
rect 11094 9148 11100 9150
rect 11164 9148 11170 9212
rect 11789 9210 11855 9213
rect 12014 9210 12020 9212
rect 11789 9208 12020 9210
rect 11789 9152 11794 9208
rect 11850 9152 12020 9208
rect 11789 9150 12020 9152
rect 11789 9147 11855 9150
rect 12014 9148 12020 9150
rect 12084 9148 12090 9212
rect 22200 9210 23000 9240
rect 19566 9150 23000 9210
rect 3969 9074 4035 9077
rect 4981 9074 5047 9077
rect 3969 9072 5047 9074
rect 3969 9016 3974 9072
rect 4030 9016 4986 9072
rect 5042 9016 5047 9072
rect 3969 9014 5047 9016
rect 3969 9011 4035 9014
rect 4981 9011 5047 9014
rect 5257 9074 5323 9077
rect 17677 9074 17743 9077
rect 5257 9072 17743 9074
rect 5257 9016 5262 9072
rect 5318 9016 17682 9072
rect 17738 9016 17743 9072
rect 5257 9014 17743 9016
rect 5257 9011 5323 9014
rect 17677 9011 17743 9014
rect 17953 9074 18019 9077
rect 19566 9074 19626 9150
rect 22200 9120 23000 9150
rect 17953 9072 19626 9074
rect 17953 9016 17958 9072
rect 18014 9016 19626 9072
rect 17953 9014 19626 9016
rect 17953 9011 18019 9014
rect 5022 8938 5028 8940
rect 3420 8878 5028 8938
rect 5022 8876 5028 8878
rect 5092 8938 5098 8940
rect 8017 8938 8083 8941
rect 12801 8938 12867 8941
rect 5092 8878 6608 8938
rect 5092 8876 5098 8878
rect 0 8802 800 8832
rect 2957 8802 3023 8805
rect 0 8800 3023 8802
rect 0 8744 2962 8800
rect 3018 8744 3023 8800
rect 0 8742 3023 8744
rect 6548 8802 6608 8878
rect 8017 8936 12867 8938
rect 8017 8880 8022 8936
rect 8078 8880 12806 8936
rect 12862 8880 12867 8936
rect 8017 8878 12867 8880
rect 8017 8875 8083 8878
rect 12801 8875 12867 8878
rect 16849 8938 16915 8941
rect 16982 8938 16988 8940
rect 16849 8936 16988 8938
rect 16849 8880 16854 8936
rect 16910 8880 16988 8936
rect 16849 8878 16988 8880
rect 16849 8875 16915 8878
rect 16982 8876 16988 8878
rect 17052 8876 17058 8940
rect 17953 8938 18019 8941
rect 17953 8936 22202 8938
rect 17953 8880 17958 8936
rect 18014 8880 22202 8936
rect 17953 8878 22202 8880
rect 17953 8875 18019 8878
rect 22142 8832 22202 8878
rect 10041 8802 10107 8805
rect 6548 8800 10107 8802
rect 6548 8744 10046 8800
rect 10102 8744 10107 8800
rect 6548 8742 10107 8744
rect 22142 8742 23000 8832
rect 0 8712 800 8742
rect 2730 8530 2790 8742
rect 2957 8739 3023 8742
rect 10041 8739 10107 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 5349 8668 5415 8669
rect 5349 8666 5396 8668
rect 5304 8664 5396 8666
rect 5304 8608 5354 8664
rect 5304 8606 5396 8608
rect 5349 8604 5396 8606
rect 5460 8604 5466 8668
rect 8201 8666 8267 8669
rect 8661 8666 8727 8669
rect 8201 8664 8727 8666
rect 8201 8608 8206 8664
rect 8262 8608 8666 8664
rect 8722 8608 8727 8664
rect 8201 8606 8727 8608
rect 5349 8603 5415 8604
rect 8201 8603 8267 8606
rect 8661 8603 8727 8606
rect 11789 8666 11855 8669
rect 11789 8664 15348 8666
rect 11789 8608 11794 8664
rect 11850 8608 15348 8664
rect 11789 8606 15348 8608
rect 11789 8603 11855 8606
rect 15142 8530 15148 8532
rect 2730 8470 15148 8530
rect 15142 8468 15148 8470
rect 15212 8468 15218 8532
rect 15288 8530 15348 8606
rect 18689 8530 18755 8533
rect 15288 8528 18755 8530
rect 15288 8472 18694 8528
rect 18750 8472 18755 8528
rect 15288 8470 18755 8472
rect 18689 8467 18755 8470
rect 0 8394 800 8424
rect 3877 8394 3943 8397
rect 0 8392 3943 8394
rect 0 8336 3882 8392
rect 3938 8336 3943 8392
rect 0 8334 3943 8336
rect 0 8304 800 8334
rect 3877 8331 3943 8334
rect 5942 8332 5948 8396
rect 6012 8394 6018 8396
rect 6085 8394 6151 8397
rect 6012 8392 6151 8394
rect 6012 8336 6090 8392
rect 6146 8336 6151 8392
rect 6012 8334 6151 8336
rect 6012 8332 6018 8334
rect 6085 8331 6151 8334
rect 6821 8394 6887 8397
rect 12525 8394 12591 8397
rect 6821 8392 12591 8394
rect 6821 8336 6826 8392
rect 6882 8336 12530 8392
rect 12586 8336 12591 8392
rect 6821 8334 12591 8336
rect 6821 8331 6887 8334
rect 12525 8331 12591 8334
rect 13721 8394 13787 8397
rect 15694 8394 15700 8396
rect 13721 8392 15700 8394
rect 13721 8336 13726 8392
rect 13782 8336 15700 8392
rect 13721 8334 15700 8336
rect 13721 8331 13787 8334
rect 15694 8332 15700 8334
rect 15764 8332 15770 8396
rect 22200 8394 23000 8424
rect 15840 8334 23000 8394
rect 10409 8258 10475 8261
rect 13077 8258 13143 8261
rect 15840 8258 15900 8334
rect 22200 8304 23000 8334
rect 10409 8256 13143 8258
rect 10409 8200 10414 8256
rect 10470 8200 13082 8256
rect 13138 8200 13143 8256
rect 10409 8198 13143 8200
rect 10409 8195 10475 8198
rect 13077 8195 13143 8198
rect 14414 8198 15900 8258
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 2630 8060 2636 8124
rect 2700 8122 2706 8124
rect 2865 8122 2931 8125
rect 2700 8120 2931 8122
rect 2700 8064 2870 8120
rect 2926 8064 2931 8120
rect 2700 8062 2931 8064
rect 2700 8060 2706 8062
rect 2865 8059 2931 8062
rect 10501 8122 10567 8125
rect 10961 8122 11027 8125
rect 10501 8120 11027 8122
rect 10501 8064 10506 8120
rect 10562 8064 10966 8120
rect 11022 8064 11027 8120
rect 10501 8062 11027 8064
rect 10501 8059 10567 8062
rect 10961 8059 11027 8062
rect 0 7986 800 8016
rect 4061 7986 4127 7989
rect 0 7984 4127 7986
rect 0 7928 4066 7984
rect 4122 7928 4127 7984
rect 0 7926 4127 7928
rect 0 7896 800 7926
rect 4061 7923 4127 7926
rect 8334 7924 8340 7988
rect 8404 7986 8410 7988
rect 9397 7986 9463 7989
rect 8404 7984 9463 7986
rect 8404 7928 9402 7984
rect 9458 7928 9463 7984
rect 8404 7926 9463 7928
rect 8404 7924 8410 7926
rect 9397 7923 9463 7926
rect 10910 7924 10916 7988
rect 10980 7986 10986 7988
rect 14414 7986 14474 8198
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 14641 8122 14707 8125
rect 14641 8120 19074 8122
rect 14641 8064 14646 8120
rect 14702 8064 19074 8120
rect 14641 8062 19074 8064
rect 14641 8059 14707 8062
rect 10980 7926 14474 7986
rect 19014 7986 19074 8062
rect 19793 7986 19859 7989
rect 20437 7986 20503 7989
rect 22200 7986 23000 8016
rect 19014 7984 20503 7986
rect 19014 7928 19798 7984
rect 19854 7928 20442 7984
rect 20498 7928 20503 7984
rect 19014 7926 20503 7928
rect 10980 7924 10986 7926
rect 19793 7923 19859 7926
rect 20437 7923 20503 7926
rect 20670 7926 23000 7986
rect 5441 7850 5507 7853
rect 9857 7850 9923 7853
rect 5441 7848 9923 7850
rect 5441 7792 5446 7848
rect 5502 7792 9862 7848
rect 9918 7792 9923 7848
rect 5441 7790 9923 7792
rect 5441 7787 5507 7790
rect 9857 7787 9923 7790
rect 10225 7850 10291 7853
rect 18137 7850 18203 7853
rect 20670 7850 20730 7926
rect 22200 7896 23000 7926
rect 10225 7848 17418 7850
rect 10225 7792 10230 7848
rect 10286 7792 17418 7848
rect 10225 7790 17418 7792
rect 10225 7787 10291 7790
rect 5717 7714 5783 7717
rect 2730 7712 5783 7714
rect 2730 7656 5722 7712
rect 5778 7656 5783 7712
rect 2730 7654 5783 7656
rect 0 7578 800 7608
rect 2730 7578 2790 7654
rect 5717 7651 5783 7654
rect 6678 7652 6684 7716
rect 6748 7714 6754 7716
rect 10133 7714 10199 7717
rect 6748 7712 10199 7714
rect 6748 7656 10138 7712
rect 10194 7656 10199 7712
rect 6748 7654 10199 7656
rect 6748 7652 6754 7654
rect 10133 7651 10199 7654
rect 11789 7714 11855 7717
rect 12341 7714 12407 7717
rect 11789 7712 15026 7714
rect 11789 7656 11794 7712
rect 11850 7656 12346 7712
rect 12402 7656 15026 7712
rect 11789 7654 15026 7656
rect 11789 7651 11855 7654
rect 12341 7651 12407 7654
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 0 7518 2790 7578
rect 7005 7578 7071 7581
rect 7557 7578 7623 7581
rect 14641 7578 14707 7581
rect 7005 7576 8770 7578
rect 7005 7520 7010 7576
rect 7066 7520 7562 7576
rect 7618 7520 8770 7576
rect 7005 7518 8770 7520
rect 0 7488 800 7518
rect 7005 7515 7071 7518
rect 7557 7515 7623 7518
rect 2313 7442 2379 7445
rect 4981 7442 5047 7445
rect 2313 7440 5047 7442
rect 2313 7384 2318 7440
rect 2374 7384 4986 7440
rect 5042 7384 5047 7440
rect 2313 7382 5047 7384
rect 2313 7379 2379 7382
rect 4981 7379 5047 7382
rect 5717 7442 5783 7445
rect 7189 7442 7255 7445
rect 8518 7442 8524 7444
rect 5717 7440 8524 7442
rect 5717 7384 5722 7440
rect 5778 7384 7194 7440
rect 7250 7384 8524 7440
rect 5717 7382 8524 7384
rect 5717 7379 5783 7382
rect 7189 7379 7255 7382
rect 8518 7380 8524 7382
rect 8588 7380 8594 7444
rect 8710 7442 8770 7518
rect 11838 7576 14707 7578
rect 11838 7520 14646 7576
rect 14702 7520 14707 7576
rect 11838 7518 14707 7520
rect 11838 7442 11898 7518
rect 14641 7515 14707 7518
rect 8710 7382 11898 7442
rect 12249 7442 12315 7445
rect 14966 7442 15026 7654
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 17166 7442 17172 7444
rect 12249 7440 14842 7442
rect 12249 7384 12254 7440
rect 12310 7384 14842 7440
rect 12249 7382 14842 7384
rect 14966 7382 17172 7442
rect 12249 7379 12315 7382
rect 3182 7244 3188 7308
rect 3252 7306 3258 7308
rect 5574 7306 5580 7308
rect 3252 7246 5580 7306
rect 3252 7244 3258 7246
rect 5574 7244 5580 7246
rect 5644 7244 5650 7308
rect 5809 7306 5875 7309
rect 14782 7306 14842 7382
rect 17166 7380 17172 7382
rect 17236 7380 17242 7444
rect 17217 7306 17283 7309
rect 5809 7304 14658 7306
rect 5809 7248 5814 7304
rect 5870 7248 14658 7304
rect 5809 7246 14658 7248
rect 14782 7304 17283 7306
rect 14782 7248 17222 7304
rect 17278 7248 17283 7304
rect 14782 7246 17283 7248
rect 17358 7306 17418 7790
rect 18137 7848 20730 7850
rect 18137 7792 18142 7848
rect 18198 7792 20730 7848
rect 18137 7790 20730 7792
rect 18137 7787 18203 7790
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 18505 7578 18571 7581
rect 22200 7578 23000 7608
rect 18505 7576 20362 7578
rect 18505 7520 18510 7576
rect 18566 7520 20362 7576
rect 18505 7518 20362 7520
rect 18505 7515 18571 7518
rect 17953 7442 18019 7445
rect 20302 7442 20362 7518
rect 22142 7488 23000 7578
rect 22142 7442 22202 7488
rect 17953 7440 20132 7442
rect 17953 7384 17958 7440
rect 18014 7384 20132 7440
rect 17953 7382 20132 7384
rect 20302 7382 22202 7442
rect 17953 7379 18019 7382
rect 17358 7246 19994 7306
rect 5809 7243 5875 7246
rect 0 7170 800 7200
rect 1209 7170 1275 7173
rect 0 7168 1275 7170
rect 0 7112 1214 7168
rect 1270 7112 1275 7168
rect 0 7110 1275 7112
rect 0 7080 800 7110
rect 1209 7107 1275 7110
rect 10726 7108 10732 7172
rect 10796 7170 10802 7172
rect 12249 7170 12315 7173
rect 10796 7168 12315 7170
rect 10796 7112 12254 7168
rect 12310 7112 12315 7168
rect 10796 7110 12315 7112
rect 14598 7170 14658 7246
rect 17217 7243 17283 7246
rect 15837 7170 15903 7173
rect 14598 7168 15903 7170
rect 14598 7112 15842 7168
rect 15898 7112 15903 7168
rect 14598 7110 15903 7112
rect 10796 7108 10802 7110
rect 12249 7107 12315 7110
rect 15837 7107 15903 7110
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 14457 7034 14523 7037
rect 17902 7034 17908 7036
rect 14457 7032 17908 7034
rect 14457 6976 14462 7032
rect 14518 6976 17908 7032
rect 14457 6974 17908 6976
rect 14457 6971 14523 6974
rect 17902 6972 17908 6974
rect 17972 6972 17978 7036
rect 3785 6898 3851 6901
rect 5073 6898 5139 6901
rect 3785 6896 5139 6898
rect 3785 6840 3790 6896
rect 3846 6840 5078 6896
rect 5134 6840 5139 6896
rect 3785 6838 5139 6840
rect 3785 6835 3851 6838
rect 5073 6835 5139 6838
rect 5758 6836 5764 6900
rect 5828 6898 5834 6900
rect 6637 6898 6703 6901
rect 5828 6896 6703 6898
rect 5828 6840 6642 6896
rect 6698 6840 6703 6896
rect 5828 6838 6703 6840
rect 5828 6836 5834 6838
rect 6637 6835 6703 6838
rect 9622 6836 9628 6900
rect 9692 6898 9698 6900
rect 12157 6898 12223 6901
rect 12985 6900 13051 6901
rect 9692 6896 12223 6898
rect 9692 6840 12162 6896
rect 12218 6840 12223 6896
rect 9692 6838 12223 6840
rect 9692 6836 9698 6838
rect 12157 6835 12223 6838
rect 12934 6836 12940 6900
rect 13004 6898 13051 6900
rect 13629 6898 13695 6901
rect 15377 6898 15443 6901
rect 13004 6896 13096 6898
rect 13046 6840 13096 6896
rect 13004 6838 13096 6840
rect 13629 6896 15443 6898
rect 13629 6840 13634 6896
rect 13690 6840 15382 6896
rect 15438 6840 15443 6896
rect 13629 6838 15443 6840
rect 13004 6836 13051 6838
rect 12985 6835 13051 6836
rect 13629 6835 13695 6838
rect 15377 6835 15443 6838
rect 17953 6898 18019 6901
rect 17953 6896 19810 6898
rect 17953 6840 17958 6896
rect 18014 6840 19810 6896
rect 17953 6838 19810 6840
rect 17953 6835 18019 6838
rect 0 6762 800 6792
rect 3785 6762 3851 6765
rect 0 6760 3851 6762
rect 0 6704 3790 6760
rect 3846 6704 3851 6760
rect 0 6702 3851 6704
rect 0 6672 800 6702
rect 3785 6699 3851 6702
rect 6269 6762 6335 6765
rect 6453 6762 6519 6765
rect 6862 6762 6868 6764
rect 6269 6760 6868 6762
rect 6269 6704 6274 6760
rect 6330 6704 6458 6760
rect 6514 6704 6868 6760
rect 6269 6702 6868 6704
rect 6269 6699 6335 6702
rect 6453 6699 6519 6702
rect 6862 6700 6868 6702
rect 6932 6700 6938 6764
rect 8753 6762 8819 6765
rect 7422 6760 8819 6762
rect 7422 6704 8758 6760
rect 8814 6704 8819 6760
rect 7422 6702 8819 6704
rect 3049 6626 3115 6629
rect 5073 6626 5139 6629
rect 6637 6628 6703 6629
rect 6637 6626 6684 6628
rect 3049 6624 5139 6626
rect 3049 6568 3054 6624
rect 3110 6568 5078 6624
rect 5134 6568 5139 6624
rect 3049 6566 5139 6568
rect 6592 6624 6684 6626
rect 6748 6626 6754 6628
rect 7422 6626 7482 6702
rect 8753 6699 8819 6702
rect 8937 6762 9003 6765
rect 8937 6760 19626 6762
rect 8937 6704 8942 6760
rect 8998 6704 19626 6760
rect 8937 6702 19626 6704
rect 8937 6699 9003 6702
rect 6592 6568 6642 6624
rect 6592 6566 6684 6568
rect 3049 6563 3115 6566
rect 5073 6563 5139 6566
rect 6637 6564 6684 6566
rect 6748 6566 7482 6626
rect 6748 6564 6754 6566
rect 7598 6564 7604 6628
rect 7668 6626 7674 6628
rect 7741 6626 7807 6629
rect 7668 6624 7807 6626
rect 7668 6568 7746 6624
rect 7802 6568 7807 6624
rect 7668 6566 7807 6568
rect 7668 6564 7674 6566
rect 6637 6563 6703 6564
rect 7741 6563 7807 6566
rect 8385 6626 8451 6629
rect 8937 6626 9003 6629
rect 9622 6626 9628 6628
rect 8385 6624 9628 6626
rect 8385 6568 8390 6624
rect 8446 6568 8942 6624
rect 8998 6568 9628 6624
rect 8385 6566 9628 6568
rect 8385 6563 8451 6566
rect 8937 6563 9003 6566
rect 9622 6564 9628 6566
rect 9692 6564 9698 6628
rect 11973 6626 12039 6629
rect 16205 6626 16271 6629
rect 11973 6624 16271 6626
rect 11973 6568 11978 6624
rect 12034 6568 16210 6624
rect 16266 6568 16271 6624
rect 11973 6566 16271 6568
rect 11973 6563 12039 6566
rect 16205 6563 16271 6566
rect 17033 6626 17099 6629
rect 19425 6626 19491 6629
rect 17033 6624 19491 6626
rect 17033 6568 17038 6624
rect 17094 6568 19430 6624
rect 19486 6568 19491 6624
rect 17033 6566 19491 6568
rect 17033 6563 17099 6566
rect 19425 6563 19491 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 3601 6490 3667 6493
rect 5349 6490 5415 6493
rect 3601 6488 5415 6490
rect 3601 6432 3606 6488
rect 3662 6432 5354 6488
rect 5410 6432 5415 6488
rect 3601 6430 5415 6432
rect 3601 6427 3667 6430
rect 5349 6427 5415 6430
rect 6637 6490 6703 6493
rect 9121 6490 9187 6493
rect 9438 6490 9444 6492
rect 6637 6488 9444 6490
rect 6637 6432 6642 6488
rect 6698 6432 9126 6488
rect 9182 6432 9444 6488
rect 6637 6430 9444 6432
rect 6637 6427 6703 6430
rect 9121 6427 9187 6430
rect 9438 6428 9444 6430
rect 9508 6428 9514 6492
rect 10869 6490 10935 6493
rect 11145 6490 11211 6493
rect 10869 6488 11211 6490
rect 10869 6432 10874 6488
rect 10930 6432 11150 6488
rect 11206 6432 11211 6488
rect 10869 6430 11211 6432
rect 0 6354 800 6384
rect 4061 6354 4127 6357
rect 0 6352 4127 6354
rect 0 6296 4066 6352
rect 4122 6296 4127 6352
rect 0 6294 4127 6296
rect 0 6264 800 6294
rect 4061 6291 4127 6294
rect 6177 6218 6243 6221
rect 2730 6216 6243 6218
rect 2730 6160 6182 6216
rect 6238 6160 6243 6216
rect 2730 6158 6243 6160
rect 9446 6218 9506 6428
rect 10869 6427 10935 6430
rect 11145 6427 11211 6430
rect 12893 6490 12959 6493
rect 16297 6490 16363 6493
rect 12893 6488 16363 6490
rect 12893 6432 12898 6488
rect 12954 6432 16302 6488
rect 16358 6432 16363 6488
rect 12893 6430 16363 6432
rect 12893 6427 12959 6430
rect 16297 6427 16363 6430
rect 9673 6354 9739 6357
rect 9673 6352 19074 6354
rect 9673 6296 9678 6352
rect 9734 6296 19074 6352
rect 9673 6294 19074 6296
rect 9673 6291 9739 6294
rect 16389 6218 16455 6221
rect 9446 6216 16455 6218
rect 9446 6160 16394 6216
rect 16450 6160 16455 6216
rect 9446 6158 16455 6160
rect 0 5946 800 5976
rect 2730 5946 2790 6158
rect 6177 6155 6243 6158
rect 16389 6155 16455 6158
rect 10133 6082 10199 6085
rect 12249 6082 12315 6085
rect 10133 6080 12315 6082
rect 10133 6024 10138 6080
rect 10194 6024 12254 6080
rect 12310 6024 12315 6080
rect 10133 6022 12315 6024
rect 10133 6019 10199 6022
rect 12249 6019 12315 6022
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 0 5886 2790 5946
rect 0 5856 800 5886
rect 5390 5884 5396 5948
rect 5460 5946 5466 5948
rect 6821 5946 6887 5949
rect 5460 5944 6887 5946
rect 5460 5888 6826 5944
rect 6882 5888 6887 5944
rect 5460 5886 6887 5888
rect 5460 5884 5466 5886
rect 6821 5883 6887 5886
rect 9121 5946 9187 5949
rect 9254 5946 9260 5948
rect 9121 5944 9260 5946
rect 9121 5888 9126 5944
rect 9182 5888 9260 5944
rect 9121 5886 9260 5888
rect 9121 5883 9187 5886
rect 9254 5884 9260 5886
rect 9324 5884 9330 5948
rect 11329 5946 11395 5949
rect 10550 5944 11395 5946
rect 10550 5888 11334 5944
rect 11390 5888 11395 5944
rect 10550 5886 11395 5888
rect 5993 5810 6059 5813
rect 8385 5810 8451 5813
rect 10550 5810 10610 5886
rect 11329 5883 11395 5886
rect 10869 5812 10935 5813
rect 10869 5810 10916 5812
rect 5993 5808 8451 5810
rect 5993 5752 5998 5808
rect 6054 5752 8390 5808
rect 8446 5752 8451 5808
rect 5993 5750 8451 5752
rect 5993 5747 6059 5750
rect 8385 5747 8451 5750
rect 9078 5750 10610 5810
rect 10824 5808 10916 5810
rect 10824 5752 10874 5808
rect 10824 5750 10916 5752
rect 4294 5614 6608 5674
rect 0 5538 800 5568
rect 3366 5538 3372 5540
rect 0 5478 3372 5538
rect 0 5448 800 5478
rect 3366 5476 3372 5478
rect 3436 5538 3442 5540
rect 4294 5538 4354 5614
rect 3436 5478 4354 5538
rect 6548 5538 6608 5614
rect 7046 5612 7052 5676
rect 7116 5674 7122 5676
rect 9078 5674 9138 5750
rect 10869 5748 10916 5750
rect 10980 5748 10986 5812
rect 15561 5810 15627 5813
rect 11102 5808 15627 5810
rect 11102 5752 15566 5808
rect 15622 5752 15627 5808
rect 11102 5750 15627 5752
rect 10869 5747 10935 5748
rect 7116 5614 9138 5674
rect 9213 5674 9279 5677
rect 9673 5674 9739 5677
rect 11102 5674 11162 5750
rect 15561 5747 15627 5750
rect 15878 5748 15884 5812
rect 15948 5810 15954 5812
rect 16113 5810 16179 5813
rect 15948 5808 16179 5810
rect 15948 5752 16118 5808
rect 16174 5752 16179 5808
rect 15948 5750 16179 5752
rect 15948 5748 15954 5750
rect 16113 5747 16179 5750
rect 16757 5810 16823 5813
rect 16982 5810 16988 5812
rect 16757 5808 16988 5810
rect 16757 5752 16762 5808
rect 16818 5752 16988 5808
rect 16757 5750 16988 5752
rect 16757 5747 16823 5750
rect 16982 5748 16988 5750
rect 17052 5748 17058 5812
rect 19014 5810 19074 6294
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 19566 5946 19626 6702
rect 19750 6354 19810 6838
rect 19934 6762 19994 7246
rect 20072 7170 20132 7382
rect 22200 7170 23000 7200
rect 20072 7110 23000 7170
rect 22200 7080 23000 7110
rect 22200 6762 23000 6792
rect 19934 6702 23000 6762
rect 22200 6672 23000 6702
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 22200 6354 23000 6384
rect 19750 6294 23000 6354
rect 22200 6264 23000 6294
rect 22200 5946 23000 5976
rect 19566 5886 23000 5946
rect 22200 5856 23000 5886
rect 20805 5810 20871 5813
rect 19014 5808 20871 5810
rect 19014 5752 20810 5808
rect 20866 5752 20871 5808
rect 19014 5750 20871 5752
rect 20805 5747 20871 5750
rect 9213 5672 11162 5674
rect 9213 5616 9218 5672
rect 9274 5616 9678 5672
rect 9734 5616 11162 5672
rect 9213 5614 11162 5616
rect 11329 5674 11395 5677
rect 17401 5674 17467 5677
rect 11329 5672 17467 5674
rect 11329 5616 11334 5672
rect 11390 5616 17406 5672
rect 17462 5616 17467 5672
rect 11329 5614 17467 5616
rect 7116 5612 7122 5614
rect 9213 5611 9279 5614
rect 9673 5611 9739 5614
rect 11329 5611 11395 5614
rect 17401 5611 17467 5614
rect 21590 5614 22202 5674
rect 10726 5538 10732 5540
rect 6548 5478 10732 5538
rect 3436 5476 3442 5478
rect 10726 5476 10732 5478
rect 10796 5538 10802 5540
rect 10869 5538 10935 5541
rect 10796 5536 10935 5538
rect 10796 5480 10874 5536
rect 10930 5480 10935 5536
rect 10796 5478 10935 5480
rect 10796 5476 10802 5478
rect 10869 5475 10935 5478
rect 17033 5538 17099 5541
rect 21590 5538 21650 5614
rect 17033 5536 21650 5538
rect 17033 5480 17038 5536
rect 17094 5480 21650 5536
rect 17033 5478 21650 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 17033 5475 17099 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 5073 5402 5139 5405
rect 5390 5402 5396 5404
rect 5073 5400 5396 5402
rect 5073 5344 5078 5400
rect 5134 5344 5396 5400
rect 5073 5342 5396 5344
rect 5073 5339 5139 5342
rect 5390 5340 5396 5342
rect 5460 5340 5466 5404
rect 6637 5402 6703 5405
rect 14825 5404 14891 5405
rect 6637 5400 10978 5402
rect 6637 5344 6642 5400
rect 6698 5344 10978 5400
rect 6637 5342 10978 5344
rect 6637 5339 6703 5342
rect 3877 5266 3943 5269
rect 10777 5266 10843 5269
rect 3877 5264 10843 5266
rect 3877 5208 3882 5264
rect 3938 5208 10782 5264
rect 10838 5208 10843 5264
rect 3877 5206 10843 5208
rect 10918 5266 10978 5342
rect 14774 5340 14780 5404
rect 14844 5402 14891 5404
rect 14844 5400 14936 5402
rect 14886 5344 14936 5400
rect 14844 5342 14936 5344
rect 14844 5340 14891 5342
rect 14825 5339 14891 5340
rect 15745 5266 15811 5269
rect 10918 5264 15811 5266
rect 10918 5208 15750 5264
rect 15806 5208 15811 5264
rect 10918 5206 15811 5208
rect 3877 5203 3943 5206
rect 10777 5203 10843 5206
rect 15745 5203 15811 5206
rect 0 5130 800 5160
rect 4889 5130 4955 5133
rect 6637 5130 6703 5133
rect 0 5070 4722 5130
rect 0 5040 800 5070
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 0 4722 800 4752
rect 3918 4722 3924 4724
rect 0 4662 3924 4722
rect 0 4632 800 4662
rect 3918 4660 3924 4662
rect 3988 4722 3994 4724
rect 4061 4722 4127 4725
rect 3988 4720 4127 4722
rect 3988 4664 4066 4720
rect 4122 4664 4127 4720
rect 3988 4662 4127 4664
rect 4662 4722 4722 5070
rect 4889 5128 6703 5130
rect 4889 5072 4894 5128
rect 4950 5072 6642 5128
rect 6698 5072 6703 5128
rect 4889 5070 6703 5072
rect 4889 5067 4955 5070
rect 6637 5067 6703 5070
rect 8201 5130 8267 5133
rect 16113 5130 16179 5133
rect 8201 5128 16179 5130
rect 8201 5072 8206 5128
rect 8262 5072 16118 5128
rect 16174 5072 16179 5128
rect 8201 5070 16179 5072
rect 8201 5067 8267 5070
rect 16113 5067 16179 5070
rect 17902 5068 17908 5132
rect 17972 5130 17978 5132
rect 22200 5130 23000 5160
rect 17972 5070 23000 5130
rect 17972 5068 17978 5070
rect 22200 5040 23000 5070
rect 5574 4932 5580 4996
rect 5644 4994 5650 4996
rect 6545 4994 6611 4997
rect 7046 4994 7052 4996
rect 5644 4992 7052 4994
rect 5644 4936 6550 4992
rect 6606 4936 7052 4992
rect 5644 4934 7052 4936
rect 5644 4932 5650 4934
rect 6545 4931 6611 4934
rect 7046 4932 7052 4934
rect 7116 4932 7122 4996
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 10685 4858 10751 4861
rect 13721 4858 13787 4861
rect 10685 4856 13787 4858
rect 10685 4800 10690 4856
rect 10746 4800 13726 4856
rect 13782 4800 13787 4856
rect 10685 4798 13787 4800
rect 10685 4795 10751 4798
rect 13721 4795 13787 4798
rect 9857 4722 9923 4725
rect 15469 4722 15535 4725
rect 4662 4720 9923 4722
rect 4662 4664 9862 4720
rect 9918 4664 9923 4720
rect 4662 4662 9923 4664
rect 3988 4660 3994 4662
rect 4061 4659 4127 4662
rect 9857 4659 9923 4662
rect 10550 4720 15535 4722
rect 10550 4664 15474 4720
rect 15530 4664 15535 4720
rect 10550 4662 15535 4664
rect 5073 4586 5139 4589
rect 5206 4586 5212 4588
rect 5073 4584 5212 4586
rect 5073 4528 5078 4584
rect 5134 4528 5212 4584
rect 5073 4526 5212 4528
rect 5073 4523 5139 4526
rect 5206 4524 5212 4526
rect 5276 4524 5282 4588
rect 9857 4586 9923 4589
rect 10550 4586 10610 4662
rect 15469 4659 15535 4662
rect 17217 4722 17283 4725
rect 22200 4722 23000 4752
rect 17217 4720 23000 4722
rect 17217 4664 17222 4720
rect 17278 4664 23000 4720
rect 17217 4662 23000 4664
rect 17217 4659 17283 4662
rect 22200 4632 23000 4662
rect 9857 4584 10610 4586
rect 9857 4528 9862 4584
rect 9918 4528 10610 4584
rect 9857 4526 10610 4528
rect 10777 4586 10843 4589
rect 13721 4586 13787 4589
rect 10777 4584 13787 4586
rect 10777 4528 10782 4584
rect 10838 4528 13726 4584
rect 13782 4528 13787 4584
rect 10777 4526 13787 4528
rect 9857 4523 9923 4526
rect 10777 4523 10843 4526
rect 13721 4523 13787 4526
rect 10317 4450 10383 4453
rect 11053 4450 11119 4453
rect 10317 4448 11119 4450
rect 10317 4392 10322 4448
rect 10378 4392 11058 4448
rect 11114 4392 11119 4448
rect 10317 4390 11119 4392
rect 10317 4387 10383 4390
rect 11053 4387 11119 4390
rect 11789 4450 11855 4453
rect 12014 4450 12020 4452
rect 11789 4448 12020 4450
rect 11789 4392 11794 4448
rect 11850 4392 12020 4448
rect 11789 4390 12020 4392
rect 11789 4387 11855 4390
rect 12014 4388 12020 4390
rect 12084 4388 12090 4452
rect 6144 4384 6460 4385
rect 0 4314 800 4344
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 22200 4314 23000 4344
rect 0 4254 4906 4314
rect 0 4224 800 4254
rect 4846 4178 4906 4254
rect 22142 4224 23000 4314
rect 8845 4178 8911 4181
rect 4846 4176 8911 4178
rect 4846 4120 8850 4176
rect 8906 4120 8911 4176
rect 4846 4118 8911 4120
rect 8845 4115 8911 4118
rect 10869 4178 10935 4181
rect 14641 4178 14707 4181
rect 10869 4176 14707 4178
rect 10869 4120 10874 4176
rect 10930 4120 14646 4176
rect 14702 4120 14707 4176
rect 10869 4118 14707 4120
rect 10869 4115 10935 4118
rect 14641 4115 14707 4118
rect 15694 4116 15700 4180
rect 15764 4178 15770 4180
rect 18045 4178 18111 4181
rect 15764 4176 18111 4178
rect 15764 4120 18050 4176
rect 18106 4120 18111 4176
rect 15764 4118 18111 4120
rect 15764 4116 15770 4118
rect 18045 4115 18111 4118
rect 18689 4178 18755 4181
rect 22142 4178 22202 4224
rect 18689 4176 22202 4178
rect 18689 4120 18694 4176
rect 18750 4120 22202 4176
rect 18689 4118 22202 4120
rect 18689 4115 18755 4118
rect 7414 3980 7420 4044
rect 7484 4042 7490 4044
rect 8109 4042 8175 4045
rect 7484 4040 8175 4042
rect 7484 3984 8114 4040
rect 8170 3984 8175 4040
rect 7484 3982 8175 3984
rect 7484 3980 7490 3982
rect 8109 3979 8175 3982
rect 8518 3980 8524 4044
rect 8588 4042 8594 4044
rect 9029 4042 9095 4045
rect 8588 4040 9095 4042
rect 8588 3984 9034 4040
rect 9090 3984 9095 4040
rect 8588 3982 9095 3984
rect 8588 3980 8594 3982
rect 9029 3979 9095 3982
rect 11697 4042 11763 4045
rect 17769 4042 17835 4045
rect 11697 4040 17835 4042
rect 11697 3984 11702 4040
rect 11758 3984 17774 4040
rect 17830 3984 17835 4040
rect 11697 3982 17835 3984
rect 11697 3979 11763 3982
rect 17769 3979 17835 3982
rect 17953 4042 18019 4045
rect 17953 4040 19626 4042
rect 17953 3984 17958 4040
rect 18014 3984 19626 4040
rect 17953 3982 19626 3984
rect 17953 3979 18019 3982
rect 0 3906 800 3936
rect 3049 3906 3115 3909
rect 0 3904 3115 3906
rect 0 3848 3054 3904
rect 3110 3848 3115 3904
rect 0 3846 3115 3848
rect 0 3816 800 3846
rect 3049 3843 3115 3846
rect 9673 3906 9739 3909
rect 11513 3906 11579 3909
rect 9673 3904 11579 3906
rect 9673 3848 9678 3904
rect 9734 3848 11518 3904
rect 11574 3848 11579 3904
rect 9673 3846 11579 3848
rect 9673 3843 9739 3846
rect 11513 3843 11579 3846
rect 11697 3906 11763 3909
rect 11830 3906 11836 3908
rect 11697 3904 11836 3906
rect 11697 3848 11702 3904
rect 11758 3848 11836 3904
rect 11697 3846 11836 3848
rect 11697 3843 11763 3846
rect 11830 3844 11836 3846
rect 11900 3844 11906 3908
rect 15142 3844 15148 3908
rect 15212 3906 15218 3908
rect 15377 3906 15443 3909
rect 15212 3904 15443 3906
rect 15212 3848 15382 3904
rect 15438 3848 15443 3904
rect 15212 3846 15443 3848
rect 19566 3906 19626 3982
rect 22200 3906 23000 3936
rect 19566 3846 23000 3906
rect 15212 3844 15218 3846
rect 15377 3843 15443 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 11053 3770 11119 3773
rect 11973 3770 12039 3773
rect 11053 3768 12039 3770
rect 11053 3712 11058 3768
rect 11114 3712 11978 3768
rect 12034 3712 12039 3768
rect 11053 3710 12039 3712
rect 11053 3707 11119 3710
rect 11973 3707 12039 3710
rect 6862 3572 6868 3636
rect 6932 3634 6938 3636
rect 9857 3634 9923 3637
rect 6932 3632 9923 3634
rect 6932 3576 9862 3632
rect 9918 3576 9923 3632
rect 6932 3574 9923 3576
rect 6932 3572 6938 3574
rect 9857 3571 9923 3574
rect 10317 3634 10383 3637
rect 15101 3634 15167 3637
rect 10317 3632 15167 3634
rect 10317 3576 10322 3632
rect 10378 3576 15106 3632
rect 15162 3576 15167 3632
rect 10317 3574 15167 3576
rect 10317 3571 10383 3574
rect 15101 3571 15167 3574
rect 0 3498 800 3528
rect 1761 3498 1827 3501
rect 0 3496 1827 3498
rect 0 3440 1766 3496
rect 1822 3440 1827 3496
rect 0 3438 1827 3440
rect 0 3408 800 3438
rect 1761 3435 1827 3438
rect 5533 3498 5599 3501
rect 5942 3498 5948 3500
rect 5533 3496 5948 3498
rect 5533 3440 5538 3496
rect 5594 3440 5948 3496
rect 5533 3438 5948 3440
rect 5533 3435 5599 3438
rect 5942 3436 5948 3438
rect 6012 3436 6018 3500
rect 6085 3498 6151 3501
rect 18413 3498 18479 3501
rect 6085 3496 18479 3498
rect 6085 3440 6090 3496
rect 6146 3440 18418 3496
rect 18474 3440 18479 3496
rect 6085 3438 18479 3440
rect 6085 3435 6151 3438
rect 18413 3435 18479 3438
rect 21541 3498 21607 3501
rect 22200 3498 23000 3528
rect 21541 3496 23000 3498
rect 21541 3440 21546 3496
rect 21602 3440 23000 3496
rect 21541 3438 23000 3440
rect 21541 3435 21607 3438
rect 22200 3408 23000 3438
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 0 3090 800 3120
rect 1853 3090 1919 3093
rect 0 3088 1919 3090
rect 0 3032 1858 3088
rect 1914 3032 1919 3088
rect 0 3030 1919 3032
rect 0 3000 800 3030
rect 1853 3027 1919 3030
rect 7230 3028 7236 3092
rect 7300 3090 7306 3092
rect 7373 3090 7439 3093
rect 7300 3088 7439 3090
rect 7300 3032 7378 3088
rect 7434 3032 7439 3088
rect 7300 3030 7439 3032
rect 7300 3028 7306 3030
rect 7373 3027 7439 3030
rect 19057 3090 19123 3093
rect 22200 3090 23000 3120
rect 19057 3088 23000 3090
rect 19057 3032 19062 3088
rect 19118 3032 23000 3088
rect 19057 3030 23000 3032
rect 19057 3027 19123 3030
rect 22200 3000 23000 3030
rect 1485 2954 1551 2957
rect 6913 2954 6979 2957
rect 8017 2954 8083 2957
rect 12709 2954 12775 2957
rect 1485 2952 12775 2954
rect 1485 2896 1490 2952
rect 1546 2896 6918 2952
rect 6974 2896 8022 2952
rect 8078 2896 12714 2952
rect 12770 2896 12775 2952
rect 1485 2894 12775 2896
rect 1485 2891 1551 2894
rect 6913 2891 6979 2894
rect 8017 2891 8083 2894
rect 12709 2891 12775 2894
rect 3545 2752 3861 2753
rect 0 2682 800 2712
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 0 2592 800 2622
rect 1577 2619 1643 2622
rect 21173 2682 21239 2685
rect 22200 2682 23000 2712
rect 21173 2680 23000 2682
rect 21173 2624 21178 2680
rect 21234 2624 23000 2680
rect 21173 2622 23000 2624
rect 21173 2619 21239 2622
rect 22200 2592 23000 2622
rect 8845 2546 8911 2549
rect 9254 2546 9260 2548
rect 8845 2544 9260 2546
rect 8845 2488 8850 2544
rect 8906 2488 9260 2544
rect 8845 2486 9260 2488
rect 8845 2483 8911 2486
rect 9254 2484 9260 2486
rect 9324 2484 9330 2548
rect 20069 2410 20135 2413
rect 20069 2408 22202 2410
rect 20069 2352 20074 2408
rect 20130 2352 22202 2408
rect 20069 2350 22202 2352
rect 20069 2347 20135 2350
rect 22142 2304 22202 2350
rect 0 2274 800 2304
rect 2773 2274 2839 2277
rect 0 2272 2839 2274
rect 0 2216 2778 2272
rect 2834 2216 2839 2272
rect 0 2214 2839 2216
rect 0 2184 800 2214
rect 2773 2211 2839 2214
rect 6637 2276 6703 2277
rect 6637 2272 6684 2276
rect 6748 2274 6754 2276
rect 6637 2216 6642 2272
rect 6637 2212 6684 2216
rect 6748 2214 6794 2274
rect 22142 2214 23000 2304
rect 6748 2212 6754 2214
rect 6637 2211 6703 2212
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 0 1866 800 1896
rect 2681 1866 2747 1869
rect 0 1864 2747 1866
rect 0 1808 2686 1864
rect 2742 1808 2747 1864
rect 0 1806 2747 1808
rect 0 1776 800 1806
rect 2681 1803 2747 1806
rect 21633 1866 21699 1869
rect 22200 1866 23000 1896
rect 21633 1864 23000 1866
rect 21633 1808 21638 1864
rect 21694 1808 23000 1864
rect 21633 1806 23000 1808
rect 21633 1803 21699 1806
rect 22200 1776 23000 1806
rect 0 1458 800 1488
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1368 800 1398
rect 3417 1395 3483 1398
rect 20345 1458 20411 1461
rect 22200 1458 23000 1488
rect 20345 1456 23000 1458
rect 20345 1400 20350 1456
rect 20406 1400 23000 1456
rect 20345 1398 23000 1400
rect 20345 1395 20411 1398
rect 22200 1368 23000 1398
rect 0 1050 800 1080
rect 4337 1050 4403 1053
rect 0 1048 4403 1050
rect 0 992 4342 1048
rect 4398 992 4403 1048
rect 0 990 4403 992
rect 0 960 800 990
rect 4337 987 4403 990
rect 22001 1050 22067 1053
rect 22200 1050 23000 1080
rect 22001 1048 23000 1050
rect 22001 992 22006 1048
rect 22062 992 23000 1048
rect 22001 990 23000 992
rect 22001 987 22067 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 3877 642 3943 645
rect 0 640 3943 642
rect 0 584 3882 640
rect 3938 584 3943 640
rect 0 582 3943 584
rect 0 552 800 582
rect 3877 579 3943 582
rect 22001 642 22067 645
rect 22200 642 23000 672
rect 22001 640 23000 642
rect 22001 584 22006 640
rect 22062 584 23000 640
rect 22001 582 23000 584
rect 22001 579 22067 582
rect 22200 552 23000 582
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 16988 19272 17052 19276
rect 16988 19216 17002 19272
rect 17002 19216 17052 19272
rect 16988 19212 17052 19216
rect 15700 19136 15764 19140
rect 15700 19080 15714 19136
rect 15714 19080 15764 19136
rect 15700 19076 15764 19080
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 8340 18668 8404 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 11836 18396 11900 18460
rect 6684 18184 6748 18188
rect 6684 18128 6698 18184
rect 6698 18128 6748 18184
rect 6684 18124 6748 18128
rect 8524 18124 8588 18188
rect 3188 17988 3252 18052
rect 9260 17988 9324 18052
rect 11836 17988 11900 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 9996 17716 10060 17780
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 5764 17036 5828 17100
rect 5028 16900 5092 16964
rect 7604 16960 7668 16964
rect 7604 16904 7654 16960
rect 7654 16904 7668 16960
rect 7604 16900 7668 16904
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 5580 16628 5644 16692
rect 6868 16492 6932 16556
rect 9444 16356 9508 16420
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 7052 15948 7116 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 2636 15600 2700 15604
rect 2636 15544 2650 15600
rect 2650 15544 2700 15600
rect 2636 15540 2700 15544
rect 3372 15540 3436 15604
rect 5212 15268 5276 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 6684 15132 6748 15196
rect 7972 14996 8036 15060
rect 5396 14860 5460 14924
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 8340 14588 8404 14652
rect 7052 14316 7116 14380
rect 3924 14240 3988 14244
rect 3924 14184 3974 14240
rect 3974 14184 3988 14240
rect 3924 14180 3988 14184
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 8156 14044 8220 14108
rect 10916 13832 10980 13836
rect 10916 13776 10930 13832
rect 10930 13776 10980 13832
rect 10916 13772 10980 13776
rect 11100 13772 11164 13836
rect 14780 13636 14844 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 11836 13228 11900 13292
rect 7420 13152 7484 13156
rect 7420 13096 7434 13152
rect 7434 13096 7484 13152
rect 7420 13092 7484 13096
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 5580 12140 5644 12204
rect 5948 12140 6012 12204
rect 5580 12064 5644 12068
rect 5580 12008 5630 12064
rect 5630 12008 5644 12064
rect 5580 12004 5644 12008
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 8340 11928 8404 11932
rect 8340 11872 8354 11928
rect 8354 11872 8404 11928
rect 8340 11868 8404 11872
rect 8524 11792 8588 11796
rect 8524 11736 8574 11792
rect 8574 11736 8588 11792
rect 8524 11732 8588 11736
rect 17172 11656 17236 11660
rect 17172 11600 17186 11656
rect 17186 11600 17236 11656
rect 17172 11596 17236 11600
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 7236 11052 7300 11116
rect 7972 11052 8036 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 17356 10372 17420 10436
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 7052 10100 7116 10164
rect 12940 10100 13004 10164
rect 5948 9964 6012 10028
rect 7052 9964 7116 10028
rect 17356 9828 17420 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 6868 9556 6932 9620
rect 8156 9556 8220 9620
rect 9996 9556 10060 9620
rect 6684 9284 6748 9348
rect 16988 9284 17052 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 5948 9148 6012 9212
rect 11100 9148 11164 9212
rect 12020 9148 12084 9212
rect 5028 8876 5092 8940
rect 16988 8876 17052 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 5396 8664 5460 8668
rect 5396 8608 5410 8664
rect 5410 8608 5460 8664
rect 5396 8604 5460 8608
rect 15148 8468 15212 8532
rect 5948 8332 6012 8396
rect 15700 8332 15764 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 2636 8060 2700 8124
rect 8340 7924 8404 7988
rect 10916 7924 10980 7988
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6684 7652 6748 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 8524 7380 8588 7444
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 3188 7244 3252 7308
rect 5580 7244 5644 7308
rect 17172 7380 17236 7444
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 10732 7108 10796 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 17908 6972 17972 7036
rect 5764 6836 5828 6900
rect 9628 6836 9692 6900
rect 12940 6896 13004 6900
rect 12940 6840 12990 6896
rect 12990 6840 13004 6896
rect 12940 6836 13004 6840
rect 6868 6700 6932 6764
rect 6684 6624 6748 6628
rect 6684 6568 6698 6624
rect 6698 6568 6748 6624
rect 6684 6564 6748 6568
rect 7604 6564 7668 6628
rect 9628 6564 9692 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 9444 6428 9508 6492
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 5396 5884 5460 5948
rect 9260 5884 9324 5948
rect 10916 5808 10980 5812
rect 10916 5752 10930 5808
rect 10930 5752 10980 5808
rect 3372 5476 3436 5540
rect 7052 5612 7116 5676
rect 10916 5748 10980 5752
rect 15884 5748 15948 5812
rect 16988 5748 17052 5812
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 10732 5476 10796 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 5396 5340 5460 5404
rect 14780 5400 14844 5404
rect 14780 5344 14830 5400
rect 14830 5344 14844 5400
rect 14780 5340 14844 5344
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 3924 4660 3988 4724
rect 17908 5068 17972 5132
rect 5580 4932 5644 4996
rect 7052 4932 7116 4996
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 5212 4524 5276 4588
rect 12020 4388 12084 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 15700 4116 15764 4180
rect 7420 3980 7484 4044
rect 8524 3980 8588 4044
rect 11836 3844 11900 3908
rect 15148 3844 15212 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6868 3572 6932 3636
rect 5948 3436 6012 3500
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 7236 3028 7300 3092
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 9260 2484 9324 2548
rect 6684 2272 6748 2276
rect 6684 2216 6698 2272
rect 6698 2216 6748 2272
rect 6684 2212 6748 2216
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3187 18052 3253 18053
rect 3187 17988 3188 18052
rect 3252 17988 3253 18052
rect 3187 17987 3253 17988
rect 2635 15604 2701 15605
rect 2635 15540 2636 15604
rect 2700 15540 2701 15604
rect 2635 15539 2701 15540
rect 2638 8125 2698 15539
rect 2635 8124 2701 8125
rect 2635 8060 2636 8124
rect 2700 8060 2701 8124
rect 2635 8059 2701 8060
rect 3190 7309 3250 17987
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8339 18732 8405 18733
rect 8339 18668 8340 18732
rect 8404 18668 8405 18732
rect 8339 18667 8405 18668
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6683 18188 6749 18189
rect 6683 18124 6684 18188
rect 6748 18124 6749 18188
rect 6683 18123 6749 18124
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5763 17100 5829 17101
rect 5763 17036 5764 17100
rect 5828 17036 5829 17100
rect 5763 17035 5829 17036
rect 5027 16964 5093 16965
rect 5027 16900 5028 16964
rect 5092 16900 5093 16964
rect 5027 16899 5093 16900
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3371 15604 3437 15605
rect 3371 15540 3372 15604
rect 3436 15540 3437 15604
rect 3371 15539 3437 15540
rect 3187 7308 3253 7309
rect 3187 7244 3188 7308
rect 3252 7244 3253 7308
rect 3187 7243 3253 7244
rect 3374 5541 3434 15539
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3923 14244 3989 14245
rect 3923 14180 3924 14244
rect 3988 14180 3989 14244
rect 3923 14179 3989 14180
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3371 5540 3437 5541
rect 3371 5476 3372 5540
rect 3436 5476 3437 5540
rect 3371 5475 3437 5476
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3926 4725 3986 14179
rect 5030 8941 5090 16899
rect 5579 16692 5645 16693
rect 5579 16628 5580 16692
rect 5644 16628 5645 16692
rect 5579 16627 5645 16628
rect 5211 15332 5277 15333
rect 5211 15268 5212 15332
rect 5276 15268 5277 15332
rect 5211 15267 5277 15268
rect 5027 8940 5093 8941
rect 5027 8876 5028 8940
rect 5092 8876 5093 8940
rect 5027 8875 5093 8876
rect 3923 4724 3989 4725
rect 3923 4660 3924 4724
rect 3988 4660 3989 4724
rect 3923 4659 3989 4660
rect 5214 4589 5274 15267
rect 5395 14924 5461 14925
rect 5395 14860 5396 14924
rect 5460 14860 5461 14924
rect 5395 14859 5461 14860
rect 5398 8669 5458 14859
rect 5582 12205 5642 16627
rect 5579 12204 5645 12205
rect 5579 12140 5580 12204
rect 5644 12140 5645 12204
rect 5579 12139 5645 12140
rect 5579 12068 5645 12069
rect 5579 12004 5580 12068
rect 5644 12004 5645 12068
rect 5579 12003 5645 12004
rect 5395 8668 5461 8669
rect 5395 8604 5396 8668
rect 5460 8604 5461 8668
rect 5395 8603 5461 8604
rect 5582 7442 5642 12003
rect 5398 7382 5642 7442
rect 5398 5949 5458 7382
rect 5579 7308 5645 7309
rect 5579 7244 5580 7308
rect 5644 7244 5645 7308
rect 5579 7243 5645 7244
rect 5395 5948 5461 5949
rect 5395 5884 5396 5948
rect 5460 5884 5461 5948
rect 5395 5883 5461 5884
rect 5398 5405 5458 5883
rect 5395 5404 5461 5405
rect 5395 5340 5396 5404
rect 5460 5340 5461 5404
rect 5395 5339 5461 5340
rect 5582 4997 5642 7243
rect 5766 6901 5826 17035
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6686 15197 6746 18123
rect 7603 16964 7669 16965
rect 7603 16900 7604 16964
rect 7668 16900 7669 16964
rect 7603 16899 7669 16900
rect 6867 16556 6933 16557
rect 6867 16492 6868 16556
rect 6932 16492 6933 16556
rect 6867 16491 6933 16492
rect 6683 15196 6749 15197
rect 6683 15132 6684 15196
rect 6748 15132 6749 15196
rect 6683 15131 6749 15132
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5947 12204 6013 12205
rect 5947 12140 5948 12204
rect 6012 12140 6013 12204
rect 5947 12139 6013 12140
rect 5950 10029 6010 12139
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5947 10028 6013 10029
rect 5947 9964 5948 10028
rect 6012 9964 6013 10028
rect 5947 9963 6013 9964
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 5947 9212 6013 9213
rect 5947 9148 5948 9212
rect 6012 9148 6013 9212
rect 5947 9147 6013 9148
rect 5950 8397 6010 9147
rect 6142 8736 6462 9760
rect 6870 9621 6930 16491
rect 7051 16012 7117 16013
rect 7051 15948 7052 16012
rect 7116 15948 7117 16012
rect 7051 15947 7117 15948
rect 7054 14381 7114 15947
rect 7051 14380 7117 14381
rect 7051 14316 7052 14380
rect 7116 14316 7117 14380
rect 7051 14315 7117 14316
rect 7054 10165 7114 14315
rect 7419 13156 7485 13157
rect 7419 13092 7420 13156
rect 7484 13092 7485 13156
rect 7419 13091 7485 13092
rect 7235 11116 7301 11117
rect 7235 11052 7236 11116
rect 7300 11052 7301 11116
rect 7235 11051 7301 11052
rect 7051 10164 7117 10165
rect 7051 10100 7052 10164
rect 7116 10100 7117 10164
rect 7051 10099 7117 10100
rect 7051 10028 7117 10029
rect 7051 9964 7052 10028
rect 7116 9964 7117 10028
rect 7051 9963 7117 9964
rect 6867 9620 6933 9621
rect 6867 9556 6868 9620
rect 6932 9556 6933 9620
rect 6867 9555 6933 9556
rect 6683 9348 6749 9349
rect 6683 9284 6684 9348
rect 6748 9284 6749 9348
rect 6683 9283 6749 9284
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 5947 8396 6013 8397
rect 5947 8332 5948 8396
rect 6012 8332 6013 8396
rect 5947 8331 6013 8332
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 5579 4996 5645 4997
rect 5579 4932 5580 4996
rect 5644 4932 5645 4996
rect 5579 4931 5645 4932
rect 5211 4588 5277 4589
rect 5211 4524 5212 4588
rect 5276 4524 5277 4588
rect 5211 4523 5277 4524
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 5950 3501 6010 8331
rect 6142 7648 6462 8672
rect 6686 7717 6746 9283
rect 7054 9210 7114 9963
rect 6870 9150 7114 9210
rect 6683 7716 6749 7717
rect 6683 7652 6684 7716
rect 6748 7652 6749 7716
rect 6683 7651 6749 7652
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6870 6765 6930 9150
rect 6867 6764 6933 6765
rect 6867 6700 6868 6764
rect 6932 6700 6933 6764
rect 6867 6699 6933 6700
rect 6683 6628 6749 6629
rect 6683 6564 6684 6628
rect 6748 6564 6749 6628
rect 6683 6563 6749 6564
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5947 3500 6013 3501
rect 5947 3436 5948 3500
rect 6012 3436 6013 3500
rect 5947 3435 6013 3436
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6686 2277 6746 6563
rect 6870 3637 6930 6699
rect 7051 5676 7117 5677
rect 7051 5612 7052 5676
rect 7116 5612 7117 5676
rect 7051 5611 7117 5612
rect 7054 4997 7114 5611
rect 7051 4996 7117 4997
rect 7051 4932 7052 4996
rect 7116 4932 7117 4996
rect 7051 4931 7117 4932
rect 6867 3636 6933 3637
rect 6867 3572 6868 3636
rect 6932 3572 6933 3636
rect 6867 3571 6933 3572
rect 7238 3093 7298 11051
rect 7422 4045 7482 13091
rect 7606 6629 7666 16899
rect 7971 15060 8037 15061
rect 7971 14996 7972 15060
rect 8036 14996 8037 15060
rect 7971 14995 8037 14996
rect 7974 11117 8034 14995
rect 8342 14653 8402 18667
rect 8523 18188 8589 18189
rect 8523 18124 8524 18188
rect 8588 18124 8589 18188
rect 8523 18123 8589 18124
rect 8339 14652 8405 14653
rect 8339 14588 8340 14652
rect 8404 14588 8405 14652
rect 8339 14587 8405 14588
rect 8155 14108 8221 14109
rect 8155 14044 8156 14108
rect 8220 14044 8221 14108
rect 8155 14043 8221 14044
rect 7971 11116 8037 11117
rect 7971 11052 7972 11116
rect 8036 11052 8037 11116
rect 7971 11051 8037 11052
rect 8158 9621 8218 14043
rect 8339 11932 8405 11933
rect 8339 11868 8340 11932
rect 8404 11868 8405 11932
rect 8339 11867 8405 11868
rect 8155 9620 8221 9621
rect 8155 9556 8156 9620
rect 8220 9556 8221 9620
rect 8155 9555 8221 9556
rect 8342 7989 8402 11867
rect 8526 11797 8586 18123
rect 8741 17984 9061 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9259 18052 9325 18053
rect 9259 17988 9260 18052
rect 9324 17988 9325 18052
rect 9259 17987 9325 17988
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8523 11796 8589 11797
rect 8523 11732 8524 11796
rect 8588 11732 8589 11796
rect 8523 11731 8589 11732
rect 8741 11456 9061 12480
rect 9262 11930 9322 17987
rect 9995 17780 10061 17781
rect 9995 17716 9996 17780
rect 10060 17716 10061 17780
rect 9995 17715 10061 17716
rect 9443 16420 9509 16421
rect 9443 16356 9444 16420
rect 9508 16356 9509 16420
rect 9443 16355 9509 16356
rect 9446 12450 9506 16355
rect 9446 12390 9690 12450
rect 9262 11870 9506 11930
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8339 7988 8405 7989
rect 8339 7924 8340 7988
rect 8404 7924 8405 7988
rect 8339 7923 8405 7924
rect 8523 7444 8589 7445
rect 8523 7380 8524 7444
rect 8588 7380 8589 7444
rect 8523 7379 8589 7380
rect 7603 6628 7669 6629
rect 7603 6564 7604 6628
rect 7668 6564 7669 6628
rect 7603 6563 7669 6564
rect 8526 4045 8586 7379
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 9446 6493 9506 11870
rect 9630 6901 9690 12390
rect 9998 9621 10058 17715
rect 11340 17440 11660 18464
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 15699 19140 15765 19141
rect 15699 19076 15700 19140
rect 15764 19076 15765 19140
rect 15699 19075 15765 19076
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 11835 18460 11901 18461
rect 11835 18396 11836 18460
rect 11900 18396 11901 18460
rect 11835 18395 11901 18396
rect 11838 18053 11898 18395
rect 11835 18052 11901 18053
rect 11835 17988 11836 18052
rect 11900 17988 11901 18052
rect 11835 17987 11901 17988
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 10915 13836 10981 13837
rect 10915 13772 10916 13836
rect 10980 13772 10981 13836
rect 10915 13771 10981 13772
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 9995 9620 10061 9621
rect 9995 9556 9996 9620
rect 10060 9556 10061 9620
rect 9995 9555 10061 9556
rect 10918 7989 10978 13771
rect 11102 9213 11162 13771
rect 11340 13088 11660 14112
rect 11838 13293 11898 17987
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 14779 13700 14845 13701
rect 14779 13636 14780 13700
rect 14844 13636 14845 13700
rect 14779 13635 14845 13636
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 11835 13292 11901 13293
rect 11835 13228 11836 13292
rect 11900 13228 11901 13292
rect 11835 13227 11901 13228
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11099 9212 11165 9213
rect 11099 9148 11100 9212
rect 11164 9148 11165 9212
rect 11099 9147 11165 9148
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 10915 7988 10981 7989
rect 10915 7924 10916 7988
rect 10980 7924 10981 7988
rect 10915 7923 10981 7924
rect 10731 7172 10797 7173
rect 10731 7108 10732 7172
rect 10796 7108 10797 7172
rect 10731 7107 10797 7108
rect 9627 6900 9693 6901
rect 9627 6836 9628 6900
rect 9692 6836 9693 6900
rect 9627 6835 9693 6836
rect 9630 6629 9690 6835
rect 9627 6628 9693 6629
rect 9627 6564 9628 6628
rect 9692 6564 9693 6628
rect 9627 6563 9693 6564
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 8523 4044 8589 4045
rect 8523 3980 8524 4044
rect 8588 3980 8589 4044
rect 8523 3979 8589 3980
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7235 3092 7301 3093
rect 7235 3028 7236 3092
rect 7300 3028 7301 3092
rect 7235 3027 7301 3028
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 6683 2276 6749 2277
rect 6683 2212 6684 2276
rect 6748 2212 6749 2276
rect 6683 2211 6749 2212
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9262 2549 9322 5883
rect 10734 5541 10794 7107
rect 10918 5813 10978 7923
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 10915 5812 10981 5813
rect 10915 5748 10916 5812
rect 10980 5748 10981 5812
rect 10915 5747 10981 5748
rect 10731 5540 10797 5541
rect 10731 5476 10732 5540
rect 10796 5476 10797 5540
rect 10731 5475 10797 5476
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11838 3909 11898 13227
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 12939 10164 13005 10165
rect 12939 10100 12940 10164
rect 13004 10100 13005 10164
rect 12939 10099 13005 10100
rect 12019 9212 12085 9213
rect 12019 9148 12020 9212
rect 12084 9148 12085 9212
rect 12019 9147 12085 9148
rect 12022 4453 12082 9147
rect 12942 6901 13002 10099
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 12939 6900 13005 6901
rect 12939 6836 12940 6900
rect 13004 6836 13005 6900
rect 12939 6835 13005 6836
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 14782 5405 14842 13635
rect 15702 12450 15762 19075
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 16987 19276 17053 19277
rect 16987 19212 16988 19276
rect 17052 19212 17053 19276
rect 16987 19211 17053 19212
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 15702 12390 15946 12450
rect 15147 8532 15213 8533
rect 15147 8468 15148 8532
rect 15212 8468 15213 8532
rect 15147 8467 15213 8468
rect 14779 5404 14845 5405
rect 14779 5340 14780 5404
rect 14844 5340 14845 5404
rect 14779 5339 14845 5340
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 12019 4452 12085 4453
rect 12019 4388 12020 4452
rect 12084 4388 12085 4452
rect 12019 4387 12085 4388
rect 11835 3908 11901 3909
rect 11835 3844 11836 3908
rect 11900 3844 11901 3908
rect 11835 3843 11901 3844
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9259 2548 9325 2549
rect 9259 2484 9260 2548
rect 9324 2484 9325 2548
rect 9259 2483 9325 2484
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 3840 14259 4864
rect 15150 3909 15210 8467
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 15702 4181 15762 8331
rect 15886 5813 15946 12390
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16990 9349 17050 19211
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 17171 11660 17237 11661
rect 17171 11596 17172 11660
rect 17236 11596 17237 11660
rect 17171 11595 17237 11596
rect 16987 9348 17053 9349
rect 16987 9284 16988 9348
rect 17052 9284 17053 9348
rect 16987 9283 17053 9284
rect 16987 8940 17053 8941
rect 16987 8876 16988 8940
rect 17052 8876 17053 8940
rect 16987 8875 17053 8876
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 15883 5812 15949 5813
rect 15883 5748 15884 5812
rect 15948 5748 15949 5812
rect 15883 5747 15949 5748
rect 16538 5472 16858 6496
rect 16990 5813 17050 8875
rect 17174 7445 17234 11595
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 17355 10436 17421 10437
rect 17355 10372 17356 10436
rect 17420 10372 17421 10436
rect 17355 10371 17421 10372
rect 17358 9893 17418 10371
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 17355 9892 17421 9893
rect 17355 9828 17356 9892
rect 17420 9828 17421 9892
rect 17355 9827 17421 9828
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 17171 7444 17237 7445
rect 17171 7380 17172 7444
rect 17236 7380 17237 7444
rect 17171 7379 17237 7380
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 17907 7036 17973 7037
rect 17907 6972 17908 7036
rect 17972 6972 17973 7036
rect 17907 6971 17973 6972
rect 16987 5812 17053 5813
rect 16987 5748 16988 5812
rect 17052 5748 17053 5812
rect 16987 5747 17053 5748
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 17910 5133 17970 6971
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 17907 5132 17973 5133
rect 17907 5068 17908 5132
rect 17972 5068 17973 5132
rect 17907 5067 17973 5068
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 15699 4180 15765 4181
rect 15699 4116 15700 4180
rect 15764 4116 15765 4180
rect 15699 4115 15765 4116
rect 15147 3908 15213 3909
rect 15147 3844 15148 3908
rect 15212 3844 15213 3908
rect 15147 3843 15213 3844
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform -1 0 2392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1649977179
transform -1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 1656 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 1656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform -1 0 2392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1649977179
transform -1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1649977179
transform 1 0 20608 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1649977179
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 21344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1649977179
transform -1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform -1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 11776 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 13892 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform -1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 14260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1649977179
transform -1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1649977179
transform -1 0 15456 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1649977179
transform -1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1649977179
transform 1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_E_FTB01_A
timestamp 1649977179
transform -1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_W_FTB01_A
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_E_FTB01_A
timestamp 1649977179
transform 1 0 18400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_N_FTB01_A
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 20700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_W_FTB01_A
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_E_FTB01_A
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_S_FTB01_A
timestamp 1649977179
transform 1 0 20148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_W_FTB01_A
timestamp 1649977179
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_delay_buf_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4048 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 3128 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 3680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4__CLK
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1649977179
transform -1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 6440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1649977179
transform 1 0 6624 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12052 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 10580 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 1472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6716 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2852 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 19136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18308 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 21160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 21620 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1649977179
transform -1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1649977179
transform 1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1649977179
transform -1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 19044 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 17848 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 19044 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 19044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 21620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 6716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1649977179
transform 1 0 3128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4048 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4048 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6256 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1649977179
transform -1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1649977179
transform -1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1649977179
transform -1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1649977179
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6348 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 13524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13064 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 11040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14904 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13064 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 21620 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_E_FTB01_A
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_W_FTB01_A
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 20148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1649977179
transform -1 0 18768 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1649977179
transform -1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_S_FTB01_A
timestamp 1649977179
transform -1 0 21620 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96
timestamp 1649977179
transform 1 0 9936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_153
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_9
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_43
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_119
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1649977179
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1649977179
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_212
timestamp 1649977179
transform 1 0 20608 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_100
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_165
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_5
timestamp 1649977179
transform 1 0 1564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_183
timestamp 1649977179
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_193
timestamp 1649977179
transform 1 0 18860 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_88
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_136
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_54
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_161
timestamp 1649977179
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_172
timestamp 1649977179
transform 1 0 16928 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_38
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_187
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_31
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1649977179
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_186
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1649977179
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_122
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1649977179
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1649977179
transform 1 0 21528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_150
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_120
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1649977179
transform 1 0 19412 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1649977179
transform 1 0 20516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_16
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_201
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_218
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_50
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1649977179
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_218
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1649977179
transform 1 0 21528 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1649977179
transform 1 0 4048 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1649977179
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_24
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_218
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_222
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_58
timestamp 1649977179
transform 1 0 6440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_179
timestamp 1649977179
transform 1 0 17572 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_201
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_41
timestamp 1649977179
transform 1 0 4876 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_124
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_143
timestamp 1649977179
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_171
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_201
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_208
timestamp 1649977179
transform 1 0 20240 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_22
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_36
timestamp 1649977179
transform 1 0 4416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_51
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1649977179
transform 1 0 6808 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_148
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1649977179
transform 1 0 16100 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1649977179
transform 1 0 2576 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_201
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_72
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_100
timestamp 1649977179
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_179
timestamp 1649977179
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1649977179
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1649977179
transform 1 0 20516 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_44
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_130
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_183
timestamp 1649977179
transform 1 0 17940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_195
timestamp 1649977179
transform 1 0 19044 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_31
timestamp 1649977179
transform 1 0 3956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1649977179
transform 1 0 7728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_94
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_14
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_100
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1649977179
transform 1 0 15364 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_81
timestamp 1649977179
transform 1 0 8556 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_150
timestamp 1649977179
transform 1 0 14904 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_162
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_186
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1649977179
transform 1 0 19412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1649977179
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_16
timestamp 1649977179
transform 1 0 2576 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 1649977179
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_156
timestamp 1649977179
transform 1 0 15456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1649977179
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_73
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_117
timestamp 1649977179
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_129
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_154
timestamp 1649977179
transform 1 0 15272 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_177
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _028_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1649977179
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1649977179
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1649977179
transform -1 0 17204 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1649977179
transform -1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform -1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform -1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1649977179
transform -1 0 1840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1649977179
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1649977179
transform -1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1649977179
transform -1 0 1840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1649977179
transform -1 0 2760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1649977179
transform -1 0 1840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1649977179
transform -1 0 3128 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1649977179
transform -1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1649977179
transform -1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform -1 0 2024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 2024 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform -1 0 1840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform -1 0 2576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform 1 0 20884 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform 1 0 21160 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform -1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform -1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1649977179
transform 1 0 10856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1649977179
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1649977179
transform -1 0 13708 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1649977179
transform -1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1649977179
transform 1 0 13156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1649977179
transform -1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1649977179
transform 1 0 14720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1649977179
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1649977179
transform -1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1649977179
transform -1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_1_E_FTB01
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_1_W_FTB01
timestamp 1649977179
transform -1 0 18216 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1649977179
transform -1 0 17112 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1649977179
transform -1 0 17664 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_16  delay_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6164 0 -1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17480 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12052 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12880 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11960 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9844 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5980 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3220 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1472 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4600 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6440 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3128 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2944 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5152 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19872 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17940 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20884 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16284 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19872 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16744 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2576 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2024 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4692 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5888 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5336 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6900 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10488 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12144 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13156 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14168 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14536 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13340 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15732 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 13064 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13616 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12788 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11868 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 11316 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 11316 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8832 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9844 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10304 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 7636 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1649977179
transform -1 0 7636 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1649977179
transform -1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8740 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10580 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9016 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8372 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12052 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12880 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13432 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13616 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16192 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6532 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5520 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3864 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2760 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1649977179
transform 1 0 1564 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7544 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5152 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5980 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5704 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3220 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3680 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16836 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1649977179
transform -1 0 15180 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18124 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20424 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1649977179
transform -1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19504 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20240 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1649977179
transform -1 0 21252 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1649977179
transform -1 0 13248 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1649977179
transform -1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20976 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1649977179
transform 1 0 19872 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 20148 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1649977179
transform -1 0 20332 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14720 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15364 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16376 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17204 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18676 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 17848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19412 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15916 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15272 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2668 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4324 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9016 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6808 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5336 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7452 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1649977179
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1649977179
transform 1 0 9108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1649977179
transform 1 0 8188 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1649977179
transform -1 0 8832 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8280 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1649977179
transform -1 0 9108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1649977179
transform -1 0 8832 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1649977179
transform 1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10488 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6900 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10764 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9384 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12972 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12972 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16192 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15916 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16284 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15364 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15640 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_E_FTB01
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_W_FTB01
timestamp 1649977179
transform -1 0 19780 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1649977179
transform 1 0 20056 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1649977179
transform 1 0 19504 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1649977179
transform -1 0 18768 0 1 19584
box -38 -48 590 592
<< labels >>
flabel metal2 s 18234 22200 18290 23000 0 FreeSans 224 90 0 0 Test_en_N_out
port 0 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 1 nsew signal input
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal2 s 3514 22200 3570 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 134 nsew signal input
flabel metal2 s 7194 22200 7250 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 135 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 136 nsew signal input
flabel metal2 s 7930 22200 7986 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 137 nsew signal input
flabel metal2 s 8298 22200 8354 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 138 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 139 nsew signal input
flabel metal2 s 9034 22200 9090 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 140 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 141 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 142 nsew signal input
flabel metal2 s 10138 22200 10194 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 143 nsew signal input
flabel metal2 s 10506 22200 10562 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 144 nsew signal input
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 145 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 146 nsew signal input
flabel metal2 s 4618 22200 4674 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 147 nsew signal input
flabel metal2 s 4986 22200 5042 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 148 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 149 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 150 nsew signal input
flabel metal2 s 6090 22200 6146 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 151 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 152 nsew signal input
flabel metal2 s 6826 22200 6882 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 153 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 154 nsew signal tristate
flabel metal2 s 14554 22200 14610 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 155 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 156 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 157 nsew signal tristate
flabel metal2 s 15658 22200 15714 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 158 nsew signal tristate
flabel metal2 s 16026 22200 16082 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 159 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 160 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 161 nsew signal tristate
flabel metal2 s 17130 22200 17186 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 162 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 163 nsew signal tristate
flabel metal2 s 17866 22200 17922 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 164 nsew signal tristate
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 165 nsew signal tristate
flabel metal2 s 11610 22200 11666 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 166 nsew signal tristate
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 167 nsew signal tristate
flabel metal2 s 12346 22200 12402 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 168 nsew signal tristate
flabel metal2 s 12714 22200 12770 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 169 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 170 nsew signal tristate
flabel metal2 s 13450 22200 13506 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 171 nsew signal tristate
flabel metal2 s 13818 22200 13874 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 172 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 173 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 clk_1_E_out
port 174 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 clk_1_N_in
port 175 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 clk_1_W_out
port 176 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 clk_2_E_out
port 177 nsew signal tristate
flabel metal2 s 18970 22200 19026 23000 0 FreeSans 224 90 0 0 clk_2_N_in
port 178 nsew signal input
flabel metal2 s 21178 22200 21234 23000 0 FreeSans 224 90 0 0 clk_2_N_out
port 179 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 clk_2_S_out
port 180 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 clk_2_W_out
port 181 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 clk_3_E_out
port 182 nsew signal tristate
flabel metal2 s 19338 22200 19394 23000 0 FreeSans 224 90 0 0 clk_3_N_in
port 183 nsew signal input
flabel metal2 s 21546 22200 21602 23000 0 FreeSans 224 90 0 0 clk_3_N_out
port 184 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 clk_3_S_out
port 185 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 clk_3_W_out
port 186 nsew signal tristate
flabel metal3 s 0 552 800 672 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 187 nsew signal input
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 188 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 189 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 190 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 191 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 192 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 193 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 194 nsew signal input
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 195 nsew signal input
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 prog_clk_1_E_out
port 196 nsew signal tristate
flabel metal2 s 20074 22200 20130 23000 0 FreeSans 224 90 0 0 prog_clk_1_N_in
port 197 nsew signal input
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 prog_clk_1_W_out
port 198 nsew signal tristate
flabel metal3 s 22200 21768 23000 21888 0 FreeSans 480 0 0 0 prog_clk_2_E_out
port 199 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_in
port 200 nsew signal input
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_out
port 201 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 prog_clk_2_S_out
port 202 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prog_clk_2_W_out
port 203 nsew signal tristate
flabel metal3 s 22200 22176 23000 22296 0 FreeSans 480 0 0 0 prog_clk_3_E_out
port 204 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_in
port 205 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 206 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 prog_clk_3_S_out
port 207 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 prog_clk_3_W_out
port 208 nsew signal tristate
flabel metal3 s 22200 552 23000 672 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 209 nsew signal input
flabel metal3 s 22200 960 23000 1080 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 210 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 211 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 212 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 213 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 214 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 215 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 216 nsew signal input
flabel metal2 s 570 22200 626 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 217 nsew signal input
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 218 nsew signal input
flabel metal2 s 1306 22200 1362 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 219 nsew signal input
flabel metal2 s 1674 22200 1730 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 220 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 221 nsew signal input
flabel metal2 s 2410 22200 2466 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 222 nsew signal input
flabel metal2 s 2778 22200 2834 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 223 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 224 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
