* NGSPICE file created from sb_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

.subckt sb_1__1_ Test_en_N_out Test_en_S_in VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] clk_1_E_out clk_1_N_in clk_1_W_out clk_2_E_out clk_2_N_in clk_2_N_out
+ clk_2_S_out clk_2_W_out clk_3_E_out clk_3_N_in clk_3_N_out clk_3_S_out clk_3_W_out
+ left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_ left_bottom_grid_pin_37_
+ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_ left_bottom_grid_pin_41_
+ prog_clk_0_N_in prog_clk_1_E_out prog_clk_1_N_in prog_clk_1_W_out prog_clk_2_E_out
+ prog_clk_2_N_in prog_clk_2_N_out prog_clk_2_S_out prog_clk_2_W_out prog_clk_3_E_out
+ prog_clk_3_N_in prog_clk_3_N_out prog_clk_3_S_out prog_clk_3_W_out right_bottom_grid_pin_34_
+ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_
+ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_ right_bottom_grid_pin_41_ top_left_grid_pin_42_
+ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_
+ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ repeater270/X mux_right_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater229/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input92_A clk_2_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_1_ input33/X _061_/A repeater237/X VGND VGND VPWR VPWR
+ mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ repeater252/X mux_left_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l1_in_3__297 VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_3_/A0
+ mux_bottom_track_33.mux_l1_in_3__297/LO sky130_fd_sc_hd__conb_1
XFILLER_18_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput220 output220/A VGND VGND VPWR VPWR prog_clk_3_N_out sky130_fd_sc_hd__buf_2
X_062_ _062_/A VGND VGND VPWR VPWR _062_/X sky130_fd_sc_hd__clkbuf_1
X_131_ _131_/A VGND VGND VPWR VPWR _131_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input55_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ repeater266/X mux_right_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_3__279 VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/A0
+ mux_right_track_0.mux_l2_in_3__279/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ repeater261/X mux_bottom_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_0_ _114_/A _105_/A mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input18_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_4__A1 _129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
Xinput120 top_left_grid_pin_49_ VGND VGND VPWR VPWR input120/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__127__A _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_3__296 VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/A0
+ mux_bottom_track_3.mux_l2_in_3__296/LO sky130_fd_sc_hd__conb_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_ repeater243/X mux_bottom_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_0.mux_l2_in_3__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input85_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_0_ _110_/A _101_/A repeater237/A VGND VGND VPWR VPWR
+ mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_3__282 VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_3_/A0
+ mux_right_track_24.mux_l2_in_3__282/LO sky130_fd_sc_hd__conb_1
Xoutput210 output210/A VGND VGND VPWR VPWR clk_3_N_out sky130_fd_sc_hd__buf_2
Xoutput221 output221/A VGND VGND VPWR VPWR prog_clk_3_S_out sky130_fd_sc_hd__buf_2
X_130_ _130_/A VGND VGND VPWR VPWR _130_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A0 _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_061_ _061_/A VGND VGND VPWR VPWR _061_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input48_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ repeater273/X mux_right_track_4.mux_l5_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xprog_clk_2_W_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR output218/A sky130_fd_sc_hd__buf_4
XANTENNA__135__A _135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _060_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input102_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ repeater247/X mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_ repeater258/X mux_top_track_16.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput110 right_bottom_grid_pin_39_ VGND VGND VPWR VPWR input110/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 _061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_3_ mux_right_track_8.mux_l2_in_3_/A0 _093_/A mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input30_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_3_ mux_top_track_0.mux_l2_in_3_/A0 _089_/A mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ repeater244/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l2_in_2__A1 _133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input78_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_3__A1 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_4_ input11/X _129_/A repeater226/A VGND VGND VPWR VPWR
+ mux_top_track_0.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xoutput200 _123_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput211 output211/A VGND VGND VPWR VPWR clk_3_S_out sky130_fd_sc_hd__buf_2
Xoutput222 output222/A VGND VGND VPWR VPWR prog_clk_3_W_out sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_060_ _060_/A VGND VGND VPWR VPWR _060_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_ repeater264/X mux_bottom_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__061__A _061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input60_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ repeater247/X mux_bottom_track_17.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclk_2_E_FTB01 input92/X VGND VGND VPWR VPWR output205/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ repeater258/X mux_top_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput111 right_bottom_grid_pin_40_ VGND VGND VPWR VPWR input111/X sky130_fd_sc_hd__clkbuf_1
Xinput100 left_bottom_grid_pin_40_ VGND VGND VPWR VPWR input100/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_8.mux_l2_in_2_ _083_/A _133_/A mux_right_track_8.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input23_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ _079_/A mux_top_track_0.mux_l1_in_4_/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ repeater243/X repeater237/X VGND VGND
+ VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_0.mux_l1_in_3__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_3_ _119_/A _069_/A repeater226/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input90_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput201 _124_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xoutput212 output212/A VGND VGND VPWR VPWR clk_3_W_out sky130_fd_sc_hd__buf_2
XANTENNA__059__A _059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_0_FTB00 input102/X VGND VGND VPWR VPWR repeater275/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ repeater264/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input53_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_3__285 VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/A0
+ mux_right_track_8.mux_l2_in_3__285/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xprog_clk_3_N_FTB01 input104/X VGND VGND VPWR VPWR output220/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_3.mux_l1_in_4__A0 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ repeater254/X mux_top_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__067__A _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput101 left_bottom_grid_pin_41_ VGND VGND VPWR VPWR input101/X sky130_fd_sc_hd__clkbuf_1
Xinput112 right_bottom_grid_pin_41_ VGND VGND VPWR VPWR input112/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input16_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l2_in_1_ _123_/A mux_right_track_8.mux_l1_in_2_/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ mux_top_track_0.mux_l1_in_3_/X mux_top_track_0.mux_l1_in_2_/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ repeater262/X mux_bottom_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater237/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 _059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A bottom_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l1_in_2_ input64/X input109/X mux_right_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_3__A1 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_2_ _059_/A input42/X repeater226/A VGND VGND VPWR VPWR
+ mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input118_A top_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input83_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput213 output213/A VGND VGND VPWR VPWR prog_clk_1_E_out sky130_fd_sc_hd__buf_2
Xoutput202 _125_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _124_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ repeater264/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l2_in_3_ mux_bottom_track_25.mux_l2_in_3_/A0 input21/X mux_bottom_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_ repeater247/X mux_bottom_track_17.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input46_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_7_ mux_right_track_4.mux_l2_in_7_/A0 _091_/A repeater227/X
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l1_in_2__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_25.mux_l2_in_3__295 VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_3_/A0
+ mux_bottom_track_25.mux_l2_in_3__295/LO sky130_fd_sc_hd__conb_1
XANTENNA_input100_A left_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ repeater259/X mux_top_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l2_in_3_ mux_bottom_track_9.mux_l2_in_3_/A0 _093_/A mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_25.mux_l4_in_0_ mux_bottom_track_25.mux_l3_in_1_/X mux_bottom_track_25.mux_l3_in_0_/X
+ mux_bottom_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _116_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 top_left_grid_pin_42_ VGND VGND VPWR VPWR input113/X sky130_fd_sc_hd__clkbuf_1
Xinput102 prog_clk_0_N_in VGND VGND VPWR VPWR input102/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l2_in_3__293 VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/A0
+ mux_bottom_track_1.mux_l2_in_3__293/LO sky130_fd_sc_hd__conb_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l3_in_1_ mux_bottom_track_25.mux_l2_in_3_/X mux_bottom_track_25.mux_l2_in_2_/X
+ mux_bottom_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l1_in_1_ input105/X _113_/A mux_right_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_1_ input119/X input117/X repeater226/X VGND VGND VPWR VPWR
+ mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input76_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput203 output203/A VGND VGND VPWR VPWR clk_1_E_out sky130_fd_sc_hd__buf_2
Xoutput214 output214/A VGND VGND VPWR VPWR prog_clk_1_W_out sky130_fd_sc_hd__buf_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ repeater262/X mux_bottom_track_5.mux_l5_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l2_in_2_ _095_/A _086_/A mux_bottom_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ repeater246/X mux_bottom_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__086__A _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_2_E_FTB01_A prog_clk_2_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_6_ _082_/A _131_/A repeater228/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l2_in_2_ input13/X _083_/A mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_2.mux_l1_in_4__A0 _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput114 top_left_grid_pin_43_ VGND VGND VPWR VPWR input114/X sky130_fd_sc_hd__clkbuf_1
Xinput103 prog_clk_1_N_in VGND VGND VPWR VPWR input103/X sky130_fd_sc_hd__clkbuf_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A0 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__094__A _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l1_in_0_ _103_/A input84/X mux_right_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ input115/X input113/X repeater226/X VGND VGND VPWR VPWR
+ mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input69_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput204 output204/A VGND VGND VPWR VPWR clk_1_W_out sky130_fd_sc_hd__buf_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput215 output215/A VGND VGND VPWR VPWR prog_clk_2_E_out sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_4.mux_l2_in_5__A1 _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclk_3_W_FTB01 input93/X VGND VGND VPWR VPWR output212/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_25.mux_l2_in_1_ input8/X mux_bottom_track_25.mux_l1_in_2_/X mux_bottom_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ repeater246/X mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xprog_clk_2_S_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR output217/A sky130_fd_sc_hd__buf_4
Xmux_right_track_4.mux_l2_in_5_ input68/X _122_/A repeater228/X VGND VGND VPWR VPWR
+ mux_right_track_4.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l2_in_3_ mux_top_track_16.mux_l2_in_3_/A0 _094_/A mux_top_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_2_ input4/X _075_/A mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_ repeater257/X mux_top_track_4.mux_l4_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l5_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l2_in_1_ input6/X mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input51_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_1
Xinput104 prog_clk_3_N_in VGND VGND VPWR VPWR input104/X sky130_fd_sc_hd__clkbuf_1
Xinput115 top_left_grid_pin_44_ VGND VGND VPWR VPWR input115/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_2.mux_l1_in_4__A1 _130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input99_A left_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A1 input44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l1_in_2_ input2/X _073_/A mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l4_in_0_ mux_top_track_16.mux_l3_in_1_/X mux_top_track_16.mux_l3_in_0_/X
+ mux_top_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input6_A bottom_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ repeater239/X mux_left_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_3_ mux_left_track_3.mux_l2_in_3_/A0 input101/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output218_A output218/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput205 output205/A VGND VGND VPWR VPWR clk_2_E_out sky130_fd_sc_hd__buf_2
Xoutput216 output216/A VGND VGND VPWR VPWR prog_clk_2_N_out sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l3_in_3_ mux_right_track_4.mux_l2_in_7_/X mux_right_track_4.mux_l2_in_6_/X
+ mux_right_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l3_in_1_ mux_top_track_16.mux_l2_in_3_/X mux_top_track_16.mux_l2_in_2_/X
+ mux_top_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input116_A top_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input81_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_7_ mux_bottom_track_5.mux_l2_in_7_/A0 _091_/A repeater236/X
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ repeater245/X mux_bottom_track_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_4_ input97/X input95/X repeater233/A VGND VGND VPWR VPWR
+ mux_left_track_3.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l2_in_4_ input112/X input111/X repeater228/A VGND VGND VPWR
+ VPWR mux_right_track_4.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l2_in_2_ _085_/A input28/X mux_top_track_16.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_1_ _066_/A input31/X mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_ repeater257/X mux_top_track_4.mux_l3_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l5_in_0_ mux_right_track_4.mux_l4_in_1_/X mux_right_track_4.mux_l4_in_0_/X
+ mux_right_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input44_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_1__A1 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput105 right_bottom_grid_pin_34_ VGND VGND VPWR VPWR input105/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput116 top_left_grid_pin_45_ VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 _065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_174 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l5_in_0_/X VGND VGND
+ VPWR VPWR _058_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_9.mux_l1_in_1_ _063_/A input44/X mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l4_in_1_ mux_right_track_4.mux_l3_in_3_/X mux_right_track_4.mux_l3_in_2_/X
+ mux_right_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_7__284 VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_7_/A0
+ mux_right_track_4.mux_l2_in_7__284/LO sky130_fd_sc_hd__conb_1
XFILLER_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ repeater239/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_2_ input99/X mux_left_track_3.mux_l1_in_4_/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput206 output206/A VGND VGND VPWR VPWR clk_2_N_out sky130_fd_sc_hd__buf_2
Xoutput217 output217/A VGND VGND VPWR VPWR prog_clk_2_S_out sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l3_in_2_ mux_right_track_4.mux_l2_in_5_/X mux_right_track_4.mux_l2_in_4_/X
+ mux_right_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input109_A right_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input74_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_6_ input28/X _082_/A repeater236/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_ repeater273/X mux_right_track_4.mux_l4_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l5_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_3_ _130_/A _121_/A repeater233/X VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A0 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_3_ mux_right_track_16.mux_l2_in_3_/A0 _094_/A mux_right_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_3_ input110/X input109/X repeater227/X VGND VGND VPWR
+ VPWR mux_right_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_16.mux_l2_in_1_ _134_/A mux_top_track_16.mux_l1_in_2_/X mux_top_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_0_ _115_/A _106_/A mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ repeater256/X repeater224/A VGND VGND
+ VPWR VPWR mux_top_track_4.mux_l3_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input37_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_4__A0 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 _065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput106 right_bottom_grid_pin_35_ VGND VGND VPWR VPWR input106/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput117 top_left_grid_pin_46_ VGND VGND VPWR VPWR input117/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_ _125_/A _074_/A mux_top_track_16.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_25.mux_l2_in_3__302 VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_3_/A0
+ mux_left_track_25.mux_l2_in_3__302/LO sky130_fd_sc_hd__conb_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l4_in_0_ mux_right_track_16.mux_l3_in_1_/X mux_right_track_16.mux_l3_in_0_/X
+ mux_right_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l1_in_0_ _113_/A _103_/A mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l1_in_1__A1 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_25.mux_l2_in_2__A0 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ repeater242/X repeater234/X VGND VGND
+ VPWR VPWR mux_left_track_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l3_in_1_ mux_right_track_16.mux_l2_in_3_/X mux_right_track_16.mux_l2_in_2_/X
+ mux_right_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput207 output207/A VGND VGND VPWR VPWR clk_2_S_out sky130_fd_sc_hd__buf_2
Xoutput218 output218/A VGND VGND VPWR VPWR prog_clk_2_W_out sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_2__A1 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input67_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_5_ input9/X input8/X repeater235/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ repeater271/X mux_right_track_4.mux_l3_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_2_ input51/X _070_/A repeater233/X VGND VGND VPWR VPWR
+ mux_left_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_2_ _085_/A _134_/A mux_right_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_4.mux_l2_in_2_ input108/X input107/X repeater227/X VGND VGND VPWR
+ VPWR mux_right_track_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A0 _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ repeater256/X mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR repeater224/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_4__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput107 right_bottom_grid_pin_36_ VGND VGND VPWR VPWR input107/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput118 top_left_grid_pin_47_ VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l1_in_1_ input37/X _065_/A mux_top_track_16.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input97_A left_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l2_in_3__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_3_ mux_bottom_track_5.mux_l2_in_7_/X mux_bottom_track_5.mux_l2_in_6_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_25.mux_l2_in_2__A1 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ repeater263/X mux_bottom_track_33.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR repeater234/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput208 output208/A VGND VGND VPWR VPWR clk_2_W_out sky130_fd_sc_hd__buf_2
Xoutput219 output219/A VGND VGND VPWR VPWR prog_clk_3_E_out sky130_fd_sc_hd__buf_2
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input4_A bottom_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A0 _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_4_ input7/X input6/X repeater236/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ repeater271/X repeater228/X VGND VGND
+ VPWR VPWR mux_right_track_4.mux_l3_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l1_in_1_ _061_/A input81/X repeater233/X VGND VGND VPWR VPWR
+ mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_7__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_16.mux_l2_in_1_ _125_/A mux_right_track_16.mux_l1_in_2_/X mux_right_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input114_A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l5_in_0_ mux_bottom_track_5.mux_l4_in_1_/X mux_bottom_track_5.mux_l4_in_0_/X
+ mux_bottom_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_2__A1 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ input106/X input105/X repeater227/X VGND VGND VPWR
+ VPWR mux_right_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_1_W_FTB01 input103/X VGND VGND VPWR VPWR output214/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ repeater256/X mux_top_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_33.mux_l1_in_3__A1 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_0.mux_l1_in_3__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_2_ input62/X input110/X mux_right_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xinput108 right_bottom_grid_pin_37_ VGND VGND VPWR VPWR input108/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l4_in_1_ mux_bottom_track_5.mux_l3_in_3_/X mux_bottom_track_5.mux_l3_in_2_/X
+ mux_bottom_track_5.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput119 top_left_grid_pin_48_ VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ input118/X input114/X mux_top_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_24.mux_l2_in_3__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput90 chany_top_in[9] VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_right_track_0.mux_l2_in_2__A0 _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_3__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l3_in_2_ mux_bottom_track_5.mux_l2_in_5_/X mux_bottom_track_5.mux_l2_in_4_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput209 output209/A VGND VGND VPWR VPWR clk_3_E_out sky130_fd_sc_hd__buf_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_33.mux_l1_in_1__A1 _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_3_ input5/X input4/X repeater235/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ repeater271/X mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR repeater228/A sky130_fd_sc_hd__dfxtp_1
Xclk_3_S_FTB01 input93/X VGND VGND VPWR VPWR output211/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_3.mux_l1_in_0_ _110_/A _101_/A repeater233/X VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ _111_/A mux_right_track_4.mux_l1_in_0_/X repeater228/X
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input107_A right_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input72_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2__A0 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_16.mux_l2_in_3__287 VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_3_/A0
+ mux_top_track_16.mux_l2_in_3__287/LO sky130_fd_sc_hd__conb_1
XANTENNA__122__A _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclk_1_E_FTB01 input91/X VGND VGND VPWR VPWR output203/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_1_ input106/X _114_/A mux_right_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput109 right_bottom_grid_pin_38_ VGND VGND VPWR VPWR input109/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_3__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input35_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_129_ _129_/A VGND VGND VPWR VPWR _129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput80 chany_top_in[18] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__clkbuf_2
Xinput91 clk_1_N_in VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_3__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__130__A _130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_2_ input3/X input2/X repeater235/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_ repeater243/X mux_bottom_track_5.mux_l4_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l5_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ repeater269/X mux_right_track_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_3__278 VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/A0
+ mux_left_track_9.mux_l2_in_3__278/LO sky130_fd_sc_hd__conb_1
XANTENNA_input65_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
Xinput1 Test_en_S_in VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_2__A1 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l1_in_0_ _105_/A input88/X mux_right_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ _102_/A input82/X mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l5_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
Xoutput190 _132_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xprog_clk_2_N_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR output216/A sky130_fd_sc_hd__buf_4
XANTENNA__133__A _133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_128_ _128_/A VGND VGND VPWR VPWR _128_/X sky130_fd_sc_hd__clkbuf_1
X_059_ _059_/A VGND VGND VPWR VPWR _059_/X sky130_fd_sc_hd__clkbuf_1
Xinput81 chany_top_in[19] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput70 chany_bottom_in[9] VGND VGND VPWR VPWR _126_/A sky130_fd_sc_hd__clkbuf_2
Xinput92 clk_2_N_in VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input95_A left_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l1_in_4__A0 _130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_1_ _071_/A input48/X repeater236/A VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_ repeater242/X mux_bottom_track_5.mux_l3_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input2_A bottom_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
Xinput2 bottom_left_grid_pin_42_ VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_33.mux_l1_in_3_ mux_bottom_track_33.mux_l1_in_3_/A0 _087_/A mux_bottom_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input112_A right_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput191 _133_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput180 _103_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_058_ _058_/A VGND VGND VPWR VPWR _058_/X sky130_fd_sc_hd__clkbuf_1
X_127_ _127_/A VGND VGND VPWR VPWR _127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput71 chany_top_in[0] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 chany_bottom_in[18] VGND VGND VPWR VPWR _135_/A sky130_fd_sc_hd__buf_2
Xinput82 chany_top_in[1] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_1
Xinput93 clk_3_N_in VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input40_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 _059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input88_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_0_ _062_/A mux_bottom_track_5.mux_l1_in_0_/X repeater236/A
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l2_in_1_ mux_bottom_track_33.mux_l1_in_3_/X mux_bottom_track_33.mux_l1_in_2_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ repeater242/X repeater235/X VGND VGND
+ VPWR VPWR mux_bottom_track_5.mux_l3_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _056_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_16.mux_l2_in_3__280 VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_3_/A0
+ mux_right_track_16.mux_l2_in_3__280/LO sky130_fd_sc_hd__conb_1
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 bottom_left_grid_pin_43_ VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_2.mux_l2_in_3__A1 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_3_ mux_top_track_24.mux_l2_in_3_/A0 _095_/A mux_top_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__062__A _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.mux_l1_in_2_ input11/X input9/X mux_bottom_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input105_A right_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input70_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_3_ mux_left_track_17.mux_l2_in_3_/A0 input99/X mux_left_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput192 _134_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
Xoutput181 _104_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xoutput170 _112_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ _057_/A VGND VGND VPWR VPWR _057_/X sky130_fd_sc_hd__clkbuf_1
X_126_ _126_/A VGND VGND VPWR VPWR _126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput72 chany_top_in[10] VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_2
Xinput61 chany_bottom_in[19] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
Xinput50 chanx_right_in[9] VGND VGND VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_2
Xinput94 left_bottom_grid_pin_34_ VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__clkbuf_1
Xinput83 chany_top_in[2] VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A0 _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input33_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l4_in_0_ mux_top_track_24.mux_l3_in_1_/X mux_top_track_24.mux_l3_in_0_/X
+ mux_top_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l2_in_3_ mux_left_track_9.mux_l2_in_3_/A0 input98/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_3_E_FTB01 input104/X VGND VGND VPWR VPWR output219/A sky130_fd_sc_hd__clkbuf_1
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.mux_l2_in_3_ mux_right_track_0.mux_l2_in_3_/A0 _089_/A mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.mux_l4_in_0_ mux_left_track_17.mux_l3_in_1_/X mux_left_track_17.mux_l3_in_0_/X
+ mux_left_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__065__A _065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l3_in_1_ mux_top_track_24.mux_l2_in_3_/X mux_top_track_24.mux_l2_in_2_/X
+ mux_top_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ repeater244/X mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR repeater236/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclk_2_W_FTB01 input92/X VGND VGND VPWR VPWR output208/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_0.mux_l1_in_4_ input57/X _129_/A repeater230/A VGND VGND VPWR VPWR
+ mux_right_track_0.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.mux_l3_in_1_ mux_left_track_17.mux_l2_in_3_/X mux_left_track_17.mux_l2_in_2_/X
+ mux_left_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l5_in_0_/X VGND
+ VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xinput4 bottom_left_grid_pin_44_ VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_2_ _086_/A input24/X mux_top_track_24.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ _111_/A _102_/A mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_1_ input5/X input41/X mux_bottom_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input63_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l2_in_2_ input95/X _134_/A mux_left_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__073__A _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput193 _135_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xmux_left_track_3.mux_l2_in_3__303 VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/A0
+ mux_left_track_3.mux_l2_in_3__303/LO sky130_fd_sc_hd__conb_1
Xoutput182 _105_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xoutput171 _113_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput160 _083_/X VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
X_125_ _125_/A VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__clkbuf_1
X_056_ _056_/A VGND VGND VPWR VPWR _056_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput73 chany_top_in[11] VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_bottom_in[0] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 chany_bottom_in[1] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
Xinput95 left_bottom_grid_pin_35_ VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput40 chanx_right_in[18] VGND VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_2
Xinput84 chany_top_in[3] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input26_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_2_ input94/X _133_/A mux_left_track_9.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_2_ _079_/A mux_right_track_0.mux_l1_in_4_/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__081__A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ repeater244/X mux_bottom_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input93_A clk_3_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_3_ _119_/A input111/X repeater230/X VGND VGND VPWR VPWR
+ mux_right_track_0.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_3_ mux_top_track_2.mux_l2_in_3_/A0 input21/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_3_ mux_right_track_24.mux_l2_in_3_/A0 _095_/A mux_right_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xinput5 bottom_left_grid_pin_45_ VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_8.mux_l1_in_1__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_1_ _135_/A mux_top_track_24.mux_l1_in_2_/X mux_top_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_0_ _067_/A _107_/A mux_bottom_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input56_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l2_in_1_ _125_/A mux_left_track_17.mux_l1_in_2_/X mux_left_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_4_ _081_/A _130_/A repeater225/X VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_4_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput161 _084_/X VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l1_in_3__A0 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput150 _092_/X VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xoutput183 _116_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput172 _114_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xoutput194 _117_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_input110_A right_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ _124_/A VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_2_ _126_/A input41/X mux_top_track_24.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput74 chany_top_in[12] VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_2
Xinput85 chany_top_in[4] VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_2
Xinput96 left_bottom_grid_pin_36_ VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__clkbuf_1
Xinput63 chany_bottom_in[2] VGND VGND VPWR VPWR _119_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 chany_bottom_in[10] VGND VGND VPWR VPWR _127_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 chanx_left_in[9] VGND VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_2
Xinput41 chanx_right_in[19] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmux_right_track_24.mux_l4_in_0_ mux_right_track_24.mux_l3_in_1_/X mux_right_track_24.mux_l3_in_0_/X
+ mux_right_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l2_in_7__277 VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_7_/A0
+ mux_left_track_5.mux_l2_in_7__277/LO sky130_fd_sc_hd__conb_1
XANTENNA_input19_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_2_ input68/X _074_/A mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A0 _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_1_ _123_/A mux_left_track_9.mux_l1_in_2_/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__079__A _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_1_ mux_right_track_0.mux_l1_in_3_/X mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_1_ mux_right_track_24.mux_l2_in_3_/X mux_right_track_24.mux_l2_in_2_/X
+ mux_right_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input86_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_2_ input64/X _073_/A mux_left_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_2_ input109/X input107/X repeater230/X VGND VGND VPWR
+ VPWR mux_right_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_2_ _090_/A mux_top_track_2.mux_l1_in_4_/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_2_ _086_/A _135_/A mux_right_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xinput6 bottom_left_grid_pin_46_ VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 _061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_3_ _121_/A _070_/A repeater225/X VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xclk_3_N_FTB01 input93/X VGND VGND VPWR VPWR output210/A sky130_fd_sc_hd__clkbuf_1
Xoutput184 _126_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput195 _118_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_7_ mux_left_track_5.mux_l2_in_7_/A0 input101/X repeater231/X
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
Xoutput173 _115_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xoutput140 _063_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput162 _085_/X VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_2.mux_l1_in_3__A1 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput151 _093_/X VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XANTENNA_input103_A prog_clk_1_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_123_ _123_/A VGND VGND VPWR VPWR _123_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_1_ _075_/A _066_/A mux_top_track_24.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput31 chanx_right_in[0] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[18] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_2
Xinput75 chany_top_in[13] VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_2
Xinput86 chany_top_in[5] VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput97 left_bottom_grid_pin_37_ VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_1
Xinput42 chanx_right_in[1] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 chany_bottom_in[3] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_bottom_in[11] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_3__290 VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_3_/A0
+ mux_top_track_32.mux_l1_in_3__290/LO sky130_fd_sc_hd__conb_1
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l2_in_3_ mux_bottom_track_1.mux_l2_in_3_/A0 _089_/A mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_1_ _065_/A _114_/A mux_left_track_17.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input31_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xrepeater270 repeater272/X VGND VGND VPWR VPWR repeater270/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l1_in_4_ input22/X input8/X repeater238/X VGND VGND VPWR VPWR
+ mux_bottom_track_1.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_1_ _063_/A _113_/A mux_left_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input79_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_1_ input105/X input81/X repeater230/X VGND VGND VPWR
+ VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ _126_/A mux_right_track_24.mux_l1_in_2_/X mux_right_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 bottom_left_grid_pin_47_ VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__A1 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ repeater255/X mux_top_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _128_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l1_in_2_ _061_/A input44/X repeater225/X VGND VGND VPWR VPWR
+ mux_top_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l2_in_3__299 VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/A0
+ mux_bottom_track_9.mux_l2_in_3__299/LO sky130_fd_sc_hd__conb_1
Xmux_right_track_24.mux_l1_in_2_ input51/X input111/X mux_right_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput185 _127_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xoutput196 _119_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xoutput152 _094_/X VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_1.mux_l1_in_3__A1 _129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput163 _096_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput174 _097_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_6_ input100/X input99/X repeater231/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
Xoutput141 _064_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput130 _072_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_17.mux_l2_in_3__294 VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_3_/A0
+ mux_bottom_track_17.mux_l2_in_3__294/LO sky130_fd_sc_hd__conb_1
XANTENNA_input61_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_122_ _122_/A VGND VGND VPWR VPWR _122_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_0_ input119/X input115/X mux_top_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ repeater265/X mux_right_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xinput10 ccff_head VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
Xinput43 chanx_right_in[2] VGND VGND VPWR VPWR _059_/A sky130_fd_sc_hd__clkbuf_2
Xinput54 chany_bottom_in[12] VGND VGND VPWR VPWR _129_/A sky130_fd_sc_hd__clkbuf_2
Xinput32 chanx_right_in[10] VGND VGND VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[19] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 chany_top_in[14] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput65 chany_bottom_in[4] VGND VGND VPWR VPWR _121_/A sky130_fd_sc_hd__clkbuf_2
Xinput98 left_bottom_grid_pin_38_ VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_1
Xinput87 chany_top_in[6] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_33.mux_l1_in_3__276 VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_3_/A0
+ mux_left_track_33.mux_l1_in_3__276/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_2_ _079_/A mux_bottom_track_1.mux_l1_in_4_/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_0_ _105_/A input88/X mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l1_in_3_ input6/X input4/X repeater238/X VGND VGND VPWR VPWR
+ mux_bottom_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xrepeater271 repeater272/X VGND VGND VPWR VPWR repeater271/X sky130_fd_sc_hd__clkbuf_1
Xrepeater260 repeater261/X VGND VGND VPWR VPWR repeater260/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l1_in_0_ input73/X _103_/A mux_left_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_0_ _109_/A _099_/A repeater230/X VGND VGND VPWR VPWR
+ mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _117_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input91_A clk_1_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 bottom_left_grid_pin_48_ VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ repeater240/X mux_left_track_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ repeater255/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_prog_clk_2_W_FTB01_A prog_clk_2_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_8.mux_l2_in_3__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l2_in_3__A0 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_1_ input120/X input118/X repeater225/X VGND VGND VPWR VPWR
+ mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_1_ input107/X _115_/A mux_right_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput153 _095_/X VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
Xoutput186 _128_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput197 _120_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput175 _098_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput164 _106_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_5_ input98/X input97/X repeater231/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
Xoutput142 _065_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput131 _073_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xmux_left_track_1.mux_l2_in_3__300 VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/A0
+ mux_left_track_1.mux_l2_in_3__300/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A0 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ _121_/A VGND VGND VPWR VPWR _121_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input54_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ repeater266/X mux_right_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xinput77 chany_top_in[15] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 chanx_left_in[1] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput44 chanx_right_in[3] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput66 chany_bottom_in[5] VGND VGND VPWR VPWR _122_/A sky130_fd_sc_hd__clkbuf_2
Xinput55 chany_bottom_in[13] VGND VGND VPWR VPWR _130_/A sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[0] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput33 chanx_right_in[11] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput88 chany_top_in[7] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__clkbuf_1
Xinput99 left_bottom_grid_pin_39_ VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A1 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_16.mux_l2_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_7__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input17_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l1_in_2_ input2/X input37/X repeater238/X VGND VGND VPWR VPWR
+ mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xrepeater250 repeater251/X VGND VGND VPWR VPWR repeater250/X sky130_fd_sc_hd__clkbuf_1
Xrepeater272 repeater273/X VGND VGND VPWR VPWR repeater272/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input9_A bottom_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater261 repeater268/X VGND VGND VPWR VPWR repeater261/X sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ repeater270/X mux_right_track_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_5.mux_l2_in_6__A0 input28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_3__281 VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/A0
+ mux_right_track_2.mux_l2_in_3__281/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l3_in_3_ mux_left_track_5.mux_l2_in_7_/X mux_left_track_5.mux_l2_in_6_/X
+ mux_left_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input119_A top_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input84_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_2_S_FTB01_A prog_clk_2_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 bottom_left_grid_pin_49_ VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ repeater239/X mux_left_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclk_2_S_FTB01 input92/X VGND VGND VPWR VPWR output207/A sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ repeater248/X repeater226/X VGND VGND
+ VPWR VPWR mux_top_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l1_in_0_ input116/X input114/X repeater225/A VGND VGND VPWR VPWR
+ mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_0_ input73/X _106_/A mux_right_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput121 output121/A VGND VGND VPWR VPWR Test_en_N_out sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_4_ input96/X input95/X repeater231/X VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
Xoutput143 _076_/X VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xoutput132 _074_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xoutput187 _129_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput198 _121_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput176 _099_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xoutput165 _107_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput154 _077_/X VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A1 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_120_ _120_/A VGND VGND VPWR VPWR _120_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input47_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ repeater272/X mux_right_track_24.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_24.mux_l2_in_2__A0 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput89 chany_top_in[8] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_2
Xinput45 chanx_right_in[4] VGND VGND VPWR VPWR _061_/A sky130_fd_sc_hd__clkbuf_2
Xinput67 chany_bottom_in[6] VGND VGND VPWR VPWR _123_/A sky130_fd_sc_hd__clkbuf_2
Xinput56 chany_bottom_in[14] VGND VGND VPWR VPWR _131_/A sky130_fd_sc_hd__buf_2
Xinput23 chanx_left_in[2] VGND VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[10] VGND VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_2
Xinput34 chanx_right_in[12] VGND VGND VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_2
Xinput78 chany_top_in[16] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__clkbuf_2
Xmux_left_track_5.mux_l5_in_0_ mux_left_track_5.mux_l4_in_1_/X mux_left_track_5.mux_l4_in_0_/X
+ mux_left_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ repeater251/X mux_left_track_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input101_A left_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_2__A0 _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A1 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l2_in_3__288 VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/A0
+ mux_top_track_2.mux_l2_in_3__288/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_16.mux_l2_in_2__A1 _134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l4_in_1_ mux_left_track_5.mux_l3_in_3_/X mux_left_track_5.mux_l3_in_2_/X
+ mux_left_track_5.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xrepeater262 repeater263/X VGND VGND VPWR VPWR repeater262/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l1_in_1_ _069_/A _059_/A repeater238/A VGND VGND VPWR VPWR
+ mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xrepeater240 repeater241/X VGND VGND VPWR VPWR repeater240/X sky130_fd_sc_hd__clkbuf_1
Xrepeater251 repeater252/X VGND VGND VPWR VPWR repeater251/X sky130_fd_sc_hd__clkbuf_1
Xrepeater273 repeater274/X VGND VGND VPWR VPWR repeater273/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ repeater270/X mux_right_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_5.mux_l2_in_6__A1 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_2_ mux_left_track_5.mux_l2_in_5_/X mux_left_track_5.mux_l2_in_4_/X
+ mux_left_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 _062_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input77_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ repeater241/X repeater233/A VGND VGND
+ VPWR VPWR mux_left_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ repeater242/X input10/X VGND VGND VPWR
+ VPWR repeater226/A sky130_fd_sc_hd__dfxtp_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput122 output122/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
Xoutput177 _100_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xoutput166 _108_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_3_ input94/X _131_/A repeater232/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xoutput155 _078_/X VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
Xoutput144 _086_/X VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xoutput133 _075_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xoutput188 _130_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xoutput199 _122_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_24.mux_l2_in_2__A0 _086_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput13 chanx_left_in[11] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_24.mux_l2_in_2__A1 _135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput46 chanx_right_in[5] VGND VGND VPWR VPWR _062_/A sky130_fd_sc_hd__clkbuf_2
Xinput57 chany_bottom_in[15] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_bottom_in[7] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_1
Xinput24 chanx_left_in[3] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chanx_right_in[13] VGND VGND VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_2
Xinput79 chany_top_in[17] VGND VGND VPWR VPWR _114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ repeater251/X mux_left_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_16.mux_l2_in_2__A1 input28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l1_in_0_ _109_/A _099_/A repeater238/A VGND VGND VPWR VPWR
+ mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xrepeater230 repeater230/A VGND VGND VPWR VPWR repeater230/X sky130_fd_sc_hd__clkbuf_2
Xrepeater241 repeater245/X VGND VGND VPWR VPWR repeater241/X sky130_fd_sc_hd__clkbuf_1
Xrepeater263 repeater264/X VGND VGND VPWR VPWR repeater263/X sky130_fd_sc_hd__clkbuf_1
Xrepeater252 repeater253/X VGND VGND VPWR VPWR repeater252/X sky130_fd_sc_hd__clkbuf_1
Xrepeater274 repeater275/X VGND VGND VPWR VPWR repeater274/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input22_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.mux_l1_in_3__A1 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ repeater270/X repeater230/A VGND VGND
+ VPWR VPWR mux_right_track_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ repeater239/X mux_left_track_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater233/A sky130_fd_sc_hd__dfxtp_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l2_in_6__A0 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1__A0 _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput189 _131_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput178 _101_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput167 _109_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_2_ _122_/A input62/X repeater232/A VGND VGND VPWR VPWR
+ mux_left_track_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput123 _056_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xoutput134 _057_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_ repeater273/X mux_right_track_24.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xoutput156 _079_/X VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
Xoutput145 _087_/X VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_3_ mux_left_track_25.mux_l2_in_3_/A0 input100/X mux_left_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_2__A1 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput25 chanx_left_in[4] VGND VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_2
Xinput14 chanx_left_in[12] VGND VGND VPWR VPWR _089_/A sky130_fd_sc_hd__buf_2
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput36 chanx_right_in[14] VGND VGND VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_2
Xinput47 chanx_right_in[6] VGND VGND VPWR VPWR _063_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 chany_bottom_in[8] VGND VGND VPWR VPWR _125_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 chany_bottom_in[16] VGND VGND VPWR VPWR _133_/A sky130_fd_sc_hd__clkbuf_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ repeater251/X mux_left_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input52_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_3__301 VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_3_/A0
+ mux_left_track_17.mux_l2_in_3__301/LO sky130_fd_sc_hd__conb_1
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l2_in_2__A1 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l4_in_0_ mux_left_track_25.mux_l3_in_1_/X mux_left_track_25.mux_l3_in_0_/X
+ mux_left_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xrepeater242 repeater243/X VGND VGND VPWR VPWR repeater242/X sky130_fd_sc_hd__clkbuf_1
Xrepeater231 repeater232/X VGND VGND VPWR VPWR repeater231/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater253 repeater254/X VGND VGND VPWR VPWR repeater253/X sky130_fd_sc_hd__clkbuf_1
Xrepeater264 repeater265/X VGND VGND VPWR VPWR repeater264/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater275 repeater275/A VGND VGND VPWR VPWR repeater275/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_32.mux_l1_in_3__A1 _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _064_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l2_in_7__298 VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_7_/A0
+ mux_bottom_track_5.mux_l2_in_7__298/LO sky130_fd_sc_hd__conb_1
XANTENNA_input15_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ repeater268/X mux_top_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR repeater230/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A bottom_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l3_in_1_ mux_left_track_25.mux_l2_in_3_/X mux_left_track_25.mux_l2_in_2_/X
+ mux_left_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l2_in_6__A1 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input117_A top_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_1_ _071_/A _062_/A repeater232/X VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput179 _102_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput168 _110_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput135 _058_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ repeater274/X mux_right_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xoutput157 _080_/X VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
Xoutput124 _066_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xoutput146 _088_/X VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_2_ input96/X _135_/A mux_left_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 chanx_left_in[5] VGND VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_2
Xinput59 chany_bottom_in[17] VGND VGND VPWR VPWR _134_/A sky130_fd_sc_hd__clkbuf_2
Xinput48 chanx_right_in[7] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 chanx_left_in[13] VGND VGND VPWR VPWR _090_/A sky130_fd_sc_hd__buf_2
Xinput37 chanx_right_in[15] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mux_left_track_17.mux_l2_in_2__A1 _134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_3_ mux_top_track_32.mux_l1_in_3_/A0 _087_/A mux_top_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ repeater250/X mux_left_track_5.mux_l5_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input45_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 _059_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ repeater241/X mux_left_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR output122/A sky130_fd_sc_hd__dfxtp_1
Xrepeater243 repeater244/X VGND VGND VPWR VPWR repeater243/X sky130_fd_sc_hd__clkbuf_1
Xrepeater232 repeater232/A VGND VGND VPWR VPWR repeater232/X sky130_fd_sc_hd__clkbuf_1
Xrepeater265 repeater266/X VGND VGND VPWR VPWR repeater265/X sky130_fd_sc_hd__clkbuf_1
Xrepeater254 repeater259/X VGND VGND VPWR VPWR repeater254/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xprog_clk_2_E_FTB01 prog_clk_2_N_in VGND VGND VPWR VPWR output215/A sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_2.mux_l1_in_3__A0 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_ repeater262/X mux_bottom_track_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__131__A _131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_3_ mux_top_track_8.mux_l2_in_3_/A0 _093_/A mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__126__A _126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l2_in_1_ mux_top_track_32.mux_l1_in_3_/X mux_top_track_32.mux_l1_in_2_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_2__A0 _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclk_1_W_FTB01 input91/X VGND VGND VPWR VPWR output204/A sky130_fd_sc_hd__clkbuf_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_25.mux_l2_in_2__A1 _135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input75_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l2_in_0_ input77/X mux_left_track_5.mux_l1_in_0_/X repeater232/A
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ repeater274/X mux_right_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xoutput125 _067_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xoutput169 _111_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput136 _059_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xoutput158 _081_/X VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xoutput147 _089_/X VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_1_ input53/X mux_left_track_25.mux_l1_in_2_/X mux_left_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 chanx_left_in[6] VGND VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_2
Xinput49 chanx_right_in[8] VGND VGND VPWR VPWR _065_/A sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[14] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_2
Xinput38 chanx_right_in[16] VGND VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_32.mux_l1_in_2_ input22/X _127_/A mux_top_track_32.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input38_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_25.mux_l1_in_2_ _126_/A _075_/A mux_left_track_25.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__134__A _134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ repeater240/X mux_left_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__129__A _129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater233 repeater233/A VGND VGND VPWR VPWR repeater233/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater244 repeater245/X VGND VGND VPWR VPWR repeater244/X sky130_fd_sc_hd__clkbuf_1
Xrepeater266 repeater267/X VGND VGND VPWR VPWR repeater266/X sky130_fd_sc_hd__clkbuf_1
Xrepeater255 repeater256/X VGND VGND VPWR VPWR repeater255/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ repeater262/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_2_ input13/X _083_/A mux_top_track_8.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input68_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput137 _060_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ repeater275/A mux_right_track_16.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xoutput159 _082_/X VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xoutput126 _068_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xoutput148 _090_/X VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.mux_l1_in_3_ mux_right_track_32.mux_l1_in_3_/A0 _087_/A mux_right_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 chanx_left_in[7] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_left_in[15] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput39 chanx_right_in[17] VGND VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_32.mux_l1_in_1_ _067_/A input31/X mux_top_track_32.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l1_in_0_ _111_/A _102_/A mux_left_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l1_in_1_ _066_/A _115_/A mux_left_track_25.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l2_in_3__286 VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/A0
+ mux_top_track_0.mux_l2_in_3__286/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ repeater249/X mux_left_track_25.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input50_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xrepeater256 repeater257/X VGND VGND VPWR VPWR repeater256/X sky130_fd_sc_hd__clkbuf_1
Xrepeater234 repeater234/A VGND VGND VPWR VPWR repeater234/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater245 repeater246/X VGND VGND VPWR VPWR repeater245/X sky130_fd_sc_hd__clkbuf_1
Xrepeater267 repeater268/X VGND VGND VPWR VPWR repeater267/X sky130_fd_sc_hd__clkbuf_1
Xrepeater223 repeater224/X VGND VGND VPWR VPWR repeater223/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input98_A left_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ repeater263/X repeater238/X VGND VGND
+ VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_1_ _133_/A mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_1_ mux_right_track_32.mux_l1_in_3_/X mux_right_track_32.mux_l1_in_2_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input13_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input5_A bottom_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_2_ _123_/A _073_/A mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l1_in_2__A1 _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput138 _061_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput127 _069_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xoutput149 _091_/X VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xmux_right_track_32.mux_l1_in_2_ input61/X _127_/A mux_right_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__063__A _063_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A top_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[16] VGND VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input80_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 chanx_left_in[8] VGND VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_2
Xmux_top_track_32.mux_l1_in_0_ input120/X input116/X mux_top_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclk_2_N_FTB01 input92/X VGND VGND VPWR VPWR output206/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l1_in_0_ _106_/A input84/X mux_left_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l2_in_7_ mux_top_track_4.mux_l2_in_7_/A0 input17/X repeater223/X
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater235 repeater236/X VGND VGND VPWR VPWR repeater235/X sky130_fd_sc_hd__dlymetal6s2s_1
Xrepeater224 repeater224/A VGND VGND VPWR VPWR repeater224/X sky130_fd_sc_hd__clkbuf_2
Xrepeater246 repeater247/X VGND VGND VPWR VPWR repeater246/X sky130_fd_sc_hd__clkbuf_1
Xrepeater268 repeater275/X VGND VGND VPWR VPWR repeater268/X sky130_fd_sc_hd__clkbuf_1
Xrepeater257 repeater258/X VGND VGND VPWR VPWR repeater257/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ repeater269/X mux_right_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR repeater238/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__066__A _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_ repeater275/X mux_right_track_16.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ input33/X _063_/A mux_top_track_8.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _120_/A sky130_fd_sc_hd__clkbuf_1
Xoutput139 _062_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput128 _070_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xmux_right_track_32.mux_l1_in_1_ input112/X input108/X mux_right_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_2.mux_l1_in_2__A0 _061_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input108_A right_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput19 chanx_left_in[17] VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input73_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
Xprog_clk_3_W_FTB01 input104/X VGND VGND VPWR VPWR output222/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_ repeater249/X mux_left_track_25.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_6_ _091_/A _082_/A repeater223/X VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_6_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__069__A _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input36_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
Xrepeater236 repeater236/A VGND VGND VPWR VPWR repeater236/X sky130_fd_sc_hd__clkbuf_2
Xrepeater269 repeater271/X VGND VGND VPWR VPWR repeater269/X sky130_fd_sc_hd__clkbuf_1
Xrepeater247 repeater261/X VGND VGND VPWR VPWR repeater247/X sky130_fd_sc_hd__clkbuf_1
Xrepeater225 repeater225/A VGND VGND VPWR VPWR repeater225/X sky130_fd_sc_hd__clkbuf_2
Xrepeater258 repeater260/X VGND VGND VPWR VPWR repeater258/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_1.mux_l2_in_3_ mux_left_track_1.mux_l2_in_3_/A0 input100/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ repeater275/X mux_right_track_16.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ input117/X input113/X mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l1_in_4_ input96/X input94/X repeater234/X VGND VGND VPWR VPWR
+ mux_left_track_1.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xoutput129 _071_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xmux_right_track_32.mux_l1_in_0_ input77/X _107_/A mux_right_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_2__A1 input44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ repeater261/X mux_top_track_32.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input66_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__090__A _090_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_4__A1 _129_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input120_A top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_3__292 VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/A0
+ mux_top_track_8.mux_l2_in_3__292/LO sky130_fd_sc_hd__conb_1
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ repeater249/X mux_left_track_25.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _057_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l2_in_5_ _131_/A _122_/A repeater224/X VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_5_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input29_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater237 repeater237/A VGND VGND VPWR VPWR repeater237/X sky130_fd_sc_hd__clkbuf_2
Xrepeater226 repeater226/A VGND VGND VPWR VPWR repeater226/X sky130_fd_sc_hd__clkbuf_2
Xrepeater248 repeater252/X VGND VGND VPWR VPWR repeater248/X sky130_fd_sc_hd__clkbuf_1
Xrepeater259 repeater260/X VGND VGND VPWR VPWR repeater259/X sky130_fd_sc_hd__clkbuf_1
Xclk_3_E_FTB01 input93/X VGND VGND VPWR VPWR output209/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_2_ input98/X mux_left_track_1.mux_l1_in_4_/X mux_left_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input96_A left_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ repeater268/X mux_right_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input11_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_2__A0 _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_3_ input61/X _129_/A repeater234/A VGND VGND VPWR VPWR
+ mux_left_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_2.mux_l2_in_3_ mux_right_track_2.mux_l2_in_3_/A0 _090_/A mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A bottom_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ repeater261/X mux_top_track_32.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_3_ mux_top_track_4.mux_l2_in_7_/X mux_top_track_4.mux_l2_in_6_/X
+ mux_top_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input59_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input113_A top_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 _065_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ repeater246/X mux_left_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l1_in_4_ _130_/A input53/X repeater229/X VGND VGND VPWR VPWR
+ mux_right_track_2.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_4_ _071_/A input48/X repeater223/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_6__A0 _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l5_in_0_ mux_top_track_4.mux_l4_in_1_/X mux_top_track_4.mux_l4_in_0_/X
+ mux_top_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xrepeater238 repeater238/A VGND VGND VPWR VPWR repeater238/X sky130_fd_sc_hd__clkbuf_2
Xrepeater227 repeater228/A VGND VGND VPWR VPWR repeater227/X sky130_fd_sc_hd__clkbuf_2
Xrepeater249 repeater250/X VGND VGND VPWR VPWR repeater249/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input41_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l4_in_1_ mux_top_track_4.mux_l3_in_3_/X mux_top_track_4.mux_l3_in_2_/X
+ mux_top_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input89_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_2_N_FTB01_A prog_clk_2_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ repeater267/X mux_right_track_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_8.mux_l2_in_2__A1 _133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l1_in_2_ _119_/A _069_/A repeater234/X VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_2_ _081_/A mux_right_track_2.mux_l1_in_4_/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_2_ mux_top_track_4.mux_l2_in_5_/X mux_top_track_4.mux_l2_in_4_/X
+ mux_top_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ repeater259/X mux_top_track_24.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2__A0 input62/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 _066_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_ repeater250/X mux_left_track_5.mux_l4_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l5_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input106_A right_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ repeater253/X mux_left_track_17.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input71_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_3_ _121_/A input112/X repeater229/A VGND VGND VPWR VPWR
+ mux_right_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_ repeater255/X mux_top_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_right_track_16.mux_l2_in_1__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_3_ _062_/A input120/X repeater223/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_6__A1 _131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater239 repeater240/X VGND VGND VPWR VPWR repeater239/X sky130_fd_sc_hd__clkbuf_1
Xrepeater228 repeater228/A VGND VGND VPWR VPWR repeater228/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input34_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_119_ _119_/A VGND VGND VPWR VPWR _119_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_3__A0 _130_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_ repeater263/X mux_bottom_track_33.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_3__283 VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_3_/A0
+ mux_right_track_32.mux_l1_in_3__283/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_24.mux_l1_in_2__A0 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l1_in_1_ _059_/A _109_/A repeater234/A VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_2__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A1 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ repeater250/X mux_left_track_5.mux_l3_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_16.mux_l2_in_1__A0 _134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input64_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_2_ input110/X input108/X repeater229/A VGND VGND VPWR
+ VPWR mux_right_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ repeater248/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_2_ input119/X input118/X repeater224/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_3_ mux_left_track_33.mux_l1_in_3_/A0 input101/X mux_left_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_135_ _135_/A VGND VGND VPWR VPWR _135_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_17.mux_l2_in_3_ mux_bottom_track_17.mux_l2_in_3_/A0 _094_/A mux_bottom_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater229 repeater229/A VGND VGND VPWR VPWR repeater229/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input27_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_118_ _118_/A VGND VGND VPWR VPWR _118_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_ repeater254/X mux_top_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ output122/A VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l1_in_2__A0 _126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ repeater265/X mux_bottom_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_3_ mux_bottom_track_3.mux_l2_in_3_/A0 _090_/A mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l4_in_0_ mux_bottom_track_17.mux_l3_in_1_/X mux_bottom_track_17.mux_l3_in_0_/X
+ mux_bottom_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l1_in_0_ _099_/A input71/X repeater234/X VGND VGND VPWR VPWR
+ mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input94_A left_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_ repeater259/X mux_top_track_24.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_16.mux_l1_in_2__A1 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_1_ mux_left_track_33.mux_l1_in_3_/X mux_left_track_33.mux_l1_in_2_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l2_in_1__A0 _135_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ repeater269/X mux_right_track_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_4_ input24/X input9/X repeater237/A VGND VGND VPWR VPWR
+ mux_bottom_track_3.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_17.mux_l3_in_1_ mux_bottom_track_17.mux_l2_in_3_/X mux_bottom_track_17.mux_l2_in_2_/X
+ mux_bottom_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_ repeater252/X mux_left_track_17.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input1_A Test_en_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ repeater240/X repeater232/X VGND VGND
+ VPWR VPWR mux_left_track_5.mux_l3_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input57_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_2.mux_l1_in_1_ input106/X _110_/A repeater229/X VGND VGND VPWR VPWR
+ mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ repeater248/X repeater225/A VGND VGND
+ VPWR VPWR mux_top_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ input117/X input116/X repeater224/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ input97/X input57/X mux_left_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _132_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input111_A right_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _133_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_3_S_FTB01 input104/X VGND VGND VPWR VPWR output221/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l2_in_2_ input17/X _085_/A mux_bottom_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_065_ _065_/A VGND VGND VPWR VPWR _065_/X sky130_fd_sc_hd__clkbuf_1
X_134_ _134_/A VGND VGND VPWR VPWR _134_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_117_ _117_/A VGND VGND VPWR VPWR _117_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_32.mux_l1_in_2__A1 _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ repeater254/X mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xprog_clk_1_E_FTB01 input103/X VGND VGND VPWR VPWR output213/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ repeater265/X mux_bottom_track_25.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_4.mux_l2_in_5__A0 _131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.mux_l2_in_7__291 VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_7_/A0
+ mux_top_track_4.mux_l2_in_7__291/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_3.mux_l2_in_2_ _081_/A mux_bottom_track_3.mux_l1_in_4_/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 input81/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ repeater260/X mux_top_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input87_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ repeater269/X mux_right_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l2_in_1__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_3_ input7/X input5/X repeater237/X VGND VGND VPWR VPWR
+ mux_bottom_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ repeater248/X mux_left_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ repeater245/X mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR repeater232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XTest_en_N_FTB01 input1/X VGND VGND VPWR VPWR output121/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l1_in_0_ _101_/A input71/X repeater229/X VGND VGND VPWR VPWR
+ mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ repeater255/X mux_top_track_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR repeater225/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_1_ _127_/A _067_/A mux_left_track_33.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_0_ input115/X mux_top_track_4.mux_l1_in_0_/X repeater224/A
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input104_A prog_clk_3_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_3__A1 _094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l5_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__clkbuf_1
X_133_ _133_/A VGND VGND VPWR VPWR _133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l2_in_1_ input7/X mux_bottom_track_17.mux_l1_in_2_/X mux_bottom_track_17.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_064_ _064_/A VGND VGND VPWR VPWR _064_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__110__A _110_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ repeater267/X mux_right_track_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_32.mux_l1_in_2__A1 _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l2_in_3__289 VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_3_/A0
+ mux_top_track_24.mux_l2_in_3__289/LO sky130_fd_sc_hd__conb_1
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_25.mux_l1_in_2__A0 _126_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ repeater253/X mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_2_ input3/X _074_/A mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l2_in_5__A1 _122_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2__A1 _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ repeater260/X mux_top_track_24.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ repeater272/X repeater229/X VGND VGND
+ VPWR VPWR mux_right_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_2_ input3/X _070_/A repeater237/X VGND VGND VPWR VPWR
+ mux_bottom_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ repeater253/X mux_left_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ repeater241/X mux_left_track_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_0_ _107_/A input82/X mux_left_track_33.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_132_ _132_/A VGND VGND VPWR VPWR _132_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_063_ _063_/A VGND VGND VPWR VPWR _063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ repeater267/X mux_right_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ input114/X input113/X mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_5.mux_l2_in_3__A1 _131_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_2__A1 _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_ repeater266/X mux_bottom_track_25.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ repeater257/X mux_top_track_4.mux_l5_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_17.mux_l1_in_1_ _065_/A input42/X mux_bottom_track_17.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input25_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ repeater258/X mux_top_track_16.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

