magic
tech sky130A
magscale 1 2
timestamp 1656943209
<< viali >>
rect 6929 17289 6963 17323
rect 7205 17289 7239 17323
rect 8493 17289 8527 17323
rect 11529 17289 11563 17323
rect 12449 17289 12483 17323
rect 13001 17289 13035 17323
rect 13369 17289 13403 17323
rect 8033 17221 8067 17255
rect 10425 17221 10459 17255
rect 10885 17221 10919 17255
rect 11989 17221 12023 17255
rect 13645 17221 13679 17255
rect 6469 17153 6503 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 7941 17153 7975 17187
rect 8677 17153 8711 17187
rect 10333 17153 10367 17187
rect 11345 17153 11379 17187
rect 13185 17153 13219 17187
rect 13553 17153 13587 17187
rect 14473 17153 14507 17187
rect 6653 17085 6687 17119
rect 8217 17085 8251 17119
rect 9229 17085 9263 17119
rect 9597 17085 9631 17119
rect 10609 17085 10643 17119
rect 12541 17085 12575 17119
rect 12633 17085 12667 17119
rect 13921 17085 13955 17119
rect 11161 17017 11195 17051
rect 14105 17017 14139 17051
rect 14289 17017 14323 17051
rect 4445 16949 4479 16983
rect 4813 16949 4847 16983
rect 5273 16949 5307 16983
rect 5641 16949 5675 16983
rect 6009 16949 6043 16983
rect 7573 16949 7607 16983
rect 8953 16949 8987 16983
rect 9321 16949 9355 16983
rect 9689 16949 9723 16983
rect 9965 16949 9999 16983
rect 11713 16949 11747 16983
rect 12081 16949 12115 16983
rect 3157 16745 3191 16779
rect 7665 16745 7699 16779
rect 13093 16745 13127 16779
rect 6561 16609 6595 16643
rect 7297 16609 7331 16643
rect 8309 16609 8343 16643
rect 10241 16609 10275 16643
rect 10977 16609 11011 16643
rect 11069 16609 11103 16643
rect 11621 16609 11655 16643
rect 12817 16609 12851 16643
rect 13553 16609 13587 16643
rect 13645 16609 13679 16643
rect 14473 16609 14507 16643
rect 15485 16609 15519 16643
rect 1777 16541 1811 16575
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 2605 16541 2639 16575
rect 2973 16541 3007 16575
rect 3341 16541 3375 16575
rect 4353 16541 4387 16575
rect 4721 16541 4755 16575
rect 5089 16541 5123 16575
rect 5457 16541 5491 16575
rect 5825 16541 5859 16575
rect 7113 16541 7147 16575
rect 8125 16541 8159 16575
rect 8585 16541 8619 16575
rect 9229 16541 9263 16575
rect 9597 16541 9631 16575
rect 10057 16541 10091 16575
rect 12633 16541 12667 16575
rect 6285 16473 6319 16507
rect 7205 16473 7239 16507
rect 11805 16473 11839 16507
rect 12725 16473 12759 16507
rect 14565 16473 14599 16507
rect 2789 16405 2823 16439
rect 3525 16405 3559 16439
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 4537 16405 4571 16439
rect 4905 16405 4939 16439
rect 5273 16405 5307 16439
rect 5641 16405 5675 16439
rect 5917 16405 5951 16439
rect 6377 16405 6411 16439
rect 6745 16405 6779 16439
rect 7757 16405 7791 16439
rect 8217 16405 8251 16439
rect 9045 16405 9079 16439
rect 9413 16405 9447 16439
rect 9689 16405 9723 16439
rect 10149 16405 10183 16439
rect 10517 16405 10551 16439
rect 10885 16405 10919 16439
rect 11713 16405 11747 16439
rect 12173 16405 12207 16439
rect 12265 16405 12299 16439
rect 13461 16405 13495 16439
rect 14197 16405 14231 16439
rect 1685 16201 1719 16235
rect 2605 16201 2639 16235
rect 3709 16201 3743 16235
rect 4905 16201 4939 16235
rect 5365 16201 5399 16235
rect 5825 16201 5859 16235
rect 9045 16201 9079 16235
rect 9413 16201 9447 16235
rect 9505 16201 9539 16235
rect 9965 16201 9999 16235
rect 10793 16201 10827 16235
rect 11161 16201 11195 16235
rect 11529 16201 11563 16235
rect 11989 16201 12023 16235
rect 12725 16201 12759 16235
rect 13185 16201 13219 16235
rect 14565 16201 14599 16235
rect 15393 16133 15427 16167
rect 1869 16065 1903 16099
rect 2789 16065 2823 16099
rect 3525 16065 3559 16099
rect 5733 16065 5767 16099
rect 6745 16065 6779 16099
rect 8677 16065 8711 16099
rect 10333 16065 10367 16099
rect 11345 16065 11379 16099
rect 11897 16065 11931 16099
rect 12633 16065 12667 16099
rect 13093 16065 13127 16099
rect 13921 16065 13955 16099
rect 15117 16065 15151 16099
rect 4997 15997 5031 16031
rect 5181 15997 5215 16031
rect 6009 15997 6043 16031
rect 6837 15997 6871 16031
rect 6929 15997 6963 16031
rect 8125 15997 8159 16031
rect 8401 15997 8435 16031
rect 8585 15997 8619 16031
rect 9321 15997 9355 16031
rect 10425 15997 10459 16031
rect 10517 15997 10551 16031
rect 12081 15997 12115 16031
rect 13277 15997 13311 16031
rect 14289 15997 14323 16031
rect 6377 15929 6411 15963
rect 7297 15929 7331 15963
rect 13553 15929 13587 15963
rect 14473 15929 14507 15963
rect 1961 15861 1995 15895
rect 2973 15861 3007 15895
rect 3893 15861 3927 15895
rect 4537 15861 4571 15895
rect 7389 15861 7423 15895
rect 7573 15861 7607 15895
rect 7941 15861 7975 15895
rect 9873 15861 9907 15895
rect 12449 15861 12483 15895
rect 15025 15861 15059 15895
rect 2605 15657 2639 15691
rect 6377 15657 6411 15691
rect 8953 15657 8987 15691
rect 10241 15657 10275 15691
rect 11253 15657 11287 15691
rect 11897 15657 11931 15691
rect 13461 15657 13495 15691
rect 4077 15589 4111 15623
rect 8033 15589 8067 15623
rect 3341 15521 3375 15555
rect 4813 15521 4847 15555
rect 5917 15521 5951 15555
rect 6929 15521 6963 15555
rect 7389 15521 7423 15555
rect 8585 15521 8619 15555
rect 9505 15521 9539 15555
rect 10793 15521 10827 15555
rect 12541 15521 12575 15555
rect 13185 15521 13219 15555
rect 2789 15453 2823 15487
rect 3617 15453 3651 15487
rect 4537 15453 4571 15487
rect 6745 15453 6779 15487
rect 9413 15453 9447 15487
rect 9781 15453 9815 15487
rect 10609 15453 10643 15487
rect 12265 15453 12299 15487
rect 7481 15385 7515 15419
rect 8493 15385 8527 15419
rect 11805 15385 11839 15419
rect 12357 15385 12391 15419
rect 2973 15317 3007 15351
rect 4169 15317 4203 15351
rect 4629 15317 4663 15351
rect 5089 15317 5123 15351
rect 6193 15317 6227 15351
rect 6837 15317 6871 15351
rect 7573 15317 7607 15351
rect 7941 15317 7975 15351
rect 8401 15317 8435 15351
rect 9321 15317 9355 15351
rect 9965 15317 9999 15351
rect 10701 15317 10735 15351
rect 11069 15317 11103 15351
rect 11529 15317 11563 15351
rect 12817 15317 12851 15351
rect 13277 15317 13311 15351
rect 14105 15317 14139 15351
rect 14565 15317 14599 15351
rect 14749 15317 14783 15351
rect 3617 15113 3651 15147
rect 4169 15113 4203 15147
rect 4445 15113 4479 15147
rect 4905 15113 4939 15147
rect 5273 15113 5307 15147
rect 5641 15113 5675 15147
rect 6561 15113 6595 15147
rect 7021 15113 7055 15147
rect 7389 15113 7423 15147
rect 7757 15113 7791 15147
rect 8677 15113 8711 15147
rect 9045 15113 9079 15147
rect 9873 15113 9907 15147
rect 9965 15113 9999 15147
rect 11253 15113 11287 15147
rect 11897 15113 11931 15147
rect 12357 15113 12391 15147
rect 12817 15113 12851 15147
rect 14381 15113 14415 15147
rect 14841 15113 14875 15147
rect 6469 15045 6503 15079
rect 8401 15045 8435 15079
rect 10333 15045 10367 15079
rect 2053 14977 2087 15011
rect 3525 14977 3559 15011
rect 4353 14977 4387 15011
rect 4813 14977 4847 15011
rect 6929 14977 6963 15011
rect 7849 14977 7883 15011
rect 12725 14977 12759 15011
rect 13553 14977 13587 15011
rect 15209 14977 15243 15011
rect 1777 14909 1811 14943
rect 3801 14909 3835 14943
rect 4997 14909 5031 14943
rect 5733 14909 5767 14943
rect 5917 14909 5951 14943
rect 7205 14909 7239 14943
rect 8033 14909 8067 14943
rect 9137 14909 9171 14943
rect 9321 14909 9355 14943
rect 10149 14909 10183 14943
rect 11713 14909 11747 14943
rect 11805 14909 11839 14943
rect 12909 14909 12943 14943
rect 13277 14909 13311 14943
rect 13461 14909 13495 14943
rect 14105 14909 14139 14943
rect 14289 14909 14323 14943
rect 15301 14909 15335 14943
rect 15393 14909 15427 14943
rect 9505 14841 9539 14875
rect 12265 14841 12299 14875
rect 3157 14773 3191 14807
rect 6193 14773 6227 14807
rect 8585 14773 8619 14807
rect 11069 14773 11103 14807
rect 13921 14773 13955 14807
rect 14749 14773 14783 14807
rect 4905 14569 4939 14603
rect 5089 14569 5123 14603
rect 5917 14569 5951 14603
rect 7297 14569 7331 14603
rect 8401 14569 8435 14603
rect 9965 14569 9999 14603
rect 11529 14569 11563 14603
rect 14933 14569 14967 14603
rect 4721 14501 4755 14535
rect 8125 14501 8159 14535
rect 9781 14501 9815 14535
rect 1685 14433 1719 14467
rect 2881 14433 2915 14467
rect 4353 14433 4387 14467
rect 5733 14433 5767 14467
rect 6469 14433 6503 14467
rect 7757 14433 7791 14467
rect 7941 14433 7975 14467
rect 14565 14433 14599 14467
rect 14657 14433 14691 14467
rect 15485 14433 15519 14467
rect 1961 14365 1995 14399
rect 4169 14365 4203 14399
rect 5457 14365 5491 14399
rect 7665 14365 7699 14399
rect 8953 14365 8987 14399
rect 11253 14365 11287 14399
rect 11437 14365 11471 14399
rect 13185 14365 13219 14399
rect 14473 14365 14507 14399
rect 3065 14297 3099 14331
rect 6377 14297 6411 14331
rect 6837 14297 6871 14331
rect 12940 14297 12974 14331
rect 15393 14297 15427 14331
rect 3157 14229 3191 14263
rect 3525 14229 3559 14263
rect 3801 14229 3835 14263
rect 4261 14229 4295 14263
rect 5549 14229 5583 14263
rect 6285 14229 6319 14263
rect 6929 14229 6963 14263
rect 8585 14229 8619 14263
rect 11805 14229 11839 14263
rect 13829 14229 13863 14263
rect 14105 14229 14139 14263
rect 15301 14229 15335 14263
rect 3617 14025 3651 14059
rect 4721 14025 4755 14059
rect 7757 14025 7791 14059
rect 8493 14025 8527 14059
rect 8861 14025 8895 14059
rect 9229 14025 9263 14059
rect 9321 14025 9355 14059
rect 9689 14025 9723 14059
rect 10149 14025 10183 14059
rect 10517 14025 10551 14059
rect 11345 14025 11379 14059
rect 12909 14025 12943 14059
rect 3433 13957 3467 13991
rect 5856 13957 5890 13991
rect 6622 13957 6656 13991
rect 10057 13957 10091 13991
rect 10885 13957 10919 13991
rect 11796 13957 11830 13991
rect 14565 13957 14599 13991
rect 15485 13957 15519 13991
rect 15577 13957 15611 13991
rect 2697 13889 2731 13923
rect 3249 13889 3283 13923
rect 4629 13889 4663 13923
rect 10977 13889 11011 13923
rect 13001 13889 13035 13923
rect 2789 13821 2823 13855
rect 2973 13821 3007 13855
rect 6101 13821 6135 13855
rect 6377 13821 6411 13855
rect 8309 13821 8343 13855
rect 8401 13821 8435 13855
rect 9137 13821 9171 13855
rect 9873 13821 9907 13855
rect 10701 13821 10735 13855
rect 11529 13821 11563 13855
rect 14473 13821 14507 13855
rect 7849 13753 7883 13787
rect 2329 13685 2363 13719
rect 5273 13481 5307 13515
rect 5549 13481 5583 13515
rect 7297 13481 7331 13515
rect 11253 13481 11287 13515
rect 12909 13481 12943 13515
rect 15163 13481 15197 13515
rect 15577 13481 15611 13515
rect 2881 13413 2915 13447
rect 5641 13413 5675 13447
rect 8769 13413 8803 13447
rect 2237 13345 2271 13379
rect 3525 13345 3559 13379
rect 7021 13345 7055 13379
rect 7389 13345 7423 13379
rect 9045 13345 9079 13379
rect 11345 13345 11379 13379
rect 14657 13345 14691 13379
rect 1961 13277 1995 13311
rect 2421 13277 2455 13311
rect 3249 13277 3283 13311
rect 3893 13277 3927 13311
rect 9781 13277 9815 13311
rect 9873 13277 9907 13311
rect 14565 13277 14599 13311
rect 15060 13277 15094 13311
rect 1685 13209 1719 13243
rect 3341 13209 3375 13243
rect 4138 13209 4172 13243
rect 6754 13209 6788 13243
rect 7656 13209 7690 13243
rect 10140 13209 10174 13243
rect 11590 13209 11624 13243
rect 2329 13141 2363 13175
rect 2789 13141 2823 13175
rect 9137 13141 9171 13175
rect 12725 13141 12759 13175
rect 14105 13141 14139 13175
rect 14473 13141 14507 13175
rect 2421 12937 2455 12971
rect 6193 12937 6227 12971
rect 7297 12937 7331 12971
rect 13369 12937 13403 12971
rect 13737 12937 13771 12971
rect 14289 12937 14323 12971
rect 14657 12937 14691 12971
rect 15117 12937 15151 12971
rect 2789 12869 2823 12903
rect 8953 12869 8987 12903
rect 11345 12869 11379 12903
rect 11774 12869 11808 12903
rect 14749 12869 14783 12903
rect 2329 12801 2363 12835
rect 2881 12801 2915 12835
rect 4454 12801 4488 12835
rect 4721 12801 4755 12835
rect 4813 12801 4847 12835
rect 5080 12801 5114 12835
rect 7389 12801 7423 12835
rect 7645 12801 7679 12835
rect 10158 12801 10192 12835
rect 10425 12801 10459 12835
rect 11529 12801 11563 12835
rect 13829 12801 13863 12835
rect 3065 12733 3099 12767
rect 13645 12733 13679 12767
rect 14841 12733 14875 12767
rect 8769 12665 8803 12699
rect 9045 12665 9079 12699
rect 12909 12665 12943 12699
rect 14197 12665 14231 12699
rect 3341 12597 3375 12631
rect 2881 12393 2915 12427
rect 6745 12393 6779 12427
rect 11253 12393 11287 12427
rect 14105 12393 14139 12427
rect 15209 12393 15243 12427
rect 11161 12325 11195 12359
rect 2237 12257 2271 12291
rect 3525 12257 3559 12291
rect 13277 12257 13311 12291
rect 13461 12257 13495 12291
rect 14749 12257 14783 12291
rect 2605 12189 2639 12223
rect 3893 12189 3927 12223
rect 4629 12189 4663 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 5457 12189 5491 12223
rect 6653 12189 6687 12223
rect 8125 12189 8159 12223
rect 8769 12189 8803 12223
rect 10333 12189 10367 12223
rect 12633 12189 12667 12223
rect 14565 12189 14599 12223
rect 3249 12121 3283 12155
rect 7880 12121 7914 12155
rect 10088 12121 10122 12155
rect 12388 12121 12422 12155
rect 14473 12121 14507 12155
rect 14933 12121 14967 12155
rect 1593 12053 1627 12087
rect 1961 12053 1995 12087
rect 2053 12053 2087 12087
rect 2789 12053 2823 12087
rect 3341 12053 3375 12087
rect 8953 12053 8987 12087
rect 12817 12053 12851 12087
rect 13185 12053 13219 12087
rect 13645 12053 13679 12087
rect 2513 11849 2547 11883
rect 3433 11849 3467 11883
rect 4077 11849 4111 11883
rect 9505 11849 9539 11883
rect 1777 11781 1811 11815
rect 3985 11781 4019 11815
rect 5190 11781 5224 11815
rect 9413 11781 9447 11815
rect 12265 11781 12299 11815
rect 1501 11713 1535 11747
rect 2605 11713 2639 11747
rect 3341 11713 3375 11747
rect 10629 11713 10663 11747
rect 10885 11713 10919 11747
rect 12357 11713 12391 11747
rect 13737 11713 13771 11747
rect 2789 11645 2823 11679
rect 3525 11645 3559 11679
rect 5457 11645 5491 11679
rect 12449 11645 12483 11679
rect 13829 11645 13863 11679
rect 14013 11645 14047 11679
rect 2145 11509 2179 11543
rect 2973 11509 3007 11543
rect 5641 11509 5675 11543
rect 5825 11509 5859 11543
rect 6009 11509 6043 11543
rect 7297 11509 7331 11543
rect 11897 11509 11931 11543
rect 13185 11509 13219 11543
rect 13369 11509 13403 11543
rect 14289 11509 14323 11543
rect 2053 11305 2087 11339
rect 5825 11305 5859 11339
rect 7297 11305 7331 11339
rect 8769 11305 8803 11339
rect 10517 11305 10551 11339
rect 15025 11305 15059 11339
rect 2881 11237 2915 11271
rect 4077 11237 4111 11271
rect 4353 11237 4387 11271
rect 9045 11237 9079 11271
rect 2605 11169 2639 11203
rect 3525 11169 3559 11203
rect 9137 11169 9171 11203
rect 10609 11169 10643 11203
rect 14565 11169 14599 11203
rect 14657 11169 14691 11203
rect 2421 11101 2455 11135
rect 3341 11101 3375 11135
rect 4445 11101 4479 11135
rect 5917 11101 5951 11135
rect 7389 11101 7423 11135
rect 9404 11101 9438 11135
rect 13461 11101 13495 11135
rect 1961 11033 1995 11067
rect 3249 11033 3283 11067
rect 3801 11033 3835 11067
rect 4690 11033 4724 11067
rect 6184 11033 6218 11067
rect 7656 11033 7690 11067
rect 10854 11033 10888 11067
rect 13194 11033 13228 11067
rect 13921 11033 13955 11067
rect 14473 11033 14507 11067
rect 2513 10965 2547 10999
rect 11989 10965 12023 10999
rect 12081 10965 12115 10999
rect 14105 10965 14139 10999
rect 1869 10761 1903 10795
rect 2237 10761 2271 10795
rect 2329 10761 2363 10795
rect 2697 10761 2731 10795
rect 3157 10761 3191 10795
rect 3525 10761 3559 10795
rect 4721 10761 4755 10795
rect 6469 10761 6503 10795
rect 8033 10761 8067 10795
rect 8861 10761 8895 10795
rect 10333 10761 10367 10795
rect 10517 10761 10551 10795
rect 11989 10761 12023 10795
rect 12633 10761 12667 10795
rect 13277 10761 13311 10795
rect 3985 10693 4019 10727
rect 5834 10693 5868 10727
rect 9220 10693 9254 10727
rect 12081 10693 12115 10727
rect 13185 10693 13219 10727
rect 3065 10625 3099 10659
rect 3893 10625 3927 10659
rect 4445 10625 4479 10659
rect 7582 10625 7616 10659
rect 7849 10625 7883 10659
rect 8953 10625 8987 10659
rect 2513 10557 2547 10591
rect 3341 10557 3375 10591
rect 4169 10557 4203 10591
rect 6101 10557 6135 10591
rect 11897 10557 11931 10591
rect 13369 10557 13403 10591
rect 4537 10421 4571 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 3157 10217 3191 10251
rect 3893 10217 3927 10251
rect 8769 10217 8803 10251
rect 10057 10217 10091 10251
rect 14381 10217 14415 10251
rect 1685 10081 1719 10115
rect 10149 10081 10183 10115
rect 13185 10081 13219 10115
rect 15117 10081 15151 10115
rect 1961 10013 1995 10047
rect 2237 10013 2271 10047
rect 2513 10013 2547 10047
rect 5006 10013 5040 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 5825 10013 5859 10047
rect 7297 10013 7331 10047
rect 7389 10013 7423 10047
rect 15025 10013 15059 10047
rect 7052 9945 7086 9979
rect 7656 9945 7690 9979
rect 10416 9945 10450 9979
rect 13001 9945 13035 9979
rect 14933 9945 14967 9979
rect 15393 9945 15427 9979
rect 2973 9877 3007 9911
rect 3433 9877 3467 9911
rect 3617 9877 3651 9911
rect 5917 9877 5951 9911
rect 11529 9877 11563 9911
rect 12633 9877 12667 9911
rect 13093 9877 13127 9911
rect 14565 9877 14599 9911
rect 5733 9673 5767 9707
rect 9597 9673 9631 9707
rect 13185 9673 13219 9707
rect 14289 9673 14323 9707
rect 14749 9673 14783 9707
rect 7604 9605 7638 9639
rect 11253 9605 11287 9639
rect 1961 9537 1995 9571
rect 2697 9537 2731 9571
rect 5374 9537 5408 9571
rect 5641 9537 5675 9571
rect 6101 9537 6135 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 8125 9537 8159 9571
rect 8381 9537 8415 9571
rect 10721 9537 10755 9571
rect 10977 9537 11011 9571
rect 12653 9537 12687 9571
rect 12909 9537 12943 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 1685 9469 1719 9503
rect 2789 9469 2823 9503
rect 2973 9469 3007 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 14841 9469 14875 9503
rect 15301 9469 15335 9503
rect 4261 9401 4295 9435
rect 11529 9401 11563 9435
rect 2329 9333 2363 9367
rect 6469 9333 6503 9367
rect 9505 9333 9539 9367
rect 2053 9129 2087 9163
rect 3985 9129 4019 9163
rect 4169 9129 4203 9163
rect 9505 9129 9539 9163
rect 9965 9129 9999 9163
rect 14105 9129 14139 9163
rect 14933 9129 14967 9163
rect 10057 9061 10091 9095
rect 12909 9061 12943 9095
rect 2513 8993 2547 9027
rect 2697 8993 2731 9027
rect 3341 8993 3375 9027
rect 3525 8993 3559 9027
rect 5917 8993 5951 9027
rect 11529 8993 11563 9027
rect 13093 8993 13127 9027
rect 14749 8993 14783 9027
rect 15485 8993 15519 9027
rect 4445 8925 4479 8959
rect 11437 8925 11471 8959
rect 11785 8925 11819 8959
rect 15301 8925 15335 8959
rect 15393 8925 15427 8959
rect 2421 8857 2455 8891
rect 3249 8857 3283 8891
rect 4690 8857 4724 8891
rect 6162 8857 6196 8891
rect 11192 8857 11226 8891
rect 13369 8857 13403 8891
rect 2881 8789 2915 8823
rect 5825 8789 5859 8823
rect 7297 8789 7331 8823
rect 13277 8789 13311 8823
rect 13737 8789 13771 8823
rect 14473 8789 14507 8823
rect 14565 8789 14599 8823
rect 1777 8585 1811 8619
rect 2237 8585 2271 8619
rect 2605 8585 2639 8619
rect 3157 8585 3191 8619
rect 3985 8585 4019 8619
rect 5549 8585 5583 8619
rect 10701 8585 10735 8619
rect 11529 8585 11563 8619
rect 12081 8585 12115 8619
rect 12725 8585 12759 8619
rect 13369 8585 13403 8619
rect 13829 8585 13863 8619
rect 14105 8585 14139 8619
rect 14381 8585 14415 8619
rect 14841 8585 14875 8619
rect 15669 8585 15703 8619
rect 2145 8517 2179 8551
rect 3065 8517 3099 8551
rect 5825 8517 5859 8551
rect 6009 8517 6043 8551
rect 6193 8517 6227 8551
rect 7205 8517 7239 8551
rect 7389 8517 7423 8551
rect 13461 8517 13495 8551
rect 13921 8517 13955 8551
rect 14749 8517 14783 8551
rect 4169 8449 4203 8483
rect 4425 8449 4459 8483
rect 8594 8449 8628 8483
rect 8861 8449 8895 8483
rect 8953 8449 8987 8483
rect 9220 8449 9254 8483
rect 2053 8381 2087 8415
rect 3341 8381 3375 8415
rect 3525 8381 3559 8415
rect 13277 8381 13311 8415
rect 14933 8381 14967 8415
rect 7481 8313 7515 8347
rect 10333 8313 10367 8347
rect 12817 8313 12851 8347
rect 2697 8245 2731 8279
rect 3801 8245 3835 8279
rect 2789 8041 2823 8075
rect 3893 8041 3927 8075
rect 7205 8041 7239 8075
rect 8953 8041 8987 8075
rect 9137 8041 9171 8075
rect 12265 8041 12299 8075
rect 13829 8041 13863 8075
rect 14473 8041 14507 8075
rect 15669 8041 15703 8075
rect 12173 7973 12207 8007
rect 14289 7973 14323 8007
rect 1685 7905 1719 7939
rect 2237 7905 2271 7939
rect 3525 7905 3559 7939
rect 6929 7905 6963 7939
rect 8677 7905 8711 7939
rect 9321 7905 9355 7939
rect 15025 7905 15059 7939
rect 1961 7837 1995 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 8410 7837 8444 7871
rect 10793 7837 10827 7871
rect 13645 7837 13679 7871
rect 14841 7837 14875 7871
rect 2329 7769 2363 7803
rect 3341 7769 3375 7803
rect 5028 7769 5062 7803
rect 6684 7769 6718 7803
rect 9588 7769 9622 7803
rect 11060 7769 11094 7803
rect 13378 7769 13412 7803
rect 2421 7701 2455 7735
rect 2881 7701 2915 7735
rect 3249 7701 3283 7735
rect 5549 7701 5583 7735
rect 7297 7701 7331 7735
rect 10701 7701 10735 7735
rect 14933 7701 14967 7735
rect 15301 7701 15335 7735
rect 2789 7497 2823 7531
rect 3157 7497 3191 7531
rect 5825 7497 5859 7531
rect 6101 7497 6135 7531
rect 6653 7497 6687 7531
rect 8217 7497 8251 7531
rect 9873 7497 9907 7531
rect 13001 7497 13035 7531
rect 14197 7497 14231 7531
rect 14289 7497 14323 7531
rect 15209 7497 15243 7531
rect 1685 7429 1719 7463
rect 11796 7429 11830 7463
rect 1961 7361 1995 7395
rect 3249 7361 3283 7395
rect 3985 7361 4019 7395
rect 5466 7361 5500 7395
rect 5733 7361 5767 7395
rect 6745 7361 6779 7395
rect 7012 7361 7046 7395
rect 9330 7361 9364 7395
rect 9597 7361 9631 7395
rect 11078 7361 11112 7395
rect 11345 7361 11379 7395
rect 11529 7361 11563 7395
rect 13369 7361 13403 7395
rect 15117 7361 15151 7395
rect 3433 7293 3467 7327
rect 4077 7293 4111 7327
rect 13461 7293 13495 7327
rect 13553 7293 13587 7327
rect 14381 7293 14415 7327
rect 15301 7293 15335 7327
rect 3801 7225 3835 7259
rect 12909 7225 12943 7259
rect 4353 7157 4387 7191
rect 8125 7157 8159 7191
rect 9965 7157 9999 7191
rect 13829 7157 13863 7191
rect 14749 7157 14783 7191
rect 15577 7157 15611 7191
rect 9045 6953 9079 6987
rect 10333 6953 10367 6987
rect 13921 6953 13955 6987
rect 7297 6885 7331 6919
rect 13737 6885 13771 6919
rect 3433 6817 3467 6851
rect 8769 6817 8803 6851
rect 14657 6817 14691 6851
rect 15393 6817 15427 6851
rect 15485 6817 15519 6851
rect 4169 6749 4203 6783
rect 4436 6749 4470 6783
rect 5917 6749 5951 6783
rect 11897 6749 11931 6783
rect 13369 6749 13403 6783
rect 13553 6749 13587 6783
rect 14473 6749 14507 6783
rect 6184 6681 6218 6715
rect 8524 6681 8558 6715
rect 11630 6681 11664 6715
rect 13102 6681 13136 6715
rect 2789 6613 2823 6647
rect 3157 6613 3191 6647
rect 3249 6613 3283 6647
rect 3893 6613 3927 6647
rect 5549 6613 5583 6647
rect 5825 6613 5859 6647
rect 7389 6613 7423 6647
rect 10517 6613 10551 6647
rect 11989 6613 12023 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 14933 6613 14967 6647
rect 15301 6613 15335 6647
rect 2973 6409 3007 6443
rect 6193 6409 6227 6443
rect 11529 6409 11563 6443
rect 11805 6409 11839 6443
rect 13185 6409 13219 6443
rect 13737 6409 13771 6443
rect 14197 6409 14231 6443
rect 14565 6409 14599 6443
rect 15393 6409 15427 6443
rect 13277 6341 13311 6375
rect 1961 6273 1995 6307
rect 2881 6273 2915 6307
rect 4454 6273 4488 6307
rect 4721 6273 4755 6307
rect 4813 6273 4847 6307
rect 5069 6273 5103 6307
rect 6469 6273 6503 6307
rect 6653 6273 6687 6307
rect 7113 6273 7147 6307
rect 7205 6273 7239 6307
rect 7472 6273 7506 6307
rect 8677 6273 8711 6307
rect 8944 6273 8978 6307
rect 14105 6273 14139 6307
rect 14933 6273 14967 6307
rect 1685 6205 1719 6239
rect 3157 6205 3191 6239
rect 13093 6205 13127 6239
rect 14381 6205 14415 6239
rect 15025 6205 15059 6239
rect 15117 6205 15151 6239
rect 13645 6137 13679 6171
rect 2513 6069 2547 6103
rect 3341 6069 3375 6103
rect 8585 6069 8619 6103
rect 10057 6069 10091 6103
rect 3433 5865 3467 5899
rect 5825 5865 5859 5899
rect 8309 5865 8343 5899
rect 8585 5865 8619 5899
rect 9597 5865 9631 5899
rect 11253 5865 11287 5899
rect 12817 5865 12851 5899
rect 14197 5865 14231 5899
rect 15485 5865 15519 5899
rect 11161 5797 11195 5831
rect 14381 5797 14415 5831
rect 2053 5729 2087 5763
rect 2145 5729 2179 5763
rect 2881 5729 2915 5763
rect 3893 5729 3927 5763
rect 7205 5729 7239 5763
rect 9781 5729 9815 5763
rect 15209 5729 15243 5763
rect 4261 5661 4295 5695
rect 4353 5661 4387 5695
rect 6949 5661 6983 5695
rect 12633 5661 12667 5695
rect 13645 5661 13679 5695
rect 14933 5661 14967 5695
rect 3065 5593 3099 5627
rect 4598 5593 4632 5627
rect 7481 5593 7515 5627
rect 10026 5593 10060 5627
rect 12388 5593 12422 5627
rect 2237 5525 2271 5559
rect 2605 5525 2639 5559
rect 2973 5525 3007 5559
rect 3525 5525 3559 5559
rect 5733 5525 5767 5559
rect 13737 5525 13771 5559
rect 2237 5321 2271 5355
rect 2881 5321 2915 5355
rect 3525 5321 3559 5355
rect 3985 5321 4019 5355
rect 4629 5321 4663 5355
rect 5457 5321 5491 5355
rect 6469 5321 6503 5355
rect 7021 5321 7055 5355
rect 7389 5321 7423 5355
rect 9781 5321 9815 5355
rect 11161 5321 11195 5355
rect 13277 5321 13311 5355
rect 2605 5253 2639 5287
rect 3893 5253 3927 5287
rect 4353 5253 4387 5287
rect 8646 5253 8680 5287
rect 13369 5253 13403 5287
rect 1869 5185 1903 5219
rect 2329 5185 2363 5219
rect 3157 5185 3191 5219
rect 4997 5185 5031 5219
rect 5825 5185 5859 5219
rect 6929 5185 6963 5219
rect 7757 5185 7791 5219
rect 8401 5185 8435 5219
rect 10241 5185 10275 5219
rect 12449 5185 12483 5219
rect 14105 5185 14139 5219
rect 14749 5185 14783 5219
rect 1593 5117 1627 5151
rect 1777 5117 1811 5151
rect 4077 5117 4111 5151
rect 5089 5117 5123 5151
rect 5273 5117 5307 5151
rect 5917 5117 5951 5151
rect 6101 5117 6135 5151
rect 7113 5117 7147 5151
rect 7849 5117 7883 5151
rect 7941 5117 7975 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 11989 5117 12023 5151
rect 12541 5117 12575 5151
rect 12633 5117 12667 5151
rect 13461 5117 13495 5151
rect 14197 5117 14231 5151
rect 14289 5117 14323 5151
rect 6561 4981 6595 5015
rect 8217 4981 8251 5015
rect 9873 4981 9907 5015
rect 12081 4981 12115 5015
rect 12909 4981 12943 5015
rect 13737 4981 13771 5015
rect 14565 4981 14599 5015
rect 1869 4777 1903 4811
rect 2881 4777 2915 4811
rect 4905 4777 4939 4811
rect 5733 4777 5767 4811
rect 6193 4777 6227 4811
rect 9137 4777 9171 4811
rect 10333 4777 10367 4811
rect 11529 4777 11563 4811
rect 13185 4777 13219 4811
rect 15025 4777 15059 4811
rect 3801 4709 3835 4743
rect 5825 4709 5859 4743
rect 8585 4709 8619 4743
rect 2513 4641 2547 4675
rect 3525 4641 3559 4675
rect 4353 4641 4387 4675
rect 6101 4641 6135 4675
rect 6653 4641 6687 4675
rect 6745 4641 6779 4675
rect 7113 4641 7147 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 8769 4641 8803 4675
rect 9781 4641 9815 4675
rect 12081 4641 12115 4675
rect 13001 4641 13035 4675
rect 13645 4641 13679 4675
rect 13737 4641 13771 4675
rect 14657 4641 14691 4675
rect 2237 4573 2271 4607
rect 7389 4573 7423 4607
rect 8953 4573 8987 4607
rect 12725 4573 12759 4607
rect 12817 4573 12851 4607
rect 14473 4573 14507 4607
rect 14565 4573 14599 4607
rect 3249 4505 3283 4539
rect 4629 4505 4663 4539
rect 11345 4505 11379 4539
rect 11897 4505 11931 4539
rect 13553 4505 13587 4539
rect 2329 4437 2363 4471
rect 3341 4437 3375 4471
rect 4169 4437 4203 4471
rect 4261 4437 4295 4471
rect 5089 4437 5123 4471
rect 5549 4437 5583 4471
rect 6561 4437 6595 4471
rect 7757 4437 7791 4471
rect 8125 4437 8159 4471
rect 8217 4437 8251 4471
rect 9873 4437 9907 4471
rect 9965 4437 9999 4471
rect 11069 4437 11103 4471
rect 11989 4437 12023 4471
rect 12357 4437 12391 4471
rect 14105 4437 14139 4471
rect 1685 4233 1719 4267
rect 2053 4233 2087 4267
rect 2973 4233 3007 4267
rect 4629 4233 4663 4267
rect 4997 4233 5031 4267
rect 5457 4233 5491 4267
rect 5825 4233 5859 4267
rect 6469 4233 6503 4267
rect 7941 4233 7975 4267
rect 8033 4233 8067 4267
rect 8401 4233 8435 4267
rect 9413 4233 9447 4267
rect 10333 4233 10367 4267
rect 10701 4233 10735 4267
rect 11529 4233 11563 4267
rect 11989 4233 12023 4267
rect 12817 4233 12851 4267
rect 13277 4233 13311 4267
rect 9505 4165 9539 4199
rect 11253 4165 11287 4199
rect 11897 4165 11931 4199
rect 2145 4097 2179 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 4169 4097 4203 4131
rect 5089 4097 5123 4131
rect 5917 4097 5951 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 12633 4097 12667 4131
rect 2329 4029 2363 4063
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 4445 4029 4479 4063
rect 5181 4029 5215 4063
rect 6009 4029 6043 4063
rect 7205 4029 7239 4063
rect 7849 4029 7883 4063
rect 9321 4029 9355 4063
rect 10793 4029 10827 4063
rect 10885 4029 10919 4063
rect 12081 4029 12115 4063
rect 6653 3961 6687 3995
rect 9873 3961 9907 3995
rect 3801 3893 3835 3927
rect 12357 3893 12391 3927
rect 2697 3689 2731 3723
rect 3617 3689 3651 3723
rect 3985 3689 4019 3723
rect 4445 3689 4479 3723
rect 5273 3689 5307 3723
rect 6009 3689 6043 3723
rect 7849 3689 7883 3723
rect 9781 3689 9815 3723
rect 10517 3689 10551 3723
rect 11345 3689 11379 3723
rect 12173 3689 12207 3723
rect 7757 3621 7791 3655
rect 13829 3621 13863 3655
rect 1777 3553 1811 3587
rect 3157 3553 3191 3587
rect 3341 3553 3375 3587
rect 4997 3553 5031 3587
rect 6561 3553 6595 3587
rect 7297 3553 7331 3587
rect 7389 3553 7423 3587
rect 8401 3553 8435 3587
rect 9137 3553 9171 3587
rect 11069 3553 11103 3587
rect 11897 3553 11931 3587
rect 12725 3553 12759 3587
rect 13645 3553 13679 3587
rect 2053 3485 2087 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 4353 3485 4387 3519
rect 4813 3485 4847 3519
rect 5549 3485 5583 3519
rect 5917 3485 5951 3519
rect 7205 3485 7239 3519
rect 8217 3485 8251 3519
rect 10885 3485 10919 3519
rect 2329 3417 2363 3451
rect 4905 3417 4939 3451
rect 6377 3417 6411 3451
rect 8309 3417 8343 3451
rect 8677 3417 8711 3451
rect 11805 3417 11839 3451
rect 12541 3417 12575 3451
rect 4169 3349 4203 3383
rect 5733 3349 5767 3383
rect 6469 3349 6503 3383
rect 6837 3349 6871 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 10149 3349 10183 3383
rect 10241 3349 10275 3383
rect 10977 3349 11011 3383
rect 11713 3349 11747 3383
rect 12633 3349 12667 3383
rect 13001 3349 13035 3383
rect 13369 3349 13403 3383
rect 13461 3349 13495 3383
rect 3157 3145 3191 3179
rect 4537 3145 4571 3179
rect 4905 3145 4939 3179
rect 5365 3145 5399 3179
rect 6377 3145 6411 3179
rect 6837 3145 6871 3179
rect 7297 3145 7331 3179
rect 9413 3145 9447 3179
rect 9781 3145 9815 3179
rect 10609 3145 10643 3179
rect 11529 3145 11563 3179
rect 13093 3145 13127 3179
rect 13461 3145 13495 3179
rect 13553 3145 13587 3179
rect 13921 3145 13955 3179
rect 14933 3145 14967 3179
rect 11897 3077 11931 3111
rect 14841 3077 14875 3111
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 2789 3009 2823 3043
rect 3341 3009 3375 3043
rect 3709 3009 3743 3043
rect 3801 3009 3835 3043
rect 4445 3009 4479 3043
rect 4997 3009 5031 3043
rect 5837 3009 5871 3043
rect 5942 3009 5976 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 8125 3009 8159 3043
rect 8953 3009 8987 3043
rect 9873 3009 9907 3043
rect 10701 3009 10735 3043
rect 11345 3009 11379 3043
rect 12633 3009 12667 3043
rect 14657 3009 14691 3043
rect 15117 3009 15151 3043
rect 2973 2941 3007 2975
rect 5089 2941 5123 2975
rect 7021 2941 7055 2975
rect 7849 2941 7883 2975
rect 8033 2941 8067 2975
rect 9045 2941 9079 2975
rect 9137 2941 9171 2975
rect 10057 2941 10091 2975
rect 10793 2941 10827 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 12817 2941 12851 2975
rect 13001 2941 13035 2975
rect 14013 2941 14047 2975
rect 14105 2941 14139 2975
rect 15393 2941 15427 2975
rect 2605 2873 2639 2907
rect 4261 2873 4295 2907
rect 5641 2873 5675 2907
rect 10241 2873 10275 2907
rect 14473 2873 14507 2907
rect 1869 2805 1903 2839
rect 2237 2805 2271 2839
rect 3525 2805 3559 2839
rect 3985 2805 4019 2839
rect 6101 2805 6135 2839
rect 7573 2805 7607 2839
rect 8493 2805 8527 2839
rect 8585 2805 8619 2839
rect 11161 2805 11195 2839
rect 12449 2805 12483 2839
rect 2145 2601 2179 2635
rect 2513 2601 2547 2635
rect 3065 2601 3099 2635
rect 3617 2601 3651 2635
rect 3249 2533 3283 2567
rect 4629 2533 4663 2567
rect 4813 2533 4847 2567
rect 5549 2533 5583 2567
rect 5825 2533 5859 2567
rect 6009 2533 6043 2567
rect 6929 2533 6963 2567
rect 7297 2533 7331 2567
rect 7757 2533 7791 2567
rect 8033 2533 8067 2567
rect 8953 2533 8987 2567
rect 10885 2533 10919 2567
rect 13553 2533 13587 2567
rect 13645 2533 13679 2567
rect 4077 2465 4111 2499
rect 7389 2465 7423 2499
rect 8493 2465 8527 2499
rect 8677 2465 8711 2499
rect 10241 2465 10275 2499
rect 11161 2465 11195 2499
rect 12449 2465 12483 2499
rect 12909 2465 12943 2499
rect 3433 2397 3467 2431
rect 4445 2397 4479 2431
rect 4997 2397 5031 2431
rect 5365 2397 5399 2431
rect 6193 2397 6227 2431
rect 6745 2397 6779 2431
rect 7113 2397 7147 2431
rect 7665 2397 7699 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 2881 2329 2915 2363
rect 8401 2329 8435 2363
rect 9137 2329 9171 2363
rect 11621 2329 11655 2363
rect 13829 2329 13863 2363
rect 3801 2261 3835 2295
rect 4261 2261 4295 2295
rect 5181 2261 5215 2295
rect 6561 2261 6595 2295
rect 9413 2261 9447 2295
rect 9689 2261 9723 2295
rect 10333 2261 10367 2295
rect 10425 2261 10459 2295
rect 10793 2261 10827 2295
rect 11713 2261 11747 2295
rect 11897 2261 11931 2295
rect 12081 2261 12115 2295
rect 12265 2261 12299 2295
rect 12633 2261 12667 2295
<< metal1 >>
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 14458 18000 14464 18012
rect 4120 17972 14464 18000
rect 4120 17960 4126 17972
rect 14458 17960 14464 17972
rect 14516 17960 14522 18012
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 11238 17864 11244 17876
rect 6052 17836 11244 17864
rect 6052 17824 6058 17836
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 14550 17796 14556 17808
rect 4120 17768 14556 17796
rect 4120 17756 4126 17768
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 12894 17728 12900 17740
rect 2746 17700 12900 17728
rect 1026 17484 1032 17536
rect 1084 17524 1090 17536
rect 2746 17524 2774 17700
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 13354 17660 13360 17672
rect 6236 17632 13360 17660
rect 6236 17620 6242 17632
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 14642 17592 14648 17604
rect 10928 17564 14648 17592
rect 10928 17552 10934 17564
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 1084 17496 2774 17524
rect 1084 17484 1090 17496
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 12986 17524 12992 17536
rect 8444 17496 12992 17524
rect 8444 17484 8450 17496
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 6914 17320 6920 17332
rect 6875 17292 6920 17320
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7193 17323 7251 17329
rect 7193 17289 7205 17323
rect 7239 17289 7251 17323
rect 7193 17283 7251 17289
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 7208 17252 7236 17283
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 8481 17323 8539 17329
rect 8481 17320 8493 17323
rect 7340 17292 8493 17320
rect 7340 17280 7346 17292
rect 8481 17289 8493 17292
rect 8527 17289 8539 17323
rect 8481 17283 8539 17289
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 9824 17292 11529 17320
rect 9824 17280 9830 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 12710 17320 12716 17332
rect 12483 17292 12716 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 12986 17320 12992 17332
rect 12947 17292 12992 17320
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 6604 17224 7236 17252
rect 6604 17212 6610 17224
rect 7742 17212 7748 17264
rect 7800 17252 7806 17264
rect 8021 17255 8079 17261
rect 8021 17252 8033 17255
rect 7800 17224 8033 17252
rect 7800 17212 7806 17224
rect 8021 17221 8033 17224
rect 8067 17252 8079 17255
rect 10413 17255 10471 17261
rect 10413 17252 10425 17255
rect 8067 17224 10425 17252
rect 8067 17221 8079 17224
rect 8021 17215 8079 17221
rect 10413 17221 10425 17224
rect 10459 17252 10471 17255
rect 10870 17252 10876 17264
rect 10459 17224 10876 17252
rect 10459 17221 10471 17224
rect 10413 17215 10471 17221
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 11977 17255 12035 17261
rect 11977 17252 11989 17255
rect 11348 17224 11989 17252
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 5592 17156 6469 17184
rect 5592 17144 5598 17156
rect 6457 17153 6469 17156
rect 6503 17184 6515 17187
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6503 17156 6745 17184
rect 6503 17153 6515 17156
rect 6457 17147 6515 17153
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17184 7987 17187
rect 8570 17184 8576 17196
rect 7975 17156 8576 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 4304 17088 6653 17116
rect 4304 17076 4310 17088
rect 6641 17085 6653 17088
rect 6687 17116 6699 17119
rect 7392 17116 7420 17147
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17184 8723 17187
rect 10321 17187 10379 17193
rect 8711 17156 9260 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 8202 17116 8208 17128
rect 6687 17088 7420 17116
rect 8163 17088 8208 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9232 17125 9260 17156
rect 10321 17153 10333 17187
rect 10367 17184 10379 17187
rect 10778 17184 10784 17196
rect 10367 17156 10784 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11348 17193 11376 17224
rect 11977 17221 11989 17224
rect 12023 17252 12035 17255
rect 12023 17224 12756 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9263 17088 9597 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 9585 17085 9597 17088
rect 9631 17116 9643 17119
rect 9766 17116 9772 17128
rect 9631 17088 9772 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17116 10655 17119
rect 10870 17116 10876 17128
rect 10643 17088 10876 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12526 17116 12532 17128
rect 12487 17088 12532 17116
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 7708 17020 11161 17048
rect 7708 17008 7714 17020
rect 11149 17017 11161 17020
rect 11195 17017 11207 17051
rect 11149 17011 11207 17017
rect 11790 17008 11796 17060
rect 11848 17048 11854 17060
rect 12636 17048 12664 17079
rect 11848 17020 12664 17048
rect 12728 17048 12756 17224
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 13446 17252 13452 17264
rect 12860 17224 13452 17252
rect 12860 17212 12866 17224
rect 13446 17212 13452 17224
rect 13504 17252 13510 17264
rect 13633 17255 13691 17261
rect 13633 17252 13645 17255
rect 13504 17224 13645 17252
rect 13504 17212 13510 17224
rect 13633 17221 13645 17224
rect 13679 17221 13691 17255
rect 13633 17215 13691 17221
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17153 13231 17187
rect 13538 17184 13544 17196
rect 13499 17156 13544 17184
rect 13173 17147 13231 17153
rect 13188 17116 13216 17147
rect 13538 17144 13544 17156
rect 13596 17184 13602 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 13596 17156 14473 17184
rect 13596 17144 13602 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 13188 17088 13676 17116
rect 13648 17060 13676 17088
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17116 13967 17119
rect 15378 17116 15384 17128
rect 13955 17088 15384 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 15378 17076 15384 17088
rect 15436 17076 15442 17128
rect 12728 17020 13584 17048
rect 11848 17008 11854 17020
rect 4430 16980 4436 16992
rect 4391 16952 4436 16980
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 4764 16952 4813 16980
rect 4764 16940 4770 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 4801 16943 4859 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16980 5687 16983
rect 5718 16980 5724 16992
rect 5675 16952 5724 16980
rect 5675 16949 5687 16952
rect 5629 16943 5687 16949
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 5994 16980 6000 16992
rect 5955 16952 6000 16980
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 7558 16980 7564 16992
rect 7519 16952 7564 16980
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 7926 16940 7932 16992
rect 7984 16980 7990 16992
rect 8941 16983 8999 16989
rect 8941 16980 8953 16983
rect 7984 16952 8953 16980
rect 7984 16940 7990 16952
rect 8941 16949 8953 16952
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 9272 16952 9321 16980
rect 9272 16940 9278 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 9582 16940 9588 16992
rect 9640 16980 9646 16992
rect 9677 16983 9735 16989
rect 9677 16980 9689 16983
rect 9640 16952 9689 16980
rect 9640 16940 9646 16952
rect 9677 16949 9689 16952
rect 9723 16949 9735 16983
rect 9950 16980 9956 16992
rect 9911 16952 9956 16980
rect 9677 16943 9735 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 12032 16952 12081 16980
rect 12032 16940 12038 16952
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 12069 16943 12127 16949
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 13170 16980 13176 16992
rect 12676 16952 13176 16980
rect 12676 16940 12682 16952
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 13556 16980 13584 17020
rect 13630 17008 13636 17060
rect 13688 17048 13694 17060
rect 14093 17051 14151 17057
rect 14093 17048 14105 17051
rect 13688 17020 14105 17048
rect 13688 17008 13694 17020
rect 14093 17017 14105 17020
rect 14139 17048 14151 17051
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 14139 17020 14289 17048
rect 14139 17017 14151 17020
rect 14093 17011 14151 17017
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 14277 17011 14335 17017
rect 14918 16980 14924 16992
rect 13556 16952 14924 16980
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3145 16779 3203 16785
rect 3145 16776 3157 16779
rect 3016 16748 3157 16776
rect 3016 16736 3022 16748
rect 3145 16745 3157 16748
rect 3191 16776 3203 16779
rect 3694 16776 3700 16788
rect 3191 16748 3700 16776
rect 3191 16745 3203 16748
rect 3145 16739 3203 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4706 16736 4712 16788
rect 4764 16776 4770 16788
rect 5166 16776 5172 16788
rect 4764 16748 5172 16776
rect 4764 16736 4770 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 7653 16779 7711 16785
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 7742 16776 7748 16788
rect 7699 16748 7748 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 11146 16776 11152 16788
rect 7984 16748 11152 16776
rect 7984 16736 7990 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12584 16748 13093 16776
rect 12584 16736 12590 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 2884 16680 4844 16708
rect 1762 16572 1768 16584
rect 1723 16544 1768 16572
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16572 2651 16575
rect 2884 16572 2912 16680
rect 3252 16612 3556 16640
rect 2639 16544 2912 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3016 16544 3061 16572
rect 3016 16532 3022 16544
rect 3142 16532 3148 16584
rect 3200 16572 3206 16584
rect 3252 16572 3280 16612
rect 3200 16544 3280 16572
rect 3200 16532 3206 16544
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 3528 16572 3556 16612
rect 4341 16575 4399 16581
rect 3384 16544 3429 16572
rect 3528 16544 4292 16572
rect 3384 16532 3390 16544
rect 3234 16464 3240 16516
rect 3292 16504 3298 16516
rect 4264 16504 4292 16544
rect 4341 16541 4353 16575
rect 4387 16572 4399 16575
rect 4430 16572 4436 16584
rect 4387 16544 4436 16572
rect 4387 16541 4399 16544
rect 4341 16535 4399 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4706 16572 4712 16584
rect 4667 16544 4712 16572
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 4816 16572 4844 16680
rect 6270 16668 6276 16720
rect 6328 16708 6334 16720
rect 9766 16708 9772 16720
rect 6328 16680 7328 16708
rect 6328 16668 6334 16680
rect 5718 16640 5724 16652
rect 5460 16612 5724 16640
rect 5077 16575 5135 16581
rect 4816 16544 5028 16572
rect 5000 16504 5028 16544
rect 5077 16541 5089 16575
rect 5123 16572 5135 16575
rect 5258 16572 5264 16584
rect 5123 16544 5264 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5460 16581 5488 16612
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 7006 16640 7012 16652
rect 6595 16612 7012 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7300 16649 7328 16680
rect 8404 16680 9772 16708
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8260 16612 8309 16640
rect 8260 16600 8266 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16541 5503 16575
rect 5445 16535 5503 16541
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16572 5871 16575
rect 5994 16572 6000 16584
rect 5859 16544 6000 16572
rect 5859 16541 5871 16544
rect 5813 16535 5871 16541
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7558 16572 7564 16584
rect 7147 16544 7564 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8404 16572 8432 16680
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 11698 16708 11704 16720
rect 10980 16680 11704 16708
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 10980 16649 11008 16680
rect 11698 16668 11704 16680
rect 11756 16708 11762 16720
rect 12618 16708 12624 16720
rect 11756 16680 12624 16708
rect 11756 16668 11762 16680
rect 12618 16668 12624 16680
rect 12676 16668 12682 16720
rect 12820 16680 13676 16708
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 9456 16612 10241 16640
rect 9456 16600 9462 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 11790 16640 11796 16652
rect 11655 16612 11796 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 8570 16572 8576 16584
rect 8159 16544 8432 16572
rect 8531 16544 8576 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 9214 16572 9220 16584
rect 9175 16544 9220 16572
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 9582 16572 9588 16584
rect 9543 16544 9588 16572
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9950 16532 9956 16584
rect 10008 16572 10014 16584
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 10008 16544 10057 16572
rect 10008 16532 10014 16544
rect 10045 16541 10057 16544
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11072 16572 11100 16603
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12820 16649 12848 16680
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12584 16612 12817 16640
rect 12584 16600 12590 16612
rect 12805 16609 12817 16612
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 13648 16649 13676 16680
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13504 16612 13553 16640
rect 13504 16600 13510 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 14458 16640 14464 16652
rect 14419 16612 14464 16640
rect 13633 16603 13691 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 10928 16544 11100 16572
rect 10928 16532 10934 16544
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 12434 16572 12440 16584
rect 11204 16544 12440 16572
rect 11204 16532 11210 16544
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 13814 16572 13820 16584
rect 12676 16544 13820 16572
rect 12676 16532 12682 16544
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 6273 16507 6331 16513
rect 3292 16476 4200 16504
rect 4264 16476 4936 16504
rect 5000 16476 5948 16504
rect 3292 16464 3298 16476
rect 1854 16396 1860 16448
rect 1912 16436 1918 16448
rect 2777 16439 2835 16445
rect 2777 16436 2789 16439
rect 1912 16408 2789 16436
rect 1912 16396 1918 16408
rect 2777 16405 2789 16408
rect 2823 16405 2835 16439
rect 2777 16399 2835 16405
rect 3513 16439 3571 16445
rect 3513 16405 3525 16439
rect 3559 16436 3571 16439
rect 3602 16436 3608 16448
rect 3559 16408 3608 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 4172 16445 4200 16476
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16405 4215 16439
rect 4157 16399 4215 16405
rect 4338 16396 4344 16448
rect 4396 16436 4402 16448
rect 4908 16445 4936 16476
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4396 16408 4537 16436
rect 4396 16396 4402 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 4893 16439 4951 16445
rect 4893 16405 4905 16439
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 5132 16408 5273 16436
rect 5132 16396 5138 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 5629 16439 5687 16445
rect 5629 16405 5641 16439
rect 5675 16436 5687 16439
rect 5810 16436 5816 16448
rect 5675 16408 5816 16436
rect 5675 16405 5687 16408
rect 5629 16399 5687 16405
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 5920 16445 5948 16476
rect 6273 16473 6285 16507
rect 6319 16504 6331 16507
rect 7193 16507 7251 16513
rect 6319 16476 6776 16504
rect 6319 16473 6331 16476
rect 6273 16467 6331 16473
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16405 5963 16439
rect 5905 16399 5963 16405
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 6748 16445 6776 16476
rect 7193 16473 7205 16507
rect 7239 16504 7251 16507
rect 7239 16476 7788 16504
rect 7239 16473 7251 16476
rect 7193 16467 7251 16473
rect 7760 16445 7788 16476
rect 8018 16464 8024 16516
rect 8076 16504 8082 16516
rect 8076 16476 9076 16504
rect 8076 16464 8082 16476
rect 6733 16439 6791 16445
rect 6420 16408 6465 16436
rect 6420 16396 6426 16408
rect 6733 16405 6745 16439
rect 6779 16405 6791 16439
rect 6733 16399 6791 16405
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16405 7803 16439
rect 7745 16399 7803 16405
rect 7926 16396 7932 16448
rect 7984 16436 7990 16448
rect 9048 16445 9076 16476
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 11793 16507 11851 16513
rect 9824 16476 10916 16504
rect 9824 16464 9830 16476
rect 8205 16439 8263 16445
rect 8205 16436 8217 16439
rect 7984 16408 8217 16436
rect 7984 16396 7990 16408
rect 8205 16405 8217 16408
rect 8251 16405 8263 16439
rect 8205 16399 8263 16405
rect 9033 16439 9091 16445
rect 9033 16405 9045 16439
rect 9079 16405 9091 16439
rect 9033 16399 9091 16405
rect 9306 16396 9312 16448
rect 9364 16436 9370 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 9364 16408 9413 16436
rect 9364 16396 9370 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9401 16399 9459 16405
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 10888 16445 10916 16476
rect 11793 16473 11805 16507
rect 11839 16504 11851 16507
rect 12713 16507 12771 16513
rect 11839 16476 12296 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 10137 16439 10195 16445
rect 10137 16405 10149 16439
rect 10183 16436 10195 16439
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10183 16408 10517 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 10505 16399 10563 16405
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16405 10931 16439
rect 11698 16436 11704 16448
rect 11659 16408 11704 16436
rect 10873 16399 10931 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12268 16445 12296 16476
rect 12713 16473 12725 16507
rect 12759 16504 12771 16507
rect 12802 16504 12808 16516
rect 12759 16476 12808 16504
rect 12759 16473 12771 16476
rect 12713 16467 12771 16473
rect 12802 16464 12808 16476
rect 12860 16504 12866 16516
rect 14553 16507 14611 16513
rect 12860 16476 14228 16504
rect 12860 16464 12866 16476
rect 12161 16439 12219 16445
rect 12161 16436 12173 16439
rect 12032 16408 12173 16436
rect 12032 16396 12038 16408
rect 12161 16405 12173 16408
rect 12207 16405 12219 16439
rect 12161 16399 12219 16405
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 13630 16436 13636 16448
rect 13495 16408 13636 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14200 16445 14228 16476
rect 14553 16473 14565 16507
rect 14599 16504 14611 16507
rect 14826 16504 14832 16516
rect 14599 16476 14832 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 14826 16464 14832 16476
rect 14884 16464 14890 16516
rect 14185 16439 14243 16445
rect 14185 16405 14197 16439
rect 14231 16436 14243 16439
rect 14642 16436 14648 16448
rect 14231 16408 14648 16436
rect 14231 16405 14243 16408
rect 14185 16399 14243 16405
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 2498 16192 2504 16244
rect 2556 16232 2562 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2556 16204 2605 16232
rect 2556 16192 2562 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 2593 16195 2651 16201
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3970 16232 3976 16244
rect 3743 16204 3976 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 4939 16204 5365 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 7466 16232 7472 16244
rect 5859 16204 7472 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9401 16235 9459 16241
rect 9401 16232 9413 16235
rect 9079 16204 9413 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9401 16201 9413 16204
rect 9447 16201 9459 16235
rect 9401 16195 9459 16201
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 9953 16235 10011 16241
rect 9953 16232 9965 16235
rect 9539 16204 9965 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 9953 16201 9965 16204
rect 9999 16201 10011 16235
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 9953 16195 10011 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11146 16232 11152 16244
rect 11107 16204 11152 16232
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 11514 16232 11520 16244
rect 11475 16204 11520 16232
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 11974 16232 11980 16244
rect 11935 16204 11980 16232
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12710 16232 12716 16244
rect 12671 16204 12716 16232
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 13173 16235 13231 16241
rect 13173 16201 13185 16235
rect 13219 16232 13231 16235
rect 13219 16204 14228 16232
rect 13219 16201 13231 16204
rect 13173 16195 13231 16201
rect 3326 16124 3332 16176
rect 3384 16164 3390 16176
rect 3786 16164 3792 16176
rect 3384 16136 3792 16164
rect 3384 16124 3390 16136
rect 3786 16124 3792 16136
rect 3844 16124 3850 16176
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 9306 16164 9312 16176
rect 4672 16136 9312 16164
rect 4672 16124 4678 16136
rect 9306 16124 9312 16136
rect 9364 16124 9370 16176
rect 11348 16136 12434 16164
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16096 2835 16099
rect 3513 16099 3571 16105
rect 2823 16068 3004 16096
rect 2823 16065 2835 16068
rect 2777 16059 2835 16065
rect 1578 15852 1584 15904
rect 1636 15892 1642 15904
rect 1872 15892 1900 16059
rect 2976 15901 3004 16068
rect 3513 16065 3525 16099
rect 3559 16096 3571 16099
rect 3602 16096 3608 16108
rect 3559 16068 3608 16096
rect 3559 16065 3571 16068
rect 3513 16059 3571 16065
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 5718 16096 5724 16108
rect 5679 16068 5724 16096
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 6779 16068 7328 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 15997 5043 16031
rect 5166 16028 5172 16040
rect 5127 16000 5172 16028
rect 4985 15991 5043 15997
rect 5000 15960 5028 15991
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 5902 15988 5908 16040
rect 5960 16028 5966 16040
rect 5997 16031 6055 16037
rect 5997 16028 6009 16031
rect 5960 16000 6009 16028
rect 5960 15988 5966 16000
rect 5997 15997 6009 16000
rect 6043 16028 6055 16031
rect 6822 16028 6828 16040
rect 6043 16000 6500 16028
rect 6783 16000 6828 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 6365 15963 6423 15969
rect 6365 15960 6377 15963
rect 5000 15932 6377 15960
rect 6365 15929 6377 15932
rect 6411 15929 6423 15963
rect 6472 15960 6500 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 6932 15960 6960 15991
rect 7300 15969 7328 16068
rect 7374 16056 7380 16108
rect 7432 16096 7438 16108
rect 7926 16096 7932 16108
rect 7432 16068 7932 16096
rect 7432 16056 7438 16068
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 8938 16096 8944 16108
rect 8711 16068 8944 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16096 10379 16099
rect 11238 16096 11244 16108
rect 10367 16068 11244 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11348 16105 11376 16136
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11882 16096 11888 16108
rect 11843 16068 11888 16096
rect 11333 16059 11391 16065
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12406 16096 12434 16136
rect 12526 16124 12532 16176
rect 12584 16164 12590 16176
rect 12584 16136 13308 16164
rect 12584 16124 12590 16136
rect 12618 16096 12624 16108
rect 12406 16068 12624 16096
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13078 16096 13084 16108
rect 13039 16068 13084 16096
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 7650 15988 7656 16040
rect 7708 16028 7714 16040
rect 8110 16028 8116 16040
rect 7708 16000 8116 16028
rect 7708 15988 7714 16000
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8846 16028 8852 16040
rect 8619 16000 8852 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 16028 9367 16031
rect 9398 16028 9404 16040
rect 9355 16000 9404 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 10284 16000 10425 16028
rect 10284 15988 10290 16000
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 10870 16028 10876 16040
rect 10551 16000 10876 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 6472 15932 6960 15960
rect 7285 15963 7343 15969
rect 6365 15923 6423 15929
rect 7285 15929 7297 15963
rect 7331 15960 7343 15963
rect 9214 15960 9220 15972
rect 7331 15932 9220 15960
rect 7331 15929 7343 15932
rect 7285 15923 7343 15929
rect 9214 15920 9220 15932
rect 9272 15920 9278 15972
rect 10520 15960 10548 15991
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 13280 16037 13308 16136
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13412 16068 13921 16096
rect 13412 16056 13418 16068
rect 13909 16065 13921 16068
rect 13955 16065 13967 16099
rect 13909 16059 13967 16065
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11480 16000 12081 16028
rect 11480 15988 11486 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 13265 16031 13323 16037
rect 13265 15997 13277 16031
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 12802 15960 12808 15972
rect 9784 15932 10548 15960
rect 10612 15932 12808 15960
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1636 15864 1961 15892
rect 1636 15852 1642 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 1949 15855 2007 15861
rect 2961 15895 3019 15901
rect 2961 15861 2973 15895
rect 3007 15892 3019 15895
rect 3418 15892 3424 15904
rect 3007 15864 3424 15892
rect 3007 15861 3019 15864
rect 2961 15855 3019 15861
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 3602 15852 3608 15904
rect 3660 15892 3666 15904
rect 3881 15895 3939 15901
rect 3881 15892 3893 15895
rect 3660 15864 3893 15892
rect 3660 15852 3666 15864
rect 3881 15861 3893 15864
rect 3927 15861 3939 15895
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 3881 15855 3939 15861
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7190 15892 7196 15904
rect 6972 15864 7196 15892
rect 6972 15852 6978 15864
rect 7190 15852 7196 15864
rect 7248 15892 7254 15904
rect 7374 15892 7380 15904
rect 7248 15864 7380 15892
rect 7248 15852 7254 15864
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 7561 15895 7619 15901
rect 7561 15892 7573 15895
rect 7524 15864 7573 15892
rect 7524 15852 7530 15864
rect 7561 15861 7573 15864
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 7834 15852 7840 15904
rect 7892 15892 7898 15904
rect 7929 15895 7987 15901
rect 7929 15892 7941 15895
rect 7892 15864 7941 15892
rect 7892 15852 7898 15864
rect 7929 15861 7941 15864
rect 7975 15861 7987 15895
rect 7929 15855 7987 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9784 15892 9812 15932
rect 8444 15864 9812 15892
rect 9861 15895 9919 15901
rect 8444 15852 8450 15864
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 9950 15892 9956 15904
rect 9907 15864 9956 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10612 15892 10640 15932
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 12894 15920 12900 15972
rect 12952 15960 12958 15972
rect 13541 15963 13599 15969
rect 13541 15960 13553 15963
rect 12952 15932 13553 15960
rect 12952 15920 12958 15932
rect 13541 15929 13553 15932
rect 13587 15929 13599 15963
rect 14200 15960 14228 16204
rect 14458 16192 14464 16244
rect 14516 16232 14522 16244
rect 14553 16235 14611 16241
rect 14553 16232 14565 16235
rect 14516 16204 14565 16232
rect 14516 16192 14522 16204
rect 14553 16201 14565 16204
rect 14599 16201 14611 16235
rect 14553 16195 14611 16201
rect 15381 16167 15439 16173
rect 15381 16133 15393 16167
rect 15427 16164 15439 16167
rect 16114 16164 16120 16176
rect 15427 16136 16120 16164
rect 15427 16133 15439 16136
rect 15381 16127 15439 16133
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 15010 16056 15016 16108
rect 15068 16096 15074 16108
rect 15105 16099 15163 16105
rect 15105 16096 15117 16099
rect 15068 16068 15117 16096
rect 15068 16056 15074 16068
rect 15105 16065 15117 16068
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 14826 16028 14832 16040
rect 14323 16000 14832 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 14461 15963 14519 15969
rect 14461 15960 14473 15963
rect 14200 15932 14473 15960
rect 13541 15923 13599 15929
rect 14461 15929 14473 15932
rect 14507 15960 14519 15963
rect 15746 15960 15752 15972
rect 14507 15932 15752 15960
rect 14507 15929 14519 15932
rect 14461 15923 14519 15929
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 10100 15864 10640 15892
rect 10100 15852 10106 15864
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 15010 15892 15016 15904
rect 12492 15864 12537 15892
rect 14971 15864 15016 15892
rect 12492 15852 12498 15864
rect 15010 15852 15016 15864
rect 15068 15852 15074 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 2130 15648 2136 15700
rect 2188 15688 2194 15700
rect 2593 15691 2651 15697
rect 2593 15688 2605 15691
rect 2188 15660 2605 15688
rect 2188 15648 2194 15660
rect 2593 15657 2605 15660
rect 2639 15657 2651 15691
rect 6178 15688 6184 15700
rect 2593 15651 2651 15657
rect 2746 15660 6184 15688
rect 1578 15580 1584 15632
rect 1636 15620 1642 15632
rect 2746 15620 2774 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6362 15688 6368 15700
rect 6323 15660 6368 15688
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 7742 15688 7748 15700
rect 6656 15660 7748 15688
rect 4062 15620 4068 15632
rect 1636 15592 2774 15620
rect 4023 15592 4068 15620
rect 1636 15580 1642 15592
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 6656 15620 6684 15660
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8938 15688 8944 15700
rect 8899 15660 8944 15688
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 11020 15660 11253 15688
rect 11020 15648 11026 15660
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 11241 15651 11299 15657
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 11756 15660 11897 15688
rect 11756 15648 11762 15660
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12952 15660 13461 15688
rect 12952 15648 12958 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 4816 15592 6684 15620
rect 6748 15592 8033 15620
rect 3326 15552 3332 15564
rect 3287 15524 3332 15552
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3878 15512 3884 15564
rect 3936 15552 3942 15564
rect 4816 15561 4844 15592
rect 4801 15555 4859 15561
rect 3936 15524 4752 15552
rect 3936 15512 3942 15524
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 3605 15487 3663 15493
rect 2832 15456 2877 15484
rect 2832 15444 2838 15456
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 4522 15484 4528 15496
rect 3651 15456 4200 15484
rect 4483 15456 4528 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 4062 15416 4068 15428
rect 1452 15388 4068 15416
rect 1452 15376 1458 15388
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2832 15320 2973 15348
rect 2832 15308 2838 15320
rect 2961 15317 2973 15320
rect 3007 15348 3019 15351
rect 3878 15348 3884 15360
rect 3007 15320 3884 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 4172 15357 4200 15456
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4724 15484 4752 15524
rect 4801 15521 4813 15555
rect 4847 15521 4859 15555
rect 5626 15552 5632 15564
rect 4801 15515 4859 15521
rect 5184 15524 5632 15552
rect 5184 15484 5212 15524
rect 5626 15512 5632 15524
rect 5684 15512 5690 15564
rect 5718 15512 5724 15564
rect 5776 15552 5782 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5776 15524 5917 15552
rect 5776 15512 5782 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 4724 15456 5212 15484
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 6362 15484 6368 15496
rect 5316 15456 6368 15484
rect 5316 15444 5322 15456
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6748 15493 6776 15592
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 11514 15620 11520 15632
rect 10744 15592 11520 15620
rect 10744 15580 10750 15592
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 12802 15620 12808 15632
rect 11624 15592 12808 15620
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 6840 15524 6929 15552
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 4430 15376 4436 15428
rect 4488 15416 4494 15428
rect 5350 15416 5356 15428
rect 4488 15388 5356 15416
rect 4488 15376 4494 15388
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 6270 15376 6276 15428
rect 6328 15416 6334 15428
rect 6840 15416 6868 15524
rect 6917 15521 6929 15524
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7392 15484 7420 15515
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 8202 15552 8208 15564
rect 7616 15524 8208 15552
rect 7616 15512 7622 15524
rect 8202 15512 8208 15524
rect 8260 15552 8266 15564
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 8260 15524 8585 15552
rect 8260 15512 8266 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 9306 15512 9312 15564
rect 9364 15552 9370 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9364 15524 9505 15552
rect 9364 15512 9370 15524
rect 9493 15521 9505 15524
rect 9539 15552 9551 15555
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 9539 15524 10793 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 8018 15484 8024 15496
rect 7392 15456 8024 15484
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8386 15444 8392 15496
rect 8444 15484 8450 15496
rect 8938 15484 8944 15496
rect 8444 15456 8944 15484
rect 8444 15444 8450 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9401 15487 9459 15493
rect 9401 15484 9413 15487
rect 9180 15456 9413 15484
rect 9180 15444 9186 15456
rect 9401 15453 9413 15456
rect 9447 15484 9459 15487
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9447 15456 9781 15484
rect 9447 15453 9459 15456
rect 9401 15447 9459 15453
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 10686 15484 10692 15496
rect 10643 15456 10692 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10686 15444 10692 15456
rect 10744 15484 10750 15496
rect 10962 15484 10968 15496
rect 10744 15456 10968 15484
rect 10744 15444 10750 15456
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 6328 15388 6868 15416
rect 6328 15376 6334 15388
rect 6914 15376 6920 15428
rect 6972 15416 6978 15428
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 6972 15388 7481 15416
rect 6972 15376 6978 15388
rect 7469 15385 7481 15388
rect 7515 15416 7527 15419
rect 7834 15416 7840 15428
rect 7515 15388 7840 15416
rect 7515 15385 7527 15388
rect 7469 15379 7527 15385
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 8481 15419 8539 15425
rect 8481 15416 8493 15419
rect 7944 15388 8493 15416
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15317 4215 15351
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4157 15311 4215 15317
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5077 15351 5135 15357
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 5442 15348 5448 15360
rect 5123 15320 5448 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 5684 15320 6193 15348
rect 5684 15308 5690 15320
rect 6181 15317 6193 15320
rect 6227 15317 6239 15351
rect 6181 15311 6239 15317
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 7561 15351 7619 15357
rect 6880 15320 6925 15348
rect 6880 15308 6886 15320
rect 7561 15317 7573 15351
rect 7607 15348 7619 15351
rect 7650 15348 7656 15360
rect 7607 15320 7656 15348
rect 7607 15317 7619 15320
rect 7561 15311 7619 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 7944 15357 7972 15388
rect 8481 15385 8493 15388
rect 8527 15385 8539 15419
rect 8481 15379 8539 15385
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 11624 15416 11652 15592
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 13136 15524 13185 15552
rect 13136 15512 13142 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12434 15484 12440 15496
rect 12299 15456 12440 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 12434 15444 12440 15456
rect 12492 15484 12498 15496
rect 12492 15456 14780 15484
rect 12492 15444 12498 15456
rect 9272 15388 11652 15416
rect 11793 15419 11851 15425
rect 9272 15376 9278 15388
rect 11793 15385 11805 15419
rect 11839 15416 11851 15419
rect 11839 15388 12020 15416
rect 11839 15385 11851 15388
rect 11793 15379 11851 15385
rect 7929 15351 7987 15357
rect 7929 15317 7941 15351
rect 7975 15317 7987 15351
rect 7929 15311 7987 15317
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 8352 15320 8401 15348
rect 8352 15308 8358 15320
rect 8389 15317 8401 15320
rect 8435 15317 8447 15351
rect 8389 15311 8447 15317
rect 9309 15351 9367 15357
rect 9309 15317 9321 15351
rect 9355 15348 9367 15351
rect 9490 15348 9496 15360
rect 9355 15320 9496 15348
rect 9355 15317 9367 15320
rect 9309 15311 9367 15317
rect 9490 15308 9496 15320
rect 9548 15348 9554 15360
rect 9953 15351 10011 15357
rect 9953 15348 9965 15351
rect 9548 15320 9965 15348
rect 9548 15308 9554 15320
rect 9953 15317 9965 15320
rect 9999 15317 10011 15351
rect 9953 15311 10011 15317
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 10652 15320 10701 15348
rect 10652 15308 10658 15320
rect 10689 15317 10701 15320
rect 10735 15348 10747 15351
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10735 15320 11069 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 11238 15308 11244 15360
rect 11296 15348 11302 15360
rect 11517 15351 11575 15357
rect 11517 15348 11529 15351
rect 11296 15320 11529 15348
rect 11296 15308 11302 15320
rect 11517 15317 11529 15320
rect 11563 15348 11575 15351
rect 11882 15348 11888 15360
rect 11563 15320 11888 15348
rect 11563 15317 11575 15320
rect 11517 15311 11575 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 11992 15348 12020 15388
rect 12066 15376 12072 15428
rect 12124 15416 12130 15428
rect 12345 15419 12403 15425
rect 12345 15416 12357 15419
rect 12124 15388 12357 15416
rect 12124 15376 12130 15388
rect 12345 15385 12357 15388
rect 12391 15385 12403 15419
rect 12345 15379 12403 15385
rect 12618 15348 12624 15360
rect 11992 15320 12624 15348
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13596 15320 14105 15348
rect 13596 15308 13602 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14553 15351 14611 15357
rect 14553 15317 14565 15351
rect 14599 15348 14611 15351
rect 14642 15348 14648 15360
rect 14599 15320 14648 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 14752 15357 14780 15456
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 15194 15348 15200 15360
rect 14783 15320 15200 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 3605 15147 3663 15153
rect 3605 15113 3617 15147
rect 3651 15144 3663 15147
rect 3970 15144 3976 15156
rect 3651 15116 3976 15144
rect 3651 15113 3663 15116
rect 3605 15107 3663 15113
rect 3970 15104 3976 15116
rect 4028 15104 4034 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 4157 15147 4215 15153
rect 4157 15144 4169 15147
rect 4120 15116 4169 15144
rect 4120 15104 4126 15116
rect 4157 15113 4169 15116
rect 4203 15113 4215 15147
rect 4157 15107 4215 15113
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 4614 15144 4620 15156
rect 4479 15116 4620 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 4939 15116 5273 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 5626 15144 5632 15156
rect 5587 15116 5632 15144
rect 5261 15107 5319 15113
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 6549 15147 6607 15153
rect 6549 15113 6561 15147
rect 6595 15144 6607 15147
rect 6822 15144 6828 15156
rect 6595 15116 6828 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 7055 15116 7389 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 8665 15147 8723 15153
rect 7791 15116 8432 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 8404 15088 8432 15116
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8846 15144 8852 15156
rect 8711 15116 8852 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9030 15144 9036 15156
rect 8991 15116 9036 15144
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9732 15116 9873 15144
rect 9732 15104 9738 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 9861 15107 9919 15113
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 11241 15147 11299 15153
rect 10008 15116 10053 15144
rect 10008 15104 10014 15116
rect 11241 15113 11253 15147
rect 11287 15144 11299 15147
rect 11330 15144 11336 15156
rect 11287 15116 11336 15144
rect 11287 15113 11299 15116
rect 11241 15107 11299 15113
rect 11330 15104 11336 15116
rect 11388 15144 11394 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11388 15116 11897 15144
rect 11388 15104 11394 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12345 15147 12403 15153
rect 12345 15144 12357 15147
rect 12124 15116 12357 15144
rect 12124 15104 12130 15116
rect 12345 15113 12357 15116
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15144 12863 15147
rect 14274 15144 14280 15156
rect 12851 15116 14280 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14369 15147 14427 15153
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 14829 15147 14887 15153
rect 14829 15144 14841 15147
rect 14415 15116 14841 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 14829 15113 14841 15116
rect 14875 15113 14887 15147
rect 14829 15107 14887 15113
rect 5442 15076 5448 15088
rect 4356 15048 5448 15076
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 3510 15008 3516 15020
rect 3471 14980 3516 15008
rect 2041 14971 2099 14977
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2056 14872 2084 14971
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 4356 15017 4384 15048
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 5810 15036 5816 15088
rect 5868 15076 5874 15088
rect 6457 15079 6515 15085
rect 6457 15076 6469 15079
rect 5868 15048 6469 15076
rect 5868 15036 5874 15048
rect 6457 15045 6469 15048
rect 6503 15076 6515 15079
rect 8202 15076 8208 15088
rect 6503 15048 8208 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 8386 15036 8392 15088
rect 8444 15076 8450 15088
rect 9048 15076 9076 15104
rect 10321 15079 10379 15085
rect 10321 15076 10333 15079
rect 8444 15048 10333 15076
rect 8444 15036 8450 15048
rect 10321 15045 10333 15048
rect 10367 15045 10379 15079
rect 10321 15039 10379 15045
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11606 15076 11612 15088
rect 11204 15048 11612 15076
rect 11204 15036 11210 15048
rect 11606 15036 11612 15048
rect 11664 15036 11670 15088
rect 11716 15048 15424 15076
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5074 15008 5080 15020
rect 4847 14980 5080 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7282 15008 7288 15020
rect 6963 14980 7288 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 15008 7895 15011
rect 7883 14980 8892 15008
rect 7883 14977 7895 14980
rect 7837 14971 7895 14977
rect 8864 14952 8892 14980
rect 3786 14940 3792 14952
rect 3747 14912 3792 14940
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5166 14940 5172 14952
rect 5031 14912 5172 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5902 14940 5908 14952
rect 5863 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 7558 14940 7564 14952
rect 7239 14912 7564 14940
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 8018 14940 8024 14952
rect 7979 14912 8024 14940
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8846 14900 8852 14952
rect 8904 14940 8910 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8904 14912 9137 14940
rect 8904 14900 8910 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9306 14940 9312 14952
rect 9267 14912 9312 14940
rect 9125 14903 9183 14909
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 10134 14940 10140 14952
rect 10095 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 11716 14949 11744 15048
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 15008 12771 15011
rect 12802 15008 12808 15020
rect 12759 14980 12808 15008
rect 12759 14977 12771 14980
rect 12713 14971 12771 14977
rect 12802 14968 12808 14980
rect 12860 15008 12866 15020
rect 13354 15008 13360 15020
rect 12860 14980 13360 15008
rect 12860 14968 12866 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 14792 14980 15209 15008
rect 14792 14968 14798 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 15197 14971 15255 14977
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 11664 14912 11713 14940
rect 11664 14900 11670 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 9493 14875 9551 14881
rect 9493 14872 9505 14875
rect 2056 14844 9505 14872
rect 9493 14841 9505 14844
rect 9539 14841 9551 14875
rect 11808 14872 11836 14903
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13262 14940 13268 14952
rect 12952 14912 12997 14940
rect 13223 14912 13268 14940
rect 12952 14900 12958 14912
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13449 14903 13507 14909
rect 13740 14912 14105 14940
rect 9493 14835 9551 14841
rect 11072 14844 11836 14872
rect 12253 14875 12311 14881
rect 11072 14816 11100 14844
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 13464 14872 13492 14903
rect 12299 14844 13492 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 3142 14804 3148 14816
rect 3103 14776 3148 14804
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5040 14776 6193 14804
rect 5040 14764 5046 14776
rect 6181 14773 6193 14776
rect 6227 14804 6239 14807
rect 7834 14804 7840 14816
rect 6227 14776 7840 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8573 14807 8631 14813
rect 8573 14773 8585 14807
rect 8619 14804 8631 14807
rect 8846 14804 8852 14816
rect 8619 14776 8852 14804
rect 8619 14773 8631 14776
rect 8573 14767 8631 14773
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 11054 14804 11060 14816
rect 11015 14776 11060 14804
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13740 14804 13768 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 14918 14940 14924 14952
rect 14323 14912 14924 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 15396 14949 15424 15048
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 15470 14940 15476 14952
rect 15427 14912 15476 14940
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 15194 14832 15200 14884
rect 15252 14872 15258 14884
rect 15304 14872 15332 14903
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 15252 14844 15332 14872
rect 15252 14832 15258 14844
rect 13320 14776 13768 14804
rect 13909 14807 13967 14813
rect 13320 14764 13326 14776
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 14458 14804 14464 14816
rect 13955 14776 14464 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14608 14776 14749 14804
rect 14608 14764 14614 14776
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 14737 14767 14795 14773
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 4890 14600 4896 14612
rect 4851 14572 4896 14600
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5074 14600 5080 14612
rect 5035 14572 5080 14600
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 5776 14572 5917 14600
rect 5776 14560 5782 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 7282 14600 7288 14612
rect 7243 14572 7288 14600
rect 5905 14563 5963 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 7892 14572 8401 14600
rect 7892 14560 7898 14572
rect 8389 14569 8401 14572
rect 8435 14600 8447 14603
rect 9490 14600 9496 14612
rect 8435 14572 9496 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 9490 14560 9496 14572
rect 9548 14600 9554 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9548 14572 9965 14600
rect 9548 14560 9554 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 10928 14572 11529 14600
rect 10928 14560 10934 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 14918 14600 14924 14612
rect 14879 14572 14924 14600
rect 11517 14563 11575 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 4709 14535 4767 14541
rect 4709 14501 4721 14535
rect 4755 14532 4767 14535
rect 5258 14532 5264 14544
rect 4755 14504 5264 14532
rect 4755 14501 4767 14504
rect 4709 14495 4767 14501
rect 1670 14464 1676 14476
rect 1631 14436 1676 14464
rect 1670 14424 1676 14436
rect 1728 14424 1734 14476
rect 2682 14424 2688 14476
rect 2740 14464 2746 14476
rect 2869 14467 2927 14473
rect 2869 14464 2881 14467
rect 2740 14436 2881 14464
rect 2740 14424 2746 14436
rect 2869 14433 2881 14436
rect 2915 14433 2927 14467
rect 2869 14427 2927 14433
rect 3142 14424 3148 14476
rect 3200 14424 3206 14476
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 3844 14436 4353 14464
rect 3844 14424 3850 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2590 14396 2596 14408
rect 1995 14368 2596 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 3160 14396 3188 14424
rect 2976 14368 3188 14396
rect 4157 14399 4215 14405
rect 2976 14260 3004 14368
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4724 14396 4752 14495
rect 5258 14492 5264 14504
rect 5316 14532 5322 14544
rect 5534 14532 5540 14544
rect 5316 14504 5540 14532
rect 5316 14492 5322 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 8113 14535 8171 14541
rect 8113 14532 8125 14535
rect 5684 14504 8125 14532
rect 5684 14492 5690 14504
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14464 5779 14467
rect 5902 14464 5908 14476
rect 5767 14436 5908 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6454 14464 6460 14476
rect 6415 14436 6460 14464
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 7760 14473 7788 14504
rect 8113 14501 8125 14504
rect 8159 14532 8171 14535
rect 9122 14532 9128 14544
rect 8159 14504 9128 14532
rect 8159 14501 8171 14504
rect 8113 14495 8171 14501
rect 9122 14492 9128 14504
rect 9180 14532 9186 14544
rect 9769 14535 9827 14541
rect 9769 14532 9781 14535
rect 9180 14504 9781 14532
rect 9180 14492 9186 14504
rect 9769 14501 9781 14504
rect 9815 14501 9827 14535
rect 9769 14495 9827 14501
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8018 14464 8024 14476
rect 7975 14436 8024 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8018 14424 8024 14436
rect 8076 14464 8082 14476
rect 9030 14464 9036 14476
rect 8076 14436 9036 14464
rect 8076 14424 8082 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 14550 14464 14556 14476
rect 14511 14436 14556 14464
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 14645 14467 14703 14473
rect 14645 14433 14657 14467
rect 14691 14433 14703 14467
rect 15470 14464 15476 14476
rect 15431 14436 15476 14464
rect 14645 14427 14703 14433
rect 4203 14368 4752 14396
rect 5445 14399 5503 14405
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 5445 14365 5457 14399
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 3053 14331 3111 14337
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 5460 14328 5488 14359
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 7653 14399 7711 14405
rect 5592 14368 6408 14396
rect 5592 14356 5598 14368
rect 5810 14328 5816 14340
rect 3099 14300 3832 14328
rect 5460 14300 5816 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 3145 14263 3203 14269
rect 3145 14260 3157 14263
rect 2976 14232 3157 14260
rect 3145 14229 3157 14232
rect 3191 14229 3203 14263
rect 3145 14223 3203 14229
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 3804 14269 3832 14300
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 6380 14337 6408 14368
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7834 14396 7840 14408
rect 7699 14368 7840 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8168 14368 8953 14396
rect 8168 14356 8174 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14396 11299 14399
rect 11330 14396 11336 14408
rect 11287 14368 11336 14396
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 11330 14356 11336 14368
rect 11388 14396 11394 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11388 14368 11437 14396
rect 11388 14356 11394 14368
rect 11425 14365 11437 14368
rect 11471 14396 11483 14399
rect 13170 14396 13176 14408
rect 11471 14368 13176 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 14458 14396 14464 14408
rect 14419 14368 14464 14396
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 12986 14337 12992 14340
rect 6365 14331 6423 14337
rect 6365 14297 6377 14331
rect 6411 14328 6423 14331
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 6411 14300 6837 14328
rect 6411 14297 6423 14300
rect 6365 14291 6423 14297
rect 6825 14297 6837 14300
rect 6871 14328 6883 14331
rect 12928 14331 12992 14337
rect 12928 14328 12940 14331
rect 6871 14300 8616 14328
rect 12899 14300 12940 14328
rect 6871 14297 6883 14300
rect 6825 14291 6883 14297
rect 3513 14263 3571 14269
rect 3513 14260 3525 14263
rect 3292 14232 3525 14260
rect 3292 14220 3298 14232
rect 3513 14229 3525 14232
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4212 14232 4261 14260
rect 4212 14220 4218 14232
rect 4249 14229 4261 14232
rect 4295 14260 4307 14263
rect 4890 14260 4896 14272
rect 4295 14232 4896 14260
rect 4295 14229 4307 14232
rect 4249 14223 4307 14229
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 5040 14232 5549 14260
rect 5040 14220 5046 14232
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 5537 14223 5595 14229
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 6273 14263 6331 14269
rect 6273 14260 6285 14263
rect 5684 14232 6285 14260
rect 5684 14220 5690 14232
rect 6273 14229 6285 14232
rect 6319 14260 6331 14263
rect 6730 14260 6736 14272
rect 6319 14232 6736 14260
rect 6319 14229 6331 14232
rect 6273 14223 6331 14229
rect 6730 14220 6736 14232
rect 6788 14260 6794 14272
rect 8588 14269 8616 14300
rect 12928 14297 12940 14300
rect 12974 14297 12992 14331
rect 12928 14291 12992 14297
rect 12986 14288 12992 14291
rect 13044 14328 13050 14340
rect 13906 14328 13912 14340
rect 13044 14300 13912 14328
rect 13044 14288 13050 14300
rect 13906 14288 13912 14300
rect 13964 14328 13970 14340
rect 14660 14328 14688 14427
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15381 14331 15439 14337
rect 15381 14328 15393 14331
rect 13964 14300 14688 14328
rect 14752 14300 15393 14328
rect 13964 14288 13970 14300
rect 6917 14263 6975 14269
rect 6917 14260 6929 14263
rect 6788 14232 6929 14260
rect 6788 14220 6794 14232
rect 6917 14229 6929 14232
rect 6963 14229 6975 14263
rect 6917 14223 6975 14229
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8846 14260 8852 14272
rect 8619 14232 8852 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 9858 14260 9864 14272
rect 9640 14232 9864 14260
rect 9640 14220 9646 14232
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 11793 14263 11851 14269
rect 11793 14229 11805 14263
rect 11839 14260 11851 14263
rect 12066 14260 12072 14272
rect 11839 14232 12072 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 13412 14232 13829 14260
rect 13412 14220 13418 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 14093 14263 14151 14269
rect 14093 14229 14105 14263
rect 14139 14260 14151 14263
rect 14458 14260 14464 14272
rect 14139 14232 14464 14260
rect 14139 14229 14151 14232
rect 14093 14223 14151 14229
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 14642 14220 14648 14272
rect 14700 14260 14706 14272
rect 14752 14260 14780 14300
rect 15381 14297 15393 14300
rect 15427 14297 15439 14331
rect 15381 14291 15439 14297
rect 14700 14232 14780 14260
rect 14700 14220 14706 14232
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 14884 14232 15301 14260
rect 14884 14220 14890 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 15289 14223 15347 14229
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3568 14028 3617 14056
rect 3568 14016 3574 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5166 14056 5172 14068
rect 4755 14028 5172 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 7742 14056 7748 14068
rect 5224 14028 6040 14056
rect 7703 14028 7748 14056
rect 5224 14016 5230 14028
rect 5902 13997 5908 14000
rect 3421 13991 3479 13997
rect 3421 13988 3433 13991
rect 2608 13960 3433 13988
rect 2406 13812 2412 13864
rect 2464 13852 2470 13864
rect 2608 13852 2636 13960
rect 3421 13957 3433 13960
rect 3467 13988 3479 13991
rect 5844 13991 5908 13997
rect 3467 13960 5764 13988
rect 3467 13957 3479 13960
rect 3421 13951 3479 13957
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 2731 13892 3249 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3237 13889 3249 13892
rect 3283 13920 3295 13923
rect 3326 13920 3332 13932
rect 3283 13892 3332 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3326 13880 3332 13892
rect 3384 13920 3390 13932
rect 3602 13920 3608 13932
rect 3384 13892 3608 13920
rect 3384 13880 3390 13892
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 5534 13920 5540 13932
rect 4663 13892 5540 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5736 13920 5764 13960
rect 5844 13957 5856 13991
rect 5890 13957 5908 13991
rect 5844 13951 5908 13957
rect 5902 13948 5908 13951
rect 5960 13948 5966 14000
rect 6012 13988 6040 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8478 14056 8484 14068
rect 8352 14028 8484 14056
rect 8352 14016 8358 14028
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 8849 14059 8907 14065
rect 8849 14025 8861 14059
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 6610 13991 6668 13997
rect 6610 13988 6622 13991
rect 6012 13960 6622 13988
rect 6610 13957 6622 13960
rect 6656 13957 6668 13991
rect 6610 13951 6668 13957
rect 6730 13948 6736 14000
rect 6788 13988 6794 14000
rect 8312 13988 8340 14016
rect 6788 13960 8340 13988
rect 8864 13988 8892 14019
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9180 14028 9229 14056
rect 9180 14016 9186 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 9490 14056 9496 14068
rect 9355 14028 9496 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9723 14028 10149 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 10137 14019 10195 14025
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 11238 14056 11244 14068
rect 10551 14028 11244 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11974 14056 11980 14068
rect 11379 14028 11980 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12897 14059 12955 14065
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 12986 14056 12992 14068
rect 12943 14028 12992 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 8864 13960 10057 13988
rect 6788 13948 6794 13960
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10870 13988 10876 14000
rect 10831 13960 10876 13988
rect 10045 13951 10103 13957
rect 10870 13948 10876 13960
rect 10928 13988 10934 14000
rect 11054 13988 11060 14000
rect 10928 13960 11060 13988
rect 10928 13948 10934 13960
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 11784 13991 11842 13997
rect 11784 13957 11796 13991
rect 11830 13988 11842 13991
rect 12802 13988 12808 14000
rect 11830 13960 12808 13988
rect 11830 13957 11842 13960
rect 11784 13951 11842 13957
rect 12802 13948 12808 13960
rect 12860 13988 12866 14000
rect 13262 13988 13268 14000
rect 12860 13960 13268 13988
rect 12860 13948 12866 13960
rect 13262 13948 13268 13960
rect 13320 13948 13326 14000
rect 14550 13988 14556 14000
rect 14511 13960 14556 13988
rect 14550 13948 14556 13960
rect 14608 13948 14614 14000
rect 15470 13988 15476 14000
rect 15431 13960 15476 13988
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 15620 13960 15665 13988
rect 15620 13948 15626 13960
rect 9582 13920 9588 13932
rect 5736 13892 9588 13920
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 10008 13892 10977 13920
rect 10008 13880 10014 13892
rect 10965 13889 10977 13892
rect 11011 13920 11023 13923
rect 11146 13920 11152 13932
rect 11011 13892 11152 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11146 13880 11152 13892
rect 11204 13920 11210 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 11204 13892 13001 13920
rect 11204 13880 11210 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2464 13824 2789 13852
rect 2464 13812 2470 13824
rect 2777 13821 2789 13824
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3786 13852 3792 13864
rect 3007 13824 3792 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4154 13852 4160 13864
rect 3896 13824 4160 13852
rect 3602 13744 3608 13796
rect 3660 13784 3666 13796
rect 3896 13784 3924 13824
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6144 13824 6377 13852
rect 6144 13812 6150 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6365 13815 6423 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8389 13855 8447 13861
rect 8389 13821 8401 13855
rect 8435 13852 8447 13855
rect 8846 13852 8852 13864
rect 8435 13824 8852 13852
rect 8435 13821 8447 13824
rect 8389 13815 8447 13821
rect 3660 13756 3924 13784
rect 3660 13744 3666 13756
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 5074 13716 5080 13728
rect 2556 13688 5080 13716
rect 2556 13676 2562 13688
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 6380 13716 6408 13815
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7432 13756 7849 13784
rect 7432 13744 7438 13756
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 8312 13784 8340 13815
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 9140 13784 9168 13815
rect 9876 13784 9904 13815
rect 9950 13784 9956 13796
rect 8312 13756 9260 13784
rect 9876 13756 9956 13784
rect 7837 13747 7895 13753
rect 7392 13716 7420 13744
rect 6380 13688 7420 13716
rect 9232 13716 9260 13756
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10704 13784 10732 13815
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 11388 13824 11529 13852
rect 11388 13812 11394 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14642 13852 14648 13864
rect 14507 13824 14648 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 10100 13756 10732 13784
rect 10100 13744 10106 13756
rect 10060 13716 10088 13744
rect 9232 13688 10088 13716
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 13814 13716 13820 13728
rect 10284 13688 13820 13716
rect 10284 13676 10290 13688
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 2682 13472 2688 13524
rect 2740 13512 2746 13524
rect 5074 13512 5080 13524
rect 2740 13484 5080 13512
rect 2740 13472 2746 13484
rect 5074 13472 5080 13484
rect 5132 13512 5138 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 5132 13484 5273 13512
rect 5132 13472 5138 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5534 13512 5540 13524
rect 5447 13484 5540 13512
rect 5261 13475 5319 13481
rect 5534 13472 5540 13484
rect 5592 13512 5598 13524
rect 6086 13512 6092 13524
rect 5592 13484 6092 13512
rect 5592 13472 5598 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 7374 13512 7380 13524
rect 7331 13484 7380 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 10226 13512 10232 13524
rect 8404 13484 10232 13512
rect 2869 13447 2927 13453
rect 2869 13444 2881 13447
rect 1964 13416 2881 13444
rect 1964 13317 1992 13416
rect 2869 13413 2881 13416
rect 2915 13413 2927 13447
rect 2869 13407 2927 13413
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 5902 13444 5908 13456
rect 5675 13416 5908 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 2682 13376 2688 13388
rect 2271 13348 2688 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 3510 13376 3516 13388
rect 3471 13348 3516 13376
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 7392 13385 7420 13472
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 7055 13348 7389 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7377 13345 7389 13348
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2372 13280 2421 13308
rect 2372 13268 2378 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 3234 13308 3240 13320
rect 3195 13280 3240 13308
rect 2409 13271 2467 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 5534 13308 5540 13320
rect 3927 13280 5540 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 1670 13240 1676 13252
rect 1631 13212 1676 13240
rect 1670 13200 1676 13212
rect 1728 13200 1734 13252
rect 3329 13243 3387 13249
rect 3329 13240 3341 13243
rect 2792 13212 3341 13240
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2792 13181 2820 13212
rect 3329 13209 3341 13212
rect 3375 13209 3387 13243
rect 3329 13203 3387 13209
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 4126 13243 4184 13249
rect 4126 13240 4138 13243
rect 3844 13212 4138 13240
rect 3844 13200 3850 13212
rect 4126 13209 4138 13212
rect 4172 13209 4184 13243
rect 4126 13203 4184 13209
rect 6454 13200 6460 13252
rect 6512 13240 6518 13252
rect 6742 13243 6800 13249
rect 6742 13240 6754 13243
rect 6512 13212 6754 13240
rect 6512 13200 6518 13212
rect 6742 13209 6754 13212
rect 6788 13209 6800 13243
rect 6742 13203 6800 13209
rect 7644 13243 7702 13249
rect 7644 13209 7656 13243
rect 7690 13240 7702 13243
rect 7742 13240 7748 13252
rect 7690 13212 7748 13240
rect 7690 13209 7702 13212
rect 7644 13203 7702 13209
rect 7742 13200 7748 13212
rect 7800 13200 7806 13252
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13141 2835 13175
rect 2777 13135 2835 13141
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 8404 13172 8432 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11606 13512 11612 13524
rect 11287 13484 11612 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12897 13515 12955 13521
rect 12124 13484 12434 13512
rect 12124 13472 12130 13484
rect 8757 13447 8815 13453
rect 8757 13413 8769 13447
rect 8803 13413 8815 13447
rect 8757 13407 8815 13413
rect 8772 13240 8800 13407
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8904 13348 9045 13376
rect 8904 13336 8910 13348
rect 9033 13345 9045 13348
rect 9079 13376 9091 13379
rect 9122 13376 9128 13388
rect 9079 13348 9128 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 11330 13376 11336 13388
rect 11291 13348 11336 13376
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 12406 13376 12434 13484
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13170 13512 13176 13524
rect 12943 13484 13176 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13998 13512 14004 13524
rect 13412 13484 14004 13512
rect 13412 13472 13418 13484
rect 13998 13472 14004 13484
rect 14056 13512 14062 13524
rect 14826 13512 14832 13524
rect 14056 13484 14832 13512
rect 14056 13472 14062 13484
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15151 13515 15209 13521
rect 15151 13481 15163 13515
rect 15197 13512 15209 13515
rect 15470 13512 15476 13524
rect 15197 13484 15476 13512
rect 15197 13481 15209 13484
rect 15151 13475 15209 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 15620 13484 15665 13512
rect 15620 13472 15626 13484
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 12406 13348 14657 13376
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9861 13311 9919 13317
rect 9861 13308 9873 13311
rect 9815 13280 9873 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9861 13277 9873 13280
rect 9907 13308 9919 13311
rect 11348 13308 11376 13336
rect 9907 13280 11376 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 14516 13280 14565 13308
rect 14516 13268 14522 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15048 13311 15106 13317
rect 15048 13308 15060 13311
rect 14976 13280 15060 13308
rect 14976 13268 14982 13280
rect 15048 13277 15060 13280
rect 15094 13277 15106 13311
rect 15048 13271 15106 13277
rect 10134 13249 10140 13252
rect 10128 13240 10140 13249
rect 8772 13212 9536 13240
rect 10095 13212 10140 13240
rect 3292 13144 8432 13172
rect 3292 13132 3298 13144
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8536 13144 9137 13172
rect 8536 13132 8542 13144
rect 9125 13141 9137 13144
rect 9171 13141 9183 13175
rect 9508 13172 9536 13212
rect 10128 13203 10140 13212
rect 10134 13200 10140 13203
rect 10192 13200 10198 13252
rect 11578 13243 11636 13249
rect 11578 13240 11590 13243
rect 10888 13212 11590 13240
rect 10888 13172 10916 13212
rect 11578 13209 11590 13212
rect 11624 13240 11636 13243
rect 12894 13240 12900 13252
rect 11624 13212 12900 13240
rect 11624 13209 11636 13212
rect 11578 13203 11636 13209
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13722 13240 13728 13252
rect 13412 13212 13728 13240
rect 13412 13200 13418 13212
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 9508 13144 10916 13172
rect 9125 13135 9183 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 12584 13144 12725 13172
rect 12584 13132 12590 13144
rect 12713 13141 12725 13144
rect 12759 13141 12771 13175
rect 12713 13135 12771 13141
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 13320 13144 14105 13172
rect 13320 13132 13326 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14240 13144 14473 13172
rect 14240 13132 14246 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 2372 12940 2421 12968
rect 2372 12928 2378 12940
rect 2409 12937 2421 12940
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 3568 12940 6193 12968
rect 3568 12928 3574 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 7374 12968 7380 12980
rect 7331 12940 7380 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 2777 12903 2835 12909
rect 2777 12869 2789 12903
rect 2823 12900 2835 12903
rect 2823 12872 3280 12900
rect 2823 12869 2835 12872
rect 2777 12863 2835 12869
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2792 12832 2820 12863
rect 2363 12804 2820 12832
rect 2869 12835 2927 12841
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3142 12832 3148 12844
rect 2915 12804 3148 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3252 12832 3280 12872
rect 3326 12860 3332 12912
rect 3384 12900 3390 12912
rect 3786 12900 3792 12912
rect 3384 12872 3792 12900
rect 3384 12860 3390 12872
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 5534 12900 5540 12912
rect 4816 12872 5540 12900
rect 3418 12832 3424 12844
rect 3252 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12832 3482 12844
rect 3970 12832 3976 12844
rect 3476 12804 3976 12832
rect 3476 12792 3482 12804
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4442 12835 4500 12841
rect 4442 12832 4454 12835
rect 4212 12804 4454 12832
rect 4212 12792 4218 12804
rect 4442 12801 4454 12804
rect 4488 12801 4500 12835
rect 4442 12795 4500 12801
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 4816 12841 4844 12872
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 5074 12841 5080 12844
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4672 12804 4721 12832
rect 4672 12792 4678 12804
rect 4709 12801 4721 12804
rect 4755 12832 4767 12835
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 4755 12804 4813 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 4801 12801 4813 12804
rect 4847 12801 4859 12835
rect 5068 12832 5080 12841
rect 5035 12804 5080 12832
rect 4801 12795 4859 12801
rect 5068 12795 5080 12804
rect 5074 12792 5080 12795
rect 5132 12792 5138 12844
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3326 12764 3332 12776
rect 3099 12736 3332 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3326 12724 3332 12736
rect 3384 12724 3390 12776
rect 6196 12764 6224 12931
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 13262 12968 13268 12980
rect 8404 12940 13268 12968
rect 7392 12841 7420 12928
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7633 12835 7691 12841
rect 7633 12832 7645 12835
rect 7377 12795 7435 12801
rect 7484 12804 7645 12832
rect 7484 12764 7512 12804
rect 7633 12801 7645 12804
rect 7679 12801 7691 12835
rect 7633 12795 7691 12801
rect 6196 12736 7512 12764
rect 2746 12668 3464 12696
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2746 12628 2774 12668
rect 3326 12628 3332 12640
rect 2648 12600 2774 12628
rect 3287 12600 3332 12628
rect 2648 12588 2654 12600
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 3436 12628 3464 12668
rect 8404 12628 8432 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13725 12971 13783 12977
rect 13412 12940 13457 12968
rect 13412 12928 13418 12940
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 13771 12940 14289 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 14277 12931 14335 12937
rect 14645 12971 14703 12977
rect 14645 12937 14657 12971
rect 14691 12968 14703 12971
rect 15010 12968 15016 12980
rect 14691 12940 15016 12968
rect 14691 12937 14703 12940
rect 14645 12931 14703 12937
rect 15010 12928 15016 12940
rect 15068 12968 15074 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 15068 12940 15117 12968
rect 15068 12928 15074 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 8754 12860 8760 12912
rect 8812 12900 8818 12912
rect 8941 12903 8999 12909
rect 8941 12900 8953 12903
rect 8812 12872 8953 12900
rect 8812 12860 8818 12872
rect 8941 12869 8953 12872
rect 8987 12900 8999 12903
rect 11330 12900 11336 12912
rect 8987 12872 10456 12900
rect 11291 12872 11336 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 9306 12832 9312 12844
rect 8772 12804 9312 12832
rect 8772 12705 8800 12804
rect 9306 12792 9312 12804
rect 9364 12832 9370 12844
rect 10428 12841 10456 12872
rect 11330 12860 11336 12872
rect 11388 12860 11394 12912
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 11762 12903 11820 12909
rect 11762 12900 11774 12903
rect 11664 12872 11774 12900
rect 11664 12860 11670 12872
rect 11762 12869 11774 12872
rect 11808 12869 11820 12903
rect 13372 12900 13400 12928
rect 14737 12903 14795 12909
rect 14737 12900 14749 12903
rect 13372 12872 14749 12900
rect 11762 12863 11820 12869
rect 14737 12869 14749 12872
rect 14783 12869 14795 12903
rect 14737 12863 14795 12869
rect 10146 12835 10204 12841
rect 10146 12832 10158 12835
rect 9364 12804 10158 12832
rect 9364 12792 9370 12804
rect 10146 12801 10158 12804
rect 10192 12801 10204 12835
rect 10146 12795 10204 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 11348 12832 11376 12860
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10459 12804 11529 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 11517 12795 11575 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13906 12764 13912 12776
rect 13679 12736 13912 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 14734 12764 14740 12776
rect 14516 12736 14740 12764
rect 14516 12724 14522 12736
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 14884 12736 14929 12764
rect 14884 12724 14890 12736
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12665 8815 12699
rect 8757 12659 8815 12665
rect 8938 12656 8944 12708
rect 8996 12696 9002 12708
rect 9033 12699 9091 12705
rect 9033 12696 9045 12699
rect 8996 12668 9045 12696
rect 8996 12656 9002 12668
rect 9033 12665 9045 12668
rect 9079 12665 9091 12699
rect 9033 12659 9091 12665
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12860 12668 12909 12696
rect 12860 12656 12866 12668
rect 12897 12665 12909 12668
rect 12943 12696 12955 12699
rect 14182 12696 14188 12708
rect 12943 12668 13768 12696
rect 14143 12668 14188 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 3436 12600 8432 12628
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10226 12628 10232 12640
rect 9824 12600 10232 12628
rect 9824 12588 9830 12600
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12158 12628 12164 12640
rect 11848 12600 12164 12628
rect 11848 12588 11854 12600
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 13740 12628 13768 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14826 12628 14832 12640
rect 13740 12600 14832 12628
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3142 12424 3148 12436
rect 2915 12396 3148 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3970 12424 3976 12436
rect 3476 12396 3976 12424
rect 3476 12384 3482 12396
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6512 12396 6745 12424
rect 6512 12384 6518 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 9122 12424 9128 12436
rect 6733 12387 6791 12393
rect 7024 12396 9128 12424
rect 5166 12356 5172 12368
rect 2240 12328 5172 12356
rect 2240 12297 2268 12328
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 7024 12356 7052 12396
rect 9122 12384 9128 12396
rect 9180 12424 9186 12436
rect 9306 12424 9312 12436
rect 9180 12396 9312 12424
rect 9180 12384 9186 12396
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 10686 12424 10692 12436
rect 9416 12396 10692 12424
rect 5500 12328 7052 12356
rect 5500 12316 5506 12328
rect 8110 12316 8116 12368
rect 8168 12356 8174 12368
rect 9416 12356 9444 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11606 12424 11612 12436
rect 11287 12396 11612 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12032 12396 13308 12424
rect 12032 12384 12038 12396
rect 8168 12328 9444 12356
rect 11149 12359 11207 12365
rect 8168 12316 8174 12328
rect 11149 12325 11161 12359
rect 11195 12356 11207 12359
rect 11330 12356 11336 12368
rect 11195 12328 11336 12356
rect 11195 12325 11207 12328
rect 11149 12319 11207 12325
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12257 2283 12291
rect 2225 12251 2283 12257
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12288 3571 12291
rect 4154 12288 4160 12300
rect 3559 12260 4160 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 8036 12260 9352 12288
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12220 2651 12223
rect 3878 12220 3884 12232
rect 2639 12192 3884 12220
rect 2639 12189 2651 12192
rect 2593 12183 2651 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4614 12220 4620 12232
rect 4527 12192 4620 12220
rect 4614 12180 4620 12192
rect 4672 12220 4678 12232
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4672 12192 4997 12220
rect 4672 12180 4678 12192
rect 4985 12189 4997 12192
rect 5031 12220 5043 12223
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 5031 12192 5181 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5169 12189 5181 12192
rect 5215 12220 5227 12223
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5215 12192 5457 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5445 12189 5457 12192
rect 5491 12220 5503 12223
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 5491 12192 6653 12220
rect 5491 12189 5503 12192
rect 5445 12183 5503 12189
rect 6641 12189 6653 12192
rect 6687 12220 6699 12223
rect 7282 12220 7288 12232
rect 6687 12192 7288 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 3237 12155 3295 12161
rect 3237 12121 3249 12155
rect 3283 12152 3295 12155
rect 4246 12152 4252 12164
rect 3283 12124 4252 12152
rect 3283 12121 3295 12124
rect 3237 12115 3295 12121
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 7868 12155 7926 12161
rect 7868 12121 7880 12155
rect 7914 12152 7926 12155
rect 8036 12152 8064 12260
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8754 12220 8760 12232
rect 8113 12183 8171 12189
rect 8266 12192 8760 12220
rect 7914 12124 8064 12152
rect 8128 12152 8156 12183
rect 8266 12152 8294 12192
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 8128 12124 8294 12152
rect 7914 12121 7926 12124
rect 7868 12115 7926 12121
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 1544 12056 1593 12084
rect 1544 12044 1550 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1581 12047 1639 12053
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2777 12087 2835 12093
rect 2096 12056 2141 12084
rect 2096 12044 2102 12056
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 3329 12087 3387 12093
rect 3329 12084 3341 12087
rect 2823 12056 3341 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3329 12053 3341 12056
rect 3375 12084 3387 12087
rect 3694 12084 3700 12096
rect 3375 12056 3700 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 8110 12084 8116 12096
rect 4028 12056 8116 12084
rect 4028 12044 4034 12056
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8352 12056 8953 12084
rect 8352 12044 8358 12056
rect 8941 12053 8953 12056
rect 8987 12084 8999 12087
rect 9030 12084 9036 12096
rect 8987 12056 9036 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9324 12084 9352 12260
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10870 12220 10876 12232
rect 10367 12192 10876 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10870 12180 10876 12192
rect 10928 12220 10934 12232
rect 11348 12220 11376 12316
rect 13280 12297 13308 12396
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13872 12396 14105 12424
rect 13872 12384 13878 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 15197 12427 15255 12433
rect 15197 12424 15209 12427
rect 15160 12396 15209 12424
rect 15160 12384 15166 12396
rect 15197 12393 15209 12396
rect 15243 12393 15255 12427
rect 15197 12387 15255 12393
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 14642 12288 14648 12300
rect 13495 12260 14648 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 14642 12248 14648 12260
rect 14700 12248 14706 12300
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 14826 12288 14832 12300
rect 14783 12260 14832 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 12618 12220 12624 12232
rect 10928 12192 12624 12220
rect 10928 12180 10934 12192
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 14550 12220 14556 12232
rect 14463 12192 14556 12220
rect 14550 12180 14556 12192
rect 14608 12220 14614 12232
rect 15102 12220 15108 12232
rect 14608 12192 15108 12220
rect 14608 12180 14614 12192
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 10076 12155 10134 12161
rect 10076 12152 10088 12155
rect 9548 12124 10088 12152
rect 9548 12112 9554 12124
rect 10076 12121 10088 12124
rect 10122 12152 10134 12155
rect 11422 12152 11428 12164
rect 10122 12124 11428 12152
rect 10122 12121 10134 12124
rect 10076 12115 10134 12121
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 12376 12155 12434 12161
rect 12376 12121 12388 12155
rect 12422 12152 12434 12155
rect 12526 12152 12532 12164
rect 12422 12124 12532 12152
rect 12422 12121 12434 12124
rect 12376 12115 12434 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 14461 12155 14519 12161
rect 12636 12124 13032 12152
rect 11790 12084 11796 12096
rect 9324 12056 11796 12084
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 11882 12044 11888 12096
rect 11940 12084 11946 12096
rect 12636 12084 12664 12124
rect 13004 12096 13032 12124
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14921 12155 14979 12161
rect 14921 12152 14933 12155
rect 14507 12124 14933 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 14921 12121 14933 12124
rect 14967 12121 14979 12155
rect 14921 12115 14979 12121
rect 12802 12084 12808 12096
rect 11940 12056 12664 12084
rect 12763 12056 12808 12084
rect 11940 12044 11946 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 13044 12056 13185 12084
rect 13044 12044 13050 12056
rect 13173 12053 13185 12056
rect 13219 12084 13231 12087
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 13219 12056 13645 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2774 11880 2780 11892
rect 2547 11852 2780 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3878 11880 3884 11892
rect 3467 11852 3884 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4154 11880 4160 11892
rect 4111 11852 4160 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 9214 11880 9220 11892
rect 5092 11852 9220 11880
rect 1762 11812 1768 11824
rect 1723 11784 1768 11812
rect 1762 11772 1768 11784
rect 1820 11772 1826 11824
rect 3973 11815 4031 11821
rect 3973 11781 3985 11815
rect 4019 11812 4031 11815
rect 4246 11812 4252 11824
rect 4019 11784 4252 11812
rect 4019 11781 4031 11784
rect 3973 11775 4031 11781
rect 4246 11772 4252 11784
rect 4304 11812 4310 11824
rect 5092 11812 5120 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 4304 11784 5120 11812
rect 4304 11772 4310 11784
rect 5166 11772 5172 11824
rect 5224 11821 5230 11824
rect 5224 11812 5236 11821
rect 5224 11784 5269 11812
rect 5224 11775 5236 11784
rect 5224 11772 5230 11775
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 5592 11784 8064 11812
rect 5592 11772 5598 11784
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 2498 11704 2504 11756
rect 2556 11744 2562 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2556 11716 2605 11744
rect 2556 11704 2562 11716
rect 2593 11713 2605 11716
rect 2639 11744 2651 11747
rect 3142 11744 3148 11756
rect 2639 11716 3148 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 4338 11744 4344 11756
rect 3375 11716 4344 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 8036 11744 8064 11784
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 9401 11815 9459 11821
rect 9401 11812 9413 11815
rect 9088 11784 9413 11812
rect 9088 11772 9094 11784
rect 9401 11781 9413 11784
rect 9447 11812 9459 11815
rect 12253 11815 12311 11821
rect 9447 11784 10916 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 10888 11756 10916 11784
rect 12253 11781 12265 11815
rect 12299 11812 12311 11815
rect 12710 11812 12716 11824
rect 12299 11784 12716 11812
rect 12299 11781 12311 11784
rect 12253 11775 12311 11781
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 9858 11744 9864 11756
rect 4457 11716 7972 11744
rect 8036 11716 9864 11744
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 2823 11648 3525 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2130 11540 2136 11552
rect 2091 11512 2136 11540
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2648 11512 2973 11540
rect 2648 11500 2654 11512
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 3436 11540 3464 11648
rect 3513 11645 3525 11648
rect 3559 11645 3571 11679
rect 3513 11639 3571 11645
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 4457 11676 4485 11716
rect 3936 11648 4485 11676
rect 5445 11679 5503 11685
rect 3936 11636 3942 11648
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5491 11648 5672 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 3510 11540 3516 11552
rect 3436 11512 3516 11540
rect 2961 11503 3019 11509
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 3694 11500 3700 11552
rect 3752 11540 3758 11552
rect 5074 11540 5080 11552
rect 3752 11512 5080 11540
rect 3752 11500 3758 11512
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5534 11540 5540 11552
rect 5316 11512 5540 11540
rect 5316 11500 5322 11512
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5644 11549 5672 11648
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5675 11512 5825 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5813 11509 5825 11512
rect 5859 11540 5871 11543
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5859 11512 6009 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5997 11509 6009 11512
rect 6043 11540 6055 11543
rect 7282 11540 7288 11552
rect 6043 11512 7288 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 7282 11500 7288 11512
rect 7340 11540 7346 11552
rect 7834 11540 7840 11552
rect 7340 11512 7840 11540
rect 7340 11500 7346 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 7944 11540 7972 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10617 11747 10675 11753
rect 10617 11713 10629 11747
rect 10663 11744 10675 11747
rect 10663 11716 10824 11744
rect 10663 11713 10675 11716
rect 10617 11707 10675 11713
rect 10796 11676 10824 11716
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 12345 11747 12403 11753
rect 10928 11716 10973 11744
rect 10928 11704 10934 11716
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12526 11744 12532 11756
rect 12391 11716 12532 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 13722 11744 13728 11756
rect 13683 11716 13728 11744
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 11606 11676 11612 11688
rect 10796 11648 11612 11676
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12124 11648 12449 11676
rect 12124 11636 12130 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13228 11648 13829 11676
rect 13228 11636 13234 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14642 11676 14648 11688
rect 14047 11648 14648 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 14016 11608 14044 11639
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 11020 11580 14044 11608
rect 11020 11568 11026 11580
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 7944 11512 11897 11540
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 13170 11540 13176 11552
rect 13131 11512 13176 11540
rect 11885 11503 11943 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 14277 11543 14335 11549
rect 14277 11540 14289 11543
rect 13780 11512 14289 11540
rect 13780 11500 13786 11512
rect 14277 11509 14289 11512
rect 14323 11540 14335 11543
rect 15562 11540 15568 11552
rect 14323 11512 15568 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2041 11339 2099 11345
rect 2041 11336 2053 11339
rect 2004 11308 2053 11336
rect 2004 11296 2010 11308
rect 2041 11305 2053 11308
rect 2087 11305 2099 11339
rect 5810 11336 5816 11348
rect 2041 11299 2099 11305
rect 3344 11308 5816 11336
rect 2869 11271 2927 11277
rect 2869 11268 2881 11271
rect 2424 11240 2881 11268
rect 2424 11141 2452 11240
rect 2869 11237 2881 11240
rect 2915 11237 2927 11271
rect 2869 11231 2927 11237
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2556 11172 2605 11200
rect 2556 11160 2562 11172
rect 2593 11169 2605 11172
rect 2639 11200 2651 11203
rect 3344 11200 3372 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 7156 11308 7297 11336
rect 7156 11296 7162 11308
rect 7285 11305 7297 11308
rect 7331 11336 7343 11339
rect 7650 11336 7656 11348
rect 7331 11308 7656 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 9398 11336 9404 11348
rect 8803 11308 9404 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10192 11308 10517 11336
rect 10192 11296 10198 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 10870 11336 10876 11348
rect 10505 11299 10563 11305
rect 10612 11308 10876 11336
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 4028 11240 4077 11268
rect 4028 11228 4034 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4338 11268 4344 11280
rect 4299 11240 4344 11268
rect 4065 11231 4123 11237
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 9030 11268 9036 11280
rect 8991 11240 9036 11268
rect 9030 11228 9036 11240
rect 9088 11268 9094 11280
rect 9088 11240 9168 11268
rect 9088 11228 9094 11240
rect 3510 11200 3516 11212
rect 2639 11172 3372 11200
rect 3471 11172 3516 11200
rect 2639 11169 2651 11172
rect 2593 11163 2651 11169
rect 3510 11160 3516 11172
rect 3568 11160 3574 11212
rect 9140 11209 9168 11240
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 10612 11209 10640 11308
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14568 11308 15025 11336
rect 14568 11209 14596 11308
rect 15013 11305 15025 11308
rect 15059 11336 15071 11339
rect 15286 11336 15292 11348
rect 15059 11308 15292 11336
rect 15059 11305 15071 11308
rect 15013 11299 15071 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10560 11172 10609 11200
rect 10560 11160 10566 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 14700 11172 14745 11200
rect 14700 11160 14706 11172
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 3326 11132 3332 11144
rect 2409 11095 2467 11101
rect 2746 11104 3332 11132
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2746 11064 2774 11104
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3528 11132 3556 11160
rect 9398 11141 9404 11144
rect 4433 11135 4491 11141
rect 3528 11104 3924 11132
rect 1995 11036 2774 11064
rect 3237 11067 3295 11073
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 3283 11036 3801 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3896 11064 3924 11104
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 4479 11104 5917 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 5905 11101 5917 11104
rect 5951 11132 5963 11135
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 5951 11104 7389 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 7377 11101 7389 11104
rect 7423 11132 7435 11135
rect 9392 11132 9404 11141
rect 7423 11104 7880 11132
rect 9359 11104 9404 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 7852 11076 7880 11104
rect 9392 11095 9404 11104
rect 9398 11092 9404 11095
rect 9456 11092 9462 11144
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 12676 11104 13461 11132
rect 12676 11092 12682 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 4678 11067 4736 11073
rect 4678 11064 4690 11067
rect 3896 11036 4690 11064
rect 3789 11027 3847 11033
rect 4678 11033 4690 11036
rect 4724 11033 4736 11067
rect 4678 11027 4736 11033
rect 6172 11067 6230 11073
rect 6172 11033 6184 11067
rect 6218 11064 6230 11067
rect 6270 11064 6276 11076
rect 6218 11036 6276 11064
rect 6218 11033 6230 11036
rect 6172 11027 6230 11033
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 7644 11067 7702 11073
rect 7644 11033 7656 11067
rect 7690 11064 7702 11067
rect 7690 11036 7788 11064
rect 7690 11033 7702 11036
rect 7644 11027 7702 11033
rect 2501 10999 2559 11005
rect 2501 10965 2513 10999
rect 2547 10996 2559 10999
rect 2590 10996 2596 11008
rect 2547 10968 2596 10996
rect 2547 10965 2559 10968
rect 2501 10959 2559 10965
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 7760 10996 7788 11036
rect 7834 11024 7840 11076
rect 7892 11024 7898 11076
rect 8938 11064 8944 11076
rect 7944 11036 8944 11064
rect 7944 10996 7972 11036
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10842 11067 10900 11073
rect 10842 11064 10854 11067
rect 10008 11036 10854 11064
rect 10008 11024 10014 11036
rect 10842 11033 10854 11036
rect 10888 11064 10900 11067
rect 10962 11064 10968 11076
rect 10888 11036 10968 11064
rect 10888 11033 10900 11036
rect 10842 11027 10900 11033
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 13182 11067 13240 11073
rect 13182 11064 13194 11067
rect 11992 11036 13194 11064
rect 7760 10968 7972 10996
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 11992 11005 12020 11036
rect 13182 11033 13194 11036
rect 13228 11033 13240 11067
rect 13182 11027 13240 11033
rect 13909 11067 13967 11073
rect 13909 11033 13921 11067
rect 13955 11064 13967 11067
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 13955 11036 14473 11064
rect 13955 11033 13967 11036
rect 13909 11027 13967 11033
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11940 10968 11989 10996
rect 11940 10956 11946 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 14090 10996 14096 11008
rect 12124 10968 12169 10996
rect 14051 10968 14096 10996
rect 12124 10956 12130 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 1857 10795 1915 10801
rect 1857 10761 1869 10795
rect 1903 10792 1915 10795
rect 2038 10792 2044 10804
rect 1903 10764 2044 10792
rect 1903 10761 1915 10764
rect 1857 10755 1915 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 2188 10764 2237 10792
rect 2188 10752 2194 10764
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2363 10764 2697 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3191 10764 3525 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 5166 10792 5172 10804
rect 4755 10764 5172 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 6328 10764 6469 10792
rect 6328 10752 6334 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8067 10764 8861 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 8849 10761 8861 10764
rect 8895 10792 8907 10795
rect 9030 10792 9036 10804
rect 8895 10764 9036 10792
rect 8895 10761 8907 10764
rect 8849 10755 8907 10761
rect 3973 10727 4031 10733
rect 3973 10693 3985 10727
rect 4019 10724 4031 10727
rect 4338 10724 4344 10736
rect 4019 10696 4344 10724
rect 4019 10693 4031 10696
rect 3973 10687 4031 10693
rect 4338 10684 4344 10696
rect 4396 10724 4402 10736
rect 5442 10724 5448 10736
rect 4396 10696 5448 10724
rect 4396 10684 4402 10696
rect 5442 10684 5448 10696
rect 5500 10684 5506 10736
rect 5626 10684 5632 10736
rect 5684 10684 5690 10736
rect 5810 10684 5816 10736
rect 5868 10733 5874 10736
rect 5868 10724 5880 10733
rect 5868 10696 5913 10724
rect 5868 10687 5880 10696
rect 5868 10684 5874 10687
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3418 10656 3424 10668
rect 3099 10628 3424 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3418 10616 3424 10628
rect 3476 10656 3482 10668
rect 3786 10656 3792 10668
rect 3476 10628 3792 10656
rect 3476 10616 3482 10628
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4062 10656 4068 10668
rect 3927 10628 4068 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4062 10616 4068 10628
rect 4120 10656 4126 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4120 10628 4445 10656
rect 4120 10616 4126 10628
rect 4433 10625 4445 10628
rect 4479 10656 4491 10659
rect 5644 10656 5672 10684
rect 4479 10628 5672 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 7558 10616 7564 10668
rect 7616 10665 7622 10668
rect 7616 10656 7628 10665
rect 7616 10628 7661 10656
rect 7616 10619 7628 10628
rect 7616 10616 7622 10619
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8036 10656 8064 10755
rect 8956 10665 8984 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10008 10764 10333 10792
rect 10008 10752 10014 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10502 10792 10508 10804
rect 10463 10764 10508 10792
rect 10321 10755 10379 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 11296 10764 11989 10792
rect 11296 10752 11302 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 12618 10792 12624 10804
rect 12579 10764 12624 10792
rect 11977 10755 12035 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 13354 10792 13360 10804
rect 13311 10764 13360 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 9208 10727 9266 10733
rect 9208 10693 9220 10727
rect 9254 10724 9266 10727
rect 10042 10724 10048 10736
rect 9254 10696 10048 10724
rect 9254 10693 9266 10696
rect 9208 10687 9266 10693
rect 10042 10684 10048 10696
rect 10100 10684 10106 10736
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10520 10724 10548 10752
rect 10192 10696 10548 10724
rect 12069 10727 12127 10733
rect 10192 10684 10198 10696
rect 12069 10693 12081 10727
rect 12115 10724 12127 10727
rect 12802 10724 12808 10736
rect 12115 10696 12808 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 13173 10727 13231 10733
rect 13173 10693 13185 10727
rect 13219 10724 13231 10727
rect 14090 10724 14096 10736
rect 13219 10696 14096 10724
rect 13219 10693 13231 10696
rect 13173 10687 13231 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 7892 10628 8064 10656
rect 8941 10659 8999 10665
rect 7892 10616 7898 10628
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3510 10588 3516 10600
rect 3375 10560 3516 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 4154 10588 4160 10600
rect 4115 10560 4160 10588
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 6089 10551 6147 10557
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5718 10452 5724 10464
rect 4571 10424 5724 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5718 10412 5724 10424
rect 5776 10452 5782 10464
rect 6104 10452 6132 10551
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 11900 10520 11928 10548
rect 13372 10520 13400 10551
rect 11900 10492 13400 10520
rect 5776 10424 6132 10452
rect 12437 10455 12495 10461
rect 5776 10412 5782 10424
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12768 10424 12817 10452
rect 12768 10412 12774 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 14550 10452 14556 10464
rect 13412 10424 14556 10452
rect 13412 10412 13418 10424
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 3568 10220 3893 10248
rect 3568 10208 3574 10220
rect 3881 10217 3893 10220
rect 3927 10217 3939 10251
rect 8754 10248 8760 10260
rect 3881 10211 3939 10217
rect 4356 10220 8412 10248
rect 8715 10220 8760 10248
rect 4356 10180 4384 10220
rect 1964 10152 4384 10180
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1964 10053 1992 10152
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 1949 10007 2007 10013
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 3878 10044 3884 10056
rect 2547 10016 3884 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4994 10047 5052 10053
rect 4994 10044 5006 10047
rect 4212 10016 5006 10044
rect 4212 10004 4218 10016
rect 4994 10013 5006 10016
rect 5040 10044 5052 10047
rect 5261 10047 5319 10053
rect 5040 10016 5111 10044
rect 5040 10013 5052 10016
rect 4994 10007 5052 10013
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2832 9880 2973 9908
rect 2832 9868 2838 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 2961 9871 3019 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 4338 9908 4344 9920
rect 3651 9880 4344 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 5083 9908 5111 10016
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5307 10016 5457 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5445 10013 5457 10016
rect 5491 10044 5503 10047
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5491 10016 5641 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5629 10013 5641 10016
rect 5675 10044 5687 10047
rect 5718 10044 5724 10056
rect 5675 10016 5724 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 5718 10004 5724 10016
rect 5776 10044 5782 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5776 10016 5825 10044
rect 5776 10004 5782 10016
rect 5813 10013 5825 10016
rect 5859 10044 5871 10047
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 5859 10016 7297 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 7285 10013 7297 10016
rect 7331 10044 7343 10047
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7331 10016 7389 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7377 10013 7389 10016
rect 7423 10044 7435 10047
rect 8110 10044 8116 10056
rect 7423 10016 8116 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8384 10044 8412 10220
rect 8754 10208 8760 10220
rect 8812 10248 8818 10260
rect 9030 10248 9036 10260
rect 8812 10220 9036 10248
rect 8812 10208 8818 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10134 10248 10140 10260
rect 10091 10220 10140 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 13814 10248 13820 10260
rect 11480 10220 13820 10248
rect 11480 10208 11486 10220
rect 13814 10208 13820 10220
rect 13872 10248 13878 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 13872 10220 14381 10248
rect 13872 10208 13878 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 10152 10121 10180 10208
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 11204 10084 13185 10112
rect 11204 10072 11210 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 14384 10044 14412 10211
rect 15102 10112 15108 10124
rect 15063 10084 15108 10112
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 8384 10016 12434 10044
rect 14384 10016 15025 10044
rect 7650 9985 7656 9988
rect 7040 9979 7098 9985
rect 7040 9945 7052 9979
rect 7086 9976 7098 9979
rect 7644 9976 7656 9985
rect 7086 9948 7512 9976
rect 7611 9948 7656 9976
rect 7086 9945 7098 9948
rect 7040 9939 7098 9945
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5083 9880 5917 9908
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 7484 9908 7512 9948
rect 7644 9939 7656 9948
rect 7650 9936 7656 9939
rect 7708 9936 7714 9988
rect 9582 9976 9588 9988
rect 7944 9948 9588 9976
rect 7944 9908 7972 9948
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 10404 9979 10462 9985
rect 10404 9945 10416 9979
rect 10450 9976 10462 9979
rect 12066 9976 12072 9988
rect 10450 9948 12072 9976
rect 10450 9945 10462 9948
rect 10404 9939 10462 9945
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 7484 9880 7972 9908
rect 11517 9911 11575 9917
rect 5905 9871 5963 9877
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11606 9908 11612 9920
rect 11563 9880 11612 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 12406 9908 12434 10016
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 14274 9976 14280 9988
rect 13035 9948 14280 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 14384 9948 14933 9976
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12406 9880 12633 9908
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 12621 9871 12679 9877
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13136 9880 13181 9908
rect 13136 9868 13142 9880
rect 13630 9868 13636 9920
rect 13688 9908 13694 9920
rect 14384 9908 14412 9948
rect 14921 9945 14933 9948
rect 14967 9976 14979 9979
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14967 9948 15393 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15381 9945 15393 9948
rect 15427 9976 15439 9979
rect 15470 9976 15476 9988
rect 15427 9948 15476 9976
rect 15427 9945 15439 9948
rect 15381 9939 15439 9945
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 14550 9908 14556 9920
rect 13688 9880 14412 9908
rect 14511 9880 14556 9908
rect 13688 9868 13694 9880
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 5718 9704 5724 9716
rect 5679 9676 5724 9704
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 9582 9704 9588 9716
rect 9495 9676 9588 9704
rect 9582 9664 9588 9676
rect 9640 9704 9646 9716
rect 11146 9704 11152 9716
rect 9640 9676 11152 9704
rect 9640 9664 9646 9676
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 13136 9676 13185 9704
rect 13136 9664 13142 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 14274 9704 14280 9716
rect 14235 9676 14280 9704
rect 13173 9667 13231 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14737 9707 14795 9713
rect 14737 9704 14749 9707
rect 14608 9676 14749 9704
rect 14608 9664 14614 9676
rect 14737 9673 14749 9676
rect 14783 9673 14795 9707
rect 14737 9667 14795 9673
rect 2406 9596 2412 9648
rect 2464 9636 2470 9648
rect 2464 9608 3004 9636
rect 2464 9596 2470 9608
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2038 9568 2044 9580
rect 1995 9540 2044 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2648 9540 2697 9568
rect 2648 9528 2654 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 2976 9509 3004 9608
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 5362 9571 5420 9577
rect 5362 9568 5374 9571
rect 3936 9540 5374 9568
rect 3936 9528 3942 9540
rect 5362 9537 5374 9540
rect 5408 9537 5420 9571
rect 5362 9531 5420 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5736 9568 5764 9664
rect 7592 9639 7650 9645
rect 7592 9605 7604 9639
rect 7638 9636 7650 9639
rect 8312 9636 8340 9664
rect 7638 9608 8340 9636
rect 7638 9605 7650 9608
rect 7592 9599 7650 9605
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 10192 9608 11253 9636
rect 10192 9596 10198 9608
rect 6089 9571 6147 9577
rect 6089 9568 6101 9571
rect 5675 9540 6101 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6089 9537 6101 9540
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7883 9540 8033 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 8021 9537 8033 9540
rect 8067 9568 8079 9571
rect 8110 9568 8116 9580
rect 8067 9540 8116 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 10980 9577 11008 9608
rect 11241 9605 11253 9608
rect 11287 9636 11299 9639
rect 11287 9608 12940 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 8369 9571 8427 9577
rect 8369 9568 8381 9571
rect 8260 9540 8381 9568
rect 8260 9528 8266 9540
rect 8369 9537 8381 9540
rect 8415 9537 8427 9571
rect 8369 9531 8427 9537
rect 10709 9571 10767 9577
rect 10709 9537 10721 9571
rect 10755 9568 10767 9571
rect 10965 9571 11023 9577
rect 10755 9540 10916 9568
rect 10755 9537 10767 9540
rect 10709 9531 10767 9537
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1452 9472 1685 9500
rect 1452 9460 1458 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 1673 9463 1731 9469
rect 2700 9472 2789 9500
rect 2700 9444 2728 9472
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 10888 9500 10916 9540
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 12641 9571 12699 9577
rect 11011 9540 11045 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 12641 9537 12653 9571
rect 12687 9568 12699 9571
rect 12802 9568 12808 9580
rect 12687 9540 12808 9568
rect 12687 9537 12699 9540
rect 12641 9531 12699 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12912 9577 12940 9608
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13814 9568 13820 9580
rect 13587 9540 13820 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14918 9568 14924 9580
rect 14691 9540 14924 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 13630 9500 13636 9512
rect 3007 9472 4292 9500
rect 10888 9472 11560 9500
rect 13591 9472 13636 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 2682 9392 2688 9444
rect 2740 9392 2746 9444
rect 4264 9441 4292 9472
rect 11532 9441 11560 9472
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 13771 9472 14841 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 15286 9500 15292 9512
rect 15247 9472 15292 9500
rect 14829 9463 14887 9469
rect 4249 9435 4307 9441
rect 4249 9401 4261 9435
rect 4295 9401 4307 9435
rect 4249 9395 4307 9401
rect 11517 9435 11575 9441
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 2317 9367 2375 9373
rect 2317 9333 2329 9367
rect 2363 9364 2375 9367
rect 2498 9364 2504 9376
rect 2363 9336 2504 9364
rect 2363 9333 2375 9336
rect 2317 9327 2375 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 6457 9367 6515 9373
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 7558 9364 7564 9376
rect 6503 9336 7564 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9582 9364 9588 9376
rect 9539 9336 9588 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 11532 9364 11560 9395
rect 13740 9364 13768 9463
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 11532 9336 13768 9364
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 3234 9160 3240 9172
rect 2188 9132 3240 9160
rect 2188 9120 2194 9132
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 4062 9160 4068 9172
rect 4019 9132 4068 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4338 9160 4344 9172
rect 4203 9132 4344 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4172 9092 4200 9123
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8938 9160 8944 9172
rect 8168 9132 8944 9160
rect 8168 9120 8174 9132
rect 8938 9120 8944 9132
rect 8996 9160 9002 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 8996 9132 9505 9160
rect 8996 9120 9002 9132
rect 9493 9129 9505 9132
rect 9539 9160 9551 9163
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9539 9132 9965 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9953 9129 9965 9132
rect 9999 9160 10011 9163
rect 10134 9160 10140 9172
rect 9999 9132 10140 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10134 9120 10140 9132
rect 10192 9160 10198 9172
rect 10686 9160 10692 9172
rect 10192 9132 10692 9160
rect 10192 9120 10198 9132
rect 10686 9120 10692 9132
rect 10744 9160 10750 9172
rect 10744 9132 11560 9160
rect 10744 9120 10750 9132
rect 10042 9092 10048 9104
rect 3344 9064 4200 9092
rect 10003 9064 10048 9092
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3344 9033 3372 9064
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 8993 3387 9027
rect 3329 8987 3387 8993
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 4154 9024 4160 9036
rect 3559 8996 4160 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 2700 8956 2728 8987
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 11532 9033 11560 9132
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13688 9132 14105 9160
rect 13688 9120 13694 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14918 9160 14924 9172
rect 14879 9132 14924 9160
rect 14093 9123 14151 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 12860 9064 12909 9092
rect 12860 9052 12866 9064
rect 12897 9061 12909 9064
rect 12943 9092 12955 9095
rect 13906 9092 13912 9104
rect 12943 9064 13912 9092
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 13906 9052 13912 9064
rect 13964 9092 13970 9104
rect 13964 9064 14780 9092
rect 13964 9052 13970 9064
rect 14752 9033 14780 9064
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5776 8996 5917 9024
rect 5776 8984 5782 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 11517 9027 11575 9033
rect 11517 8993 11529 9027
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 9024 14795 9027
rect 15102 9024 15108 9036
rect 14783 8996 15108 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 4433 8959 4491 8965
rect 2700 8928 4384 8956
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 3050 8888 3056 8900
rect 2455 8860 3056 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 4062 8888 4068 8900
rect 3283 8860 4068 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 4356 8888 4384 8928
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 5736 8956 5764 8984
rect 4479 8928 5764 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5994 8916 6000 8968
rect 6052 8956 6058 8968
rect 11330 8956 11336 8968
rect 6052 8928 11336 8956
rect 6052 8916 6058 8928
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8956 11483 8959
rect 11532 8956 11560 8987
rect 11471 8928 11560 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 11773 8959 11831 8965
rect 11773 8956 11785 8959
rect 11664 8928 11785 8956
rect 11664 8916 11670 8928
rect 11773 8925 11785 8928
rect 11819 8956 11831 8959
rect 13096 8956 13124 8987
rect 15102 8984 15108 8996
rect 15160 9024 15166 9036
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 15160 8996 15485 9024
rect 15160 8984 15166 8996
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 14918 8956 14924 8968
rect 11819 8928 14924 8956
rect 11819 8925 11831 8928
rect 11773 8919 11831 8925
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15746 8956 15752 8968
rect 15427 8928 15752 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 4678 8891 4736 8897
rect 4678 8888 4690 8891
rect 4356 8860 4690 8888
rect 4678 8857 4690 8860
rect 4724 8888 4736 8891
rect 5534 8888 5540 8900
rect 4724 8860 5540 8888
rect 4724 8857 4736 8860
rect 4678 8851 4736 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 6150 8891 6208 8897
rect 6150 8888 6162 8891
rect 5828 8860 6162 8888
rect 2869 8823 2927 8829
rect 2869 8789 2881 8823
rect 2915 8820 2927 8823
rect 3142 8820 3148 8832
rect 2915 8792 3148 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 5828 8829 5856 8860
rect 6150 8857 6162 8860
rect 6196 8857 6208 8891
rect 6150 8851 6208 8857
rect 11180 8891 11238 8897
rect 11180 8857 11192 8891
rect 11226 8888 11238 8891
rect 12066 8888 12072 8900
rect 11226 8860 12072 8888
rect 11226 8857 11238 8860
rect 11180 8851 11238 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 12768 8860 13369 8888
rect 12768 8848 12774 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 14642 8888 14648 8900
rect 13403 8860 14648 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5684 8792 5825 8820
rect 5684 8780 5690 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 7282 8820 7288 8832
rect 7243 8792 7288 8820
rect 5813 8783 5871 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 12860 8792 13277 8820
rect 12860 8780 12866 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13722 8820 13728 8832
rect 13683 8792 13728 8820
rect 13265 8783 13323 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14458 8820 14464 8832
rect 14419 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14608 8792 14653 8820
rect 14608 8780 14614 8792
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 1811 8588 2237 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2225 8585 2237 8588
rect 2271 8616 2283 8619
rect 2314 8616 2320 8628
rect 2271 8588 2320 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 3142 8616 3148 8628
rect 3103 8588 3148 8616
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3292 8588 3985 8616
rect 3292 8576 3298 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 5534 8616 5540 8628
rect 5495 8588 5540 8616
rect 3973 8579 4031 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 10686 8616 10692 8628
rect 10647 8588 10692 8616
rect 10686 8576 10692 8588
rect 10744 8616 10750 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 10744 8588 11529 8616
rect 10744 8576 10750 8588
rect 11517 8585 11529 8588
rect 11563 8616 11575 8619
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11563 8588 12081 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12710 8616 12716 8628
rect 12671 8588 12716 8616
rect 12069 8579 12127 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13722 8616 13728 8628
rect 13403 8588 13728 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 13872 8588 13917 8616
rect 13872 8576 13878 8588
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 14056 8588 14105 8616
rect 14056 8576 14062 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14550 8616 14556 8628
rect 14415 8588 14556 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 2130 8548 2136 8560
rect 2091 8520 2136 8548
rect 2130 8508 2136 8520
rect 2188 8508 2194 8560
rect 3053 8551 3111 8557
rect 3053 8517 3065 8551
rect 3099 8548 3111 8551
rect 3418 8548 3424 8560
rect 3099 8520 3424 8548
rect 3099 8517 3111 8520
rect 3053 8511 3111 8517
rect 3418 8508 3424 8520
rect 3476 8548 3482 8560
rect 3786 8548 3792 8560
rect 3476 8520 3792 8548
rect 3476 8508 3482 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 5813 8551 5871 8557
rect 5813 8548 5825 8551
rect 4172 8520 5825 8548
rect 3878 8480 3884 8492
rect 3344 8452 3884 8480
rect 3344 8421 3372 8452
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4172 8489 4200 8520
rect 5813 8517 5825 8520
rect 5859 8548 5871 8551
rect 5997 8551 6055 8557
rect 5997 8548 6009 8551
rect 5859 8520 6009 8548
rect 5859 8517 5871 8520
rect 5813 8511 5871 8517
rect 5997 8517 6009 8520
rect 6043 8548 6055 8551
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 6043 8520 6193 8548
rect 6043 8517 6055 8520
rect 5997 8511 6055 8517
rect 6181 8517 6193 8520
rect 6227 8548 6239 8551
rect 7190 8548 7196 8560
rect 6227 8520 7196 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 7190 8508 7196 8520
rect 7248 8548 7254 8560
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 7248 8520 7389 8548
rect 7248 8508 7254 8520
rect 7377 8517 7389 8520
rect 7423 8548 7435 8551
rect 7423 8520 8892 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4413 8483 4471 8489
rect 4413 8480 4425 8483
rect 4157 8443 4215 8449
rect 4264 8452 4425 8480
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8381 2099 8415
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 2041 8375 2099 8381
rect 2240 8384 3341 8412
rect 2056 8344 2084 8375
rect 2240 8344 2268 8384
rect 3329 8381 3341 8384
rect 3375 8381 3387 8415
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3329 8375 3387 8381
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 4264 8412 4292 8452
rect 4413 8449 4425 8452
rect 4459 8449 4471 8483
rect 4413 8443 4471 8449
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 8864 8489 8892 8520
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 13449 8551 13507 8557
rect 13449 8548 13461 8551
rect 13320 8520 13461 8548
rect 13320 8508 13326 8520
rect 13449 8517 13461 8520
rect 13495 8548 13507 8551
rect 13538 8548 13544 8560
rect 13495 8520 13544 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13538 8508 13544 8520
rect 13596 8548 13602 8560
rect 13909 8551 13967 8557
rect 13909 8548 13921 8551
rect 13596 8520 13921 8548
rect 13596 8508 13602 8520
rect 13909 8517 13921 8520
rect 13955 8517 13967 8551
rect 14108 8548 14136 8579
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14826 8616 14832 8628
rect 14787 8588 14832 8616
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 15746 8616 15752 8628
rect 15703 8588 15752 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 14108 8520 14749 8548
rect 13909 8511 13967 8517
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 8582 8483 8640 8489
rect 8582 8480 8594 8483
rect 7524 8452 8594 8480
rect 7524 8440 7530 8452
rect 8582 8449 8594 8452
rect 8628 8449 8640 8483
rect 8582 8443 8640 8449
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 8938 8480 8944 8492
rect 8895 8452 8944 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 9214 8489 9220 8492
rect 9208 8443 9220 8489
rect 9272 8480 9278 8492
rect 9272 8452 9308 8480
rect 9214 8440 9220 8443
rect 9272 8440 9278 8452
rect 3620 8384 4292 8412
rect 13265 8415 13323 8421
rect 2056 8316 2268 8344
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 3620 8344 3648 8384
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13906 8412 13912 8424
rect 13311 8384 13912 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 14976 8384 15021 8412
rect 14976 8372 14982 8384
rect 2464 8316 3648 8344
rect 2464 8304 2470 8316
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 7156 8316 7481 8344
rect 7156 8304 7162 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 11790 8344 11796 8356
rect 10367 8316 11796 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 2685 8279 2743 8285
rect 2685 8276 2697 8279
rect 2556 8248 2697 8276
rect 2556 8236 2562 8248
rect 2685 8245 2697 8248
rect 2731 8245 2743 8279
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 2685 8239 2743 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 10962 8276 10968 8288
rect 5408 8248 10968 8276
rect 5408 8236 5414 8248
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11606 8276 11612 8288
rect 11112 8248 11612 8276
rect 11112 8236 11118 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14366 8276 14372 8288
rect 13872 8248 14372 8276
rect 13872 8236 13878 8248
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 3142 8072 3148 8084
rect 2823 8044 3148 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 7190 8072 7196 8084
rect 7151 8044 7196 8072
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8072 9002 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8996 8044 9137 8072
rect 8996 8032 9002 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2406 7936 2412 7948
rect 2271 7908 2412 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3476 7908 3525 7936
rect 3476 7896 3482 7908
rect 3513 7905 3525 7908
rect 3559 7936 3571 7939
rect 3896 7936 3924 8032
rect 3559 7908 3924 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7208 7936 7236 8032
rect 6972 7908 7236 7936
rect 8665 7939 8723 7945
rect 6972 7896 6978 7908
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 9140 7936 9168 8035
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12124 8044 12265 8072
rect 12124 8032 12130 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 13814 8072 13820 8084
rect 13775 8044 13820 8072
rect 12253 8035 12311 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14458 8072 14464 8084
rect 14419 8044 14464 8072
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 15746 8072 15752 8084
rect 15703 8044 15752 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 12161 8007 12219 8013
rect 12161 7973 12173 8007
rect 12207 8004 12219 8007
rect 12618 8004 12624 8016
rect 12207 7976 12624 8004
rect 12207 7973 12219 7976
rect 12161 7967 12219 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 14274 8004 14280 8016
rect 14187 7976 14280 8004
rect 14274 7964 14280 7976
rect 14332 8004 14338 8016
rect 14734 8004 14740 8016
rect 14332 7976 14740 8004
rect 14332 7964 14338 7976
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8711 7908 9321 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 5166 7868 5172 7880
rect 1995 7840 5172 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5307 7840 5457 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5445 7837 5457 7840
rect 5491 7868 5503 7871
rect 6932 7868 6960 7896
rect 5491 7840 6960 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 8398 7871 8456 7877
rect 8398 7868 8410 7871
rect 7340 7840 8410 7868
rect 7340 7828 7346 7840
rect 8398 7837 8410 7840
rect 8444 7837 8456 7871
rect 9324 7868 9352 7899
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15013 7939 15071 7945
rect 15013 7936 15025 7939
rect 14976 7908 15025 7936
rect 14976 7896 14982 7908
rect 15013 7905 15025 7908
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 9858 7868 9864 7880
rect 9324 7840 9864 7868
rect 8398 7831 8456 7837
rect 9858 7828 9864 7840
rect 9916 7868 9922 7880
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 9916 7840 10793 7868
rect 9916 7828 9922 7840
rect 10781 7837 10793 7840
rect 10827 7868 10839 7871
rect 11330 7868 11336 7880
rect 10827 7840 11336 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 11330 7828 11336 7840
rect 11388 7868 11394 7880
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 11388 7840 13645 7868
rect 11388 7828 11394 7840
rect 13633 7837 13645 7840
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14550 7868 14556 7880
rect 13872 7840 14556 7868
rect 13872 7828 13878 7840
rect 14550 7828 14556 7840
rect 14608 7868 14614 7880
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 14608 7840 14841 7868
rect 14608 7828 14614 7840
rect 14829 7837 14841 7840
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 2317 7803 2375 7809
rect 2317 7769 2329 7803
rect 2363 7800 2375 7803
rect 3329 7803 3387 7809
rect 2363 7772 2912 7800
rect 2363 7769 2375 7772
rect 2317 7763 2375 7769
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2884 7741 2912 7772
rect 3329 7769 3341 7803
rect 3375 7800 3387 7803
rect 3970 7800 3976 7812
rect 3375 7772 3976 7800
rect 3375 7769 3387 7772
rect 3329 7763 3387 7769
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 5016 7803 5074 7809
rect 5016 7800 5028 7803
rect 4212 7772 5028 7800
rect 4212 7760 4218 7772
rect 5016 7769 5028 7772
rect 5062 7800 5074 7803
rect 5062 7772 5672 7800
rect 5062 7769 5074 7772
rect 5016 7763 5074 7769
rect 2869 7735 2927 7741
rect 2464 7704 2509 7732
rect 2464 7692 2470 7704
rect 2869 7701 2881 7735
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 4246 7732 4252 7744
rect 3283 7704 4252 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 5537 7735 5595 7741
rect 5537 7732 5549 7735
rect 5500 7704 5549 7732
rect 5500 7692 5506 7704
rect 5537 7701 5549 7704
rect 5583 7701 5595 7735
rect 5644 7732 5672 7772
rect 5718 7760 5724 7812
rect 5776 7800 5782 7812
rect 9582 7809 9588 7812
rect 6672 7803 6730 7809
rect 6672 7800 6684 7803
rect 5776 7772 6684 7800
rect 5776 7760 5782 7772
rect 6672 7769 6684 7772
rect 6718 7800 6730 7803
rect 9576 7800 9588 7809
rect 6718 7772 7328 7800
rect 9543 7772 9588 7800
rect 6718 7769 6730 7772
rect 6672 7763 6730 7769
rect 7006 7732 7012 7744
rect 5644 7704 7012 7732
rect 5537 7695 5595 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7300 7741 7328 7772
rect 9576 7763 9588 7772
rect 9582 7760 9588 7763
rect 9640 7760 9646 7812
rect 11048 7803 11106 7809
rect 11048 7800 11060 7803
rect 10704 7772 11060 7800
rect 10704 7741 10732 7772
rect 11048 7769 11060 7772
rect 11094 7800 11106 7803
rect 11094 7772 12434 7800
rect 11094 7769 11106 7772
rect 11048 7763 11106 7769
rect 7285 7735 7343 7741
rect 7285 7701 7297 7735
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7701 10747 7735
rect 12406 7732 12434 7772
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 13078 7800 13084 7812
rect 12676 7772 13084 7800
rect 12676 7760 12682 7772
rect 13078 7760 13084 7772
rect 13136 7800 13142 7812
rect 13366 7803 13424 7809
rect 13366 7800 13378 7803
rect 13136 7772 13378 7800
rect 13136 7760 13142 7772
rect 13366 7769 13378 7772
rect 13412 7769 13424 7803
rect 15102 7800 15108 7812
rect 13366 7763 13424 7769
rect 13740 7772 15108 7800
rect 13740 7732 13768 7772
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 12406 7704 13768 7732
rect 14921 7735 14979 7741
rect 10689 7695 10747 7701
rect 14921 7701 14933 7735
rect 14967 7732 14979 7735
rect 15010 7732 15016 7744
rect 14967 7704 15016 7732
rect 14967 7701 14979 7704
rect 14921 7695 14979 7701
rect 15010 7692 15016 7704
rect 15068 7732 15074 7744
rect 15194 7732 15200 7744
rect 15068 7704 15200 7732
rect 15068 7692 15074 7704
rect 15194 7692 15200 7704
rect 15252 7732 15258 7744
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 15252 7704 15301 7732
rect 15252 7692 15258 7704
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2777 7531 2835 7537
rect 2777 7528 2789 7531
rect 2464 7500 2789 7528
rect 2464 7488 2470 7500
rect 2777 7497 2789 7500
rect 2823 7497 2835 7531
rect 2777 7491 2835 7497
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3510 7528 3516 7540
rect 3191 7500 3516 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 5718 7528 5724 7540
rect 3752 7500 5724 7528
rect 3752 7488 3758 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5859 7500 6101 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 6089 7497 6101 7500
rect 6135 7528 6147 7531
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6135 7500 6653 7528
rect 6135 7497 6147 7500
rect 6089 7491 6147 7497
rect 6641 7497 6653 7500
rect 6687 7528 6699 7531
rect 6914 7528 6920 7540
rect 6687 7500 6920 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 1673 7463 1731 7469
rect 1673 7460 1685 7463
rect 1636 7432 1685 7460
rect 1636 7420 1642 7432
rect 1673 7429 1685 7432
rect 1719 7429 1731 7463
rect 1673 7423 1731 7429
rect 2746 7432 5672 7460
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2746 7392 2774 7432
rect 1995 7364 2774 7392
rect 3237 7395 3295 7401
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3326 7392 3332 7404
rect 3283 7364 3332 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3326 7352 3332 7364
rect 3384 7392 3390 7404
rect 3384 7364 3924 7392
rect 3384 7352 3390 7364
rect 3896 7336 3924 7364
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4028 7364 4073 7392
rect 4028 7352 4034 7364
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 5442 7392 5448 7404
rect 5500 7401 5506 7404
rect 4212 7364 5448 7392
rect 4212 7352 4218 7364
rect 5442 7352 5448 7364
rect 5500 7355 5512 7401
rect 5500 7352 5506 7355
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3936 7296 4077 7324
rect 3936 7284 3942 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 5644 7324 5672 7432
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 5828 7392 5856 7491
rect 6748 7401 6776 7500
rect 6914 7488 6920 7500
rect 6972 7488 6978 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 7064 7500 8217 7528
rect 7064 7488 7070 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 8205 7491 8263 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 12989 7531 13047 7537
rect 12989 7528 13001 7531
rect 9968 7500 13001 7528
rect 6840 7432 9536 7460
rect 5767 7364 5856 7392
rect 6733 7395 6791 7401
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6840 7324 6868 7432
rect 7006 7401 7012 7404
rect 7000 7355 7012 7401
rect 7064 7392 7070 7404
rect 7064 7364 7100 7392
rect 7006 7352 7012 7355
rect 7064 7352 7070 7364
rect 9306 7352 9312 7404
rect 9364 7401 9370 7404
rect 9364 7392 9376 7401
rect 9364 7364 9409 7392
rect 9364 7355 9376 7364
rect 9364 7352 9370 7355
rect 5644 7296 6868 7324
rect 9508 7324 9536 7432
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 9876 7392 9904 7488
rect 9631 7364 9904 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 9968 7324 9996 7500
rect 12989 7497 13001 7500
rect 13035 7497 13047 7531
rect 12989 7491 13047 7497
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 13964 7500 14197 7528
rect 13964 7488 13970 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 14185 7491 14243 7497
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14332 7500 14377 7528
rect 14332 7488 14338 7500
rect 14826 7488 14832 7540
rect 14884 7528 14890 7540
rect 15197 7531 15255 7537
rect 15197 7528 15209 7531
rect 14884 7500 15209 7528
rect 14884 7488 14890 7500
rect 15197 7497 15209 7500
rect 15243 7528 15255 7531
rect 15746 7528 15752 7540
rect 15243 7500 15752 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 11790 7469 11796 7472
rect 11784 7460 11796 7469
rect 11751 7432 11796 7460
rect 11784 7423 11796 7432
rect 11848 7460 11854 7472
rect 12802 7460 12808 7472
rect 11848 7432 12808 7460
rect 11790 7420 11796 7423
rect 11848 7420 11854 7432
rect 12802 7420 12808 7432
rect 12860 7420 12866 7472
rect 11054 7392 11060 7404
rect 11112 7401 11118 7404
rect 11024 7364 11060 7392
rect 11054 7352 11060 7364
rect 11112 7355 11124 7401
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11112 7352 11118 7355
rect 11330 7352 11336 7364
rect 11388 7392 11394 7404
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 11388 7364 11529 7392
rect 11388 7352 11394 7364
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 13357 7395 13415 7401
rect 12124 7364 13032 7392
rect 12124 7352 12130 7364
rect 9508 7296 9996 7324
rect 4065 7287 4123 7293
rect 3789 7259 3847 7265
rect 3789 7225 3801 7259
rect 3835 7256 3847 7259
rect 4246 7256 4252 7268
rect 3835 7228 4252 7256
rect 3835 7225 3847 7228
rect 3789 7219 3847 7225
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 12894 7256 12900 7268
rect 9640 7228 10088 7256
rect 12855 7228 12900 7256
rect 9640 7216 9646 7228
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4430 7188 4436 7200
rect 4387 7160 4436 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 7006 7188 7012 7200
rect 5868 7160 7012 7188
rect 5868 7148 5874 7160
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7892 7160 8125 7188
rect 7892 7148 7898 7160
rect 8113 7157 8125 7160
rect 8159 7188 8171 7191
rect 8202 7188 8208 7200
rect 8159 7160 8208 7188
rect 8159 7157 8171 7160
rect 8113 7151 8171 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 9950 7188 9956 7200
rect 9911 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10060 7188 10088 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13004 7256 13032 7364
rect 13357 7361 13369 7395
rect 13403 7392 13415 7395
rect 13722 7392 13728 7404
rect 13403 7364 13728 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15378 7392 15384 7404
rect 15151 7364 15384 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 13446 7324 13452 7336
rect 13407 7296 13452 7324
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 13556 7256 13584 7287
rect 14384 7256 14412 7287
rect 13004 7228 13584 7256
rect 13648 7228 14412 7256
rect 13648 7188 13676 7228
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 15304 7256 15332 7287
rect 15160 7228 15332 7256
rect 15160 7216 15166 7228
rect 13814 7188 13820 7200
rect 10060 7160 13676 7188
rect 13775 7160 13820 7188
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15565 7191 15623 7197
rect 15565 7188 15577 7191
rect 15344 7160 15577 7188
rect 15344 7148 15350 7160
rect 15565 7157 15577 7160
rect 15611 7157 15623 7191
rect 15565 7151 15623 7157
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9858 6984 9864 6996
rect 9079 6956 9864 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 3510 6876 3516 6928
rect 3568 6916 3574 6928
rect 3970 6916 3976 6928
rect 3568 6888 3976 6916
rect 3568 6876 3574 6888
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 7285 6919 7343 6925
rect 7285 6885 7297 6919
rect 7331 6885 7343 6919
rect 7285 6879 7343 6885
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 4172 6848 4200 6876
rect 3467 6820 4200 6848
rect 7300 6848 7328 6879
rect 8757 6851 8815 6857
rect 7300 6820 7788 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4424 6783 4482 6789
rect 4424 6749 4436 6783
rect 4470 6749 4482 6783
rect 4424 6743 4482 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 7760 6780 7788 6820
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8846 6848 8852 6860
rect 8803 6820 8852 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8846 6808 8852 6820
rect 8904 6848 8910 6860
rect 9048 6848 9076 6947
rect 9858 6944 9864 6956
rect 9916 6984 9922 6996
rect 10321 6987 10379 6993
rect 10321 6984 10333 6987
rect 9916 6956 10333 6984
rect 9916 6944 9922 6956
rect 10321 6953 10333 6956
rect 10367 6953 10379 6987
rect 10321 6947 10379 6953
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13909 6987 13967 6993
rect 13136 6956 13400 6984
rect 13136 6944 13142 6956
rect 8904 6820 9076 6848
rect 8904 6808 8910 6820
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10870 6848 10876 6860
rect 10008 6820 10876 6848
rect 10008 6808 10014 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 13372 6848 13400 6956
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 14090 6984 14096 6996
rect 13955 6956 14096 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14090 6944 14096 6956
rect 14148 6984 14154 6996
rect 14550 6984 14556 6996
rect 14148 6956 14556 6984
rect 14148 6944 14154 6956
rect 14550 6944 14556 6956
rect 14608 6984 14614 6996
rect 14608 6956 15056 6984
rect 14608 6944 14614 6956
rect 13725 6919 13783 6925
rect 13725 6885 13737 6919
rect 13771 6916 13783 6919
rect 13998 6916 14004 6928
rect 13771 6888 14004 6916
rect 13771 6885 13783 6888
rect 13725 6879 13783 6885
rect 13998 6876 14004 6888
rect 14056 6916 14062 6928
rect 14458 6916 14464 6928
rect 14056 6888 14464 6916
rect 14056 6876 14062 6888
rect 14458 6876 14464 6888
rect 14516 6876 14522 6928
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 13372 6820 14657 6848
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 15028 6848 15056 6956
rect 15102 6876 15108 6928
rect 15160 6916 15166 6928
rect 15160 6888 15516 6916
rect 15160 6876 15166 6888
rect 15488 6857 15516 6888
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15028 6820 15393 6848
rect 14645 6811 14703 6817
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 9398 6780 9404 6792
rect 7760 6752 9404 6780
rect 5905 6743 5963 6749
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3142 6644 3148 6656
rect 2832 6616 2877 6644
rect 3103 6616 3148 6644
rect 2832 6604 2838 6616
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3418 6644 3424 6656
rect 3283 6616 3424 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4172 6644 4200 6743
rect 4338 6672 4344 6724
rect 4396 6712 4402 6724
rect 4448 6712 4476 6743
rect 5920 6712 5948 6743
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11388 6752 11897 6780
rect 11388 6740 11394 6752
rect 11885 6749 11897 6752
rect 11931 6780 11943 6783
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 11931 6752 13369 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13357 6743 13415 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13906 6780 13912 6792
rect 13648 6752 13912 6780
rect 4396 6684 4476 6712
rect 4540 6684 5948 6712
rect 4396 6672 4402 6684
rect 4540 6644 4568 6684
rect 5534 6644 5540 6656
rect 4172 6616 4568 6644
rect 5495 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5813 6647 5871 6653
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 5920 6644 5948 6684
rect 6172 6715 6230 6721
rect 6172 6681 6184 6715
rect 6218 6712 6230 6715
rect 8512 6715 8570 6721
rect 6218 6684 8432 6712
rect 6218 6681 6230 6684
rect 6172 6675 6230 6681
rect 6454 6644 6460 6656
rect 5859 6616 6460 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7466 6644 7472 6656
rect 7423 6616 7472 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7466 6604 7472 6616
rect 7524 6644 7530 6656
rect 8110 6644 8116 6656
rect 7524 6616 8116 6644
rect 7524 6604 7530 6616
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8404 6644 8432 6684
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 11238 6712 11244 6724
rect 8558 6684 11244 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11618 6715 11676 6721
rect 11618 6712 11630 6715
rect 11348 6684 11630 6712
rect 9766 6644 9772 6656
rect 8404 6616 9772 6644
rect 9766 6604 9772 6616
rect 9824 6644 9830 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 9824 6616 10517 6644
rect 9824 6604 9830 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11348 6644 11376 6684
rect 11618 6681 11630 6684
rect 11664 6681 11676 6715
rect 11618 6675 11676 6681
rect 11900 6684 12848 6712
rect 11900 6656 11928 6684
rect 10928 6616 11376 6644
rect 10928 6604 10934 6616
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 11977 6647 12035 6653
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12526 6644 12532 6656
rect 12023 6616 12532 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12820 6644 12848 6684
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13090 6715 13148 6721
rect 13090 6712 13102 6715
rect 12952 6684 13102 6712
rect 12952 6672 12958 6684
rect 13090 6681 13102 6684
rect 13136 6712 13148 6715
rect 13648 6712 13676 6752
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14734 6780 14740 6792
rect 14507 6752 14740 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 13136 6684 13676 6712
rect 13136 6681 13148 6684
rect 13090 6675 13148 6681
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 13780 6684 13952 6712
rect 13780 6672 13786 6684
rect 13538 6644 13544 6656
rect 12820 6616 13544 6644
rect 13538 6604 13544 6616
rect 13596 6604 13602 6656
rect 13924 6644 13952 6684
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13924 6616 14105 6644
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14608 6616 14653 6644
rect 14608 6604 14614 6616
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14792 6616 14933 6644
rect 14792 6604 14798 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 15286 6644 15292 6656
rect 15247 6616 15292 6644
rect 14921 6607 14979 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2961 6443 3019 6449
rect 2740 6400 2774 6440
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3878 6440 3884 6452
rect 3007 6412 3884 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3878 6400 3884 6412
rect 3936 6440 3942 6452
rect 6086 6440 6092 6452
rect 3936 6412 6092 6440
rect 3936 6400 3942 6412
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 9122 6440 9128 6452
rect 6236 6412 9128 6440
rect 6236 6400 6242 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11388 6412 11529 6440
rect 11388 6400 11394 6412
rect 11517 6409 11529 6412
rect 11563 6440 11575 6443
rect 11790 6440 11796 6452
rect 11563 6412 11796 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13219 6412 13737 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13872 6412 14197 6440
rect 13872 6400 13878 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14185 6403 14243 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 15378 6440 15384 6452
rect 15339 6412 15384 6440
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 2746 6372 2774 6400
rect 8846 6372 8852 6384
rect 2746 6344 4660 6372
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6304 2007 6307
rect 2774 6304 2780 6316
rect 1995 6276 2780 6304
rect 1995 6273 2007 6276
rect 1949 6267 2007 6273
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 3878 6304 3884 6316
rect 2915 6276 3884 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4430 6264 4436 6316
rect 4488 6313 4494 6316
rect 4488 6304 4500 6313
rect 4488 6276 4533 6304
rect 4488 6267 4500 6276
rect 4488 6264 4494 6267
rect 1670 6236 1676 6248
rect 1631 6208 1676 6236
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 4632 6236 4660 6344
rect 4816 6344 6500 6372
rect 4816 6313 4844 6344
rect 6472 6316 6500 6344
rect 7208 6344 8852 6372
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4755 6276 4813 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 5057 6307 5115 6313
rect 5057 6304 5069 6307
rect 4801 6267 4859 6273
rect 4908 6276 5069 6304
rect 4908 6236 4936 6276
rect 5057 6273 5069 6276
rect 5103 6304 5115 6307
rect 5534 6304 5540 6316
rect 5103 6276 5540 6304
rect 5103 6273 5115 6276
rect 5057 6267 5115 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6454 6304 6460 6316
rect 6367 6276 6460 6304
rect 6454 6264 6460 6276
rect 6512 6304 6518 6316
rect 7208 6313 7236 6344
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 6512 6276 6653 6304
rect 6512 6264 6518 6276
rect 6641 6273 6653 6276
rect 6687 6304 6699 6307
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6687 6276 7113 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 7101 6273 7113 6276
rect 7147 6304 7159 6307
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 7147 6276 7205 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7460 6307 7518 6313
rect 7460 6273 7472 6307
rect 7506 6304 7518 6307
rect 7926 6304 7932 6316
rect 7506 6276 7932 6304
rect 7506 6273 7518 6276
rect 7460 6267 7518 6273
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 8680 6313 8708 6344
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 14734 6372 14740 6384
rect 13311 6344 14740 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 15010 6372 15016 6384
rect 14844 6344 15016 6372
rect 8938 6313 8944 6316
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8932 6304 8944 6313
rect 8899 6276 8944 6304
rect 8665 6267 8723 6273
rect 8932 6267 8944 6276
rect 8938 6264 8944 6267
rect 8996 6264 9002 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13872 6276 14105 6304
rect 13872 6264 13878 6276
rect 14093 6273 14105 6276
rect 14139 6304 14151 6307
rect 14844 6304 14872 6344
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 14139 6276 14872 6304
rect 14921 6307 14979 6313
rect 14139 6273 14151 6276
rect 14093 6267 14151 6273
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15470 6304 15476 6316
rect 14967 6276 15476 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 13078 6236 13084 6248
rect 3191 6208 3372 6236
rect 4632 6208 4936 6236
rect 13039 6208 13084 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 3344 6109 3372 6208
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 13504 6140 13645 6168
rect 13504 6128 13510 6140
rect 13633 6137 13645 6140
rect 13679 6137 13691 6171
rect 13633 6131 13691 6137
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14090 6168 14096 6180
rect 13780 6140 14096 6168
rect 13780 6128 13786 6140
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 14384 6168 14412 6199
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 15013 6239 15071 6245
rect 15013 6236 15025 6239
rect 14700 6208 15025 6236
rect 14700 6196 14706 6208
rect 15013 6205 15025 6208
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15160 6208 15205 6236
rect 15160 6196 15166 6208
rect 15120 6168 15148 6196
rect 14384 6140 15148 6168
rect 3329 6103 3387 6109
rect 3329 6069 3341 6103
rect 3375 6100 3387 6103
rect 4338 6100 4344 6112
rect 3375 6072 4344 6100
rect 3375 6069 3387 6072
rect 3329 6063 3387 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8260 6072 8585 6100
rect 8260 6060 8266 6072
rect 8573 6069 8585 6072
rect 8619 6100 8631 6103
rect 8938 6100 8944 6112
rect 8619 6072 8944 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9732 6072 10057 6100
rect 9732 6060 9738 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 12894 6060 12900 6112
rect 12952 6100 12958 6112
rect 13998 6100 14004 6112
rect 12952 6072 14004 6100
rect 12952 6060 12958 6072
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 3418 5896 3424 5908
rect 3379 5868 3424 5896
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 5810 5896 5816 5908
rect 5771 5868 5816 5896
rect 5810 5856 5816 5868
rect 5868 5896 5874 5908
rect 6270 5896 6276 5908
rect 5868 5868 6276 5896
rect 5868 5856 5874 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 8294 5896 8300 5908
rect 8207 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5896 8358 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 8352 5868 8585 5896
rect 8352 5856 8358 5868
rect 8573 5865 8585 5868
rect 8619 5896 8631 5899
rect 8846 5896 8852 5908
rect 8619 5868 8852 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8846 5856 8852 5868
rect 8904 5896 8910 5908
rect 9585 5899 9643 5905
rect 9585 5896 9597 5899
rect 8904 5868 9597 5896
rect 8904 5856 8910 5868
rect 9585 5865 9597 5868
rect 9631 5865 9643 5899
rect 11238 5896 11244 5908
rect 11199 5868 11244 5896
rect 9585 5859 9643 5865
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5760 2191 5763
rect 2222 5760 2228 5772
rect 2179 5732 2228 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 2056 5692 2084 5723
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 3694 5760 3700 5772
rect 2915 5732 3700 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 3878 5760 3884 5772
rect 3839 5732 3884 5760
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8294 5760 8300 5772
rect 7239 5732 8300 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9600 5760 9628 5859
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 11348 5868 12817 5896
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11149 5831 11207 5837
rect 11149 5828 11161 5831
rect 11112 5800 11161 5828
rect 11112 5788 11118 5800
rect 11149 5797 11161 5800
rect 11195 5797 11207 5831
rect 11149 5791 11207 5797
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9600 5732 9781 5760
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 4062 5692 4068 5704
rect 2056 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4295 5664 4353 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 5718 5692 5724 5704
rect 4387 5664 5724 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 5718 5652 5724 5664
rect 5776 5692 5782 5704
rect 6454 5692 6460 5704
rect 5776 5664 6460 5692
rect 5776 5652 5782 5664
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6937 5695 6995 5701
rect 6937 5661 6949 5695
rect 6983 5692 6995 5695
rect 7098 5692 7104 5704
rect 6983 5664 7104 5692
rect 6983 5661 6995 5664
rect 6937 5655 6995 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 11348 5692 11376 5868
rect 12805 5865 12817 5868
rect 12851 5896 12863 5899
rect 13630 5896 13636 5908
rect 12851 5868 13636 5896
rect 12851 5865 12863 5868
rect 12805 5859 12863 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 14182 5896 14188 5908
rect 14095 5868 14188 5896
rect 14182 5856 14188 5868
rect 14240 5896 14246 5908
rect 14734 5896 14740 5908
rect 14240 5868 14740 5896
rect 14240 5856 14246 5868
rect 14734 5856 14740 5868
rect 14792 5896 14798 5908
rect 14918 5896 14924 5908
rect 14792 5868 14924 5896
rect 14792 5856 14798 5868
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15470 5896 15476 5908
rect 15431 5868 15476 5896
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 13648 5828 13676 5856
rect 14369 5831 14427 5837
rect 14369 5828 14381 5831
rect 13648 5800 14381 5828
rect 14369 5797 14381 5800
rect 14415 5828 14427 5831
rect 14642 5828 14648 5840
rect 14415 5800 14648 5828
rect 14415 5797 14427 5800
rect 14369 5791 14427 5797
rect 14642 5788 14648 5800
rect 14700 5788 14706 5840
rect 15194 5760 15200 5772
rect 15155 5732 15200 5760
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 7708 5664 11376 5692
rect 7708 5652 7714 5664
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11848 5664 12633 5692
rect 11848 5652 11854 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5692 13691 5695
rect 14458 5692 14464 5704
rect 13679 5664 14464 5692
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 3053 5627 3111 5633
rect 3053 5624 3065 5627
rect 2746 5596 3065 5624
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 2406 5556 2412 5568
rect 2271 5528 2412 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2593 5559 2651 5565
rect 2593 5525 2605 5559
rect 2639 5556 2651 5559
rect 2746 5556 2774 5596
rect 3053 5593 3065 5596
rect 3099 5593 3111 5627
rect 4586 5627 4644 5633
rect 4586 5624 4598 5627
rect 3053 5587 3111 5593
rect 3528 5596 4598 5624
rect 2958 5556 2964 5568
rect 2639 5528 2774 5556
rect 2919 5528 2964 5556
rect 2639 5525 2651 5528
rect 2593 5519 2651 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 3528 5565 3556 5596
rect 4586 5593 4598 5596
rect 4632 5593 4644 5627
rect 4586 5587 4644 5593
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 7282 5624 7288 5636
rect 5408 5596 7288 5624
rect 5408 5584 5414 5596
rect 7282 5584 7288 5596
rect 7340 5584 7346 5636
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 9122 5624 9128 5636
rect 7515 5596 9128 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 3513 5559 3571 5565
rect 3513 5556 3525 5559
rect 3476 5528 3525 5556
rect 3476 5516 3482 5528
rect 3513 5525 3525 5528
rect 3559 5525 3571 5559
rect 3513 5519 3571 5525
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 5368 5556 5396 5584
rect 4120 5528 5396 5556
rect 5721 5559 5779 5565
rect 4120 5516 4126 5528
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 7006 5556 7012 5568
rect 5767 5528 7012 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 7484 5556 7512 5587
rect 9122 5584 9128 5596
rect 9180 5584 9186 5636
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10014 5627 10072 5633
rect 10014 5624 10026 5627
rect 9732 5596 10026 5624
rect 9732 5584 9738 5596
rect 10014 5593 10026 5596
rect 10060 5593 10072 5627
rect 10014 5587 10072 5593
rect 12376 5627 12434 5633
rect 12376 5593 12388 5627
rect 12422 5624 12434 5627
rect 12526 5624 12532 5636
rect 12422 5596 12532 5624
rect 12422 5593 12434 5596
rect 12376 5587 12434 5593
rect 12526 5584 12532 5596
rect 12584 5584 12590 5636
rect 14936 5624 14964 5655
rect 12636 5596 14964 5624
rect 7248 5528 7512 5556
rect 7248 5516 7254 5528
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 9858 5556 9864 5568
rect 7984 5528 9864 5556
rect 7984 5516 7990 5528
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 12636 5556 12664 5596
rect 10192 5528 12664 5556
rect 10192 5516 10198 5528
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 13136 5528 13737 5556
rect 13136 5516 13142 5528
rect 13725 5525 13737 5528
rect 13771 5556 13783 5559
rect 13814 5556 13820 5568
rect 13771 5528 13820 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5321 2283 5355
rect 2225 5315 2283 5321
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2240 5216 2268 5315
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2869 5355 2927 5361
rect 2869 5352 2881 5355
rect 2372 5324 2881 5352
rect 2372 5312 2378 5324
rect 2869 5321 2881 5324
rect 2915 5321 2927 5355
rect 2869 5315 2927 5321
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3513 5355 3571 5361
rect 3513 5352 3525 5355
rect 3016 5324 3525 5352
rect 3016 5312 3022 5324
rect 3513 5321 3525 5324
rect 3559 5321 3571 5355
rect 3513 5315 3571 5321
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4019 5324 4629 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5224 5324 5457 5352
rect 5224 5312 5230 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 6454 5352 6460 5364
rect 6415 5324 6460 5352
rect 5445 5315 5503 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6914 5312 6920 5364
rect 6972 5312 6978 5364
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5352 7067 5355
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7055 5324 7389 5352
rect 7055 5321 7067 5324
rect 7009 5315 7067 5321
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 9858 5352 9864 5364
rect 9815 5324 9864 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 10686 5352 10692 5364
rect 10284 5324 10692 5352
rect 10284 5312 10290 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 11790 5352 11796 5364
rect 11195 5324 11796 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 14182 5352 14188 5364
rect 13311 5324 14188 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 2590 5284 2596 5296
rect 2551 5256 2596 5284
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 3234 5244 3240 5296
rect 3292 5284 3298 5296
rect 3881 5287 3939 5293
rect 3881 5284 3893 5287
rect 3292 5256 3893 5284
rect 3292 5244 3298 5256
rect 3881 5253 3893 5256
rect 3927 5284 3939 5287
rect 4341 5287 4399 5293
rect 4341 5284 4353 5287
rect 3927 5256 4353 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4341 5253 4353 5256
rect 4387 5284 4399 5287
rect 4798 5284 4804 5296
rect 4387 5256 4804 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 6932 5284 6960 5312
rect 7834 5284 7840 5296
rect 6932 5256 7840 5284
rect 7834 5244 7840 5256
rect 7892 5284 7898 5296
rect 8634 5287 8692 5293
rect 8634 5284 8646 5287
rect 7892 5256 8646 5284
rect 7892 5244 7898 5256
rect 8634 5253 8646 5256
rect 8680 5253 8692 5287
rect 8634 5247 8692 5253
rect 13357 5287 13415 5293
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 13630 5284 13636 5296
rect 13403 5256 13636 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 13630 5244 13636 5256
rect 13688 5244 13694 5296
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2240 5188 2329 5216
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 2317 5179 2375 5185
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 2464 5188 3157 5216
rect 2464 5176 2470 5188
rect 3145 5185 3157 5188
rect 3191 5216 3203 5219
rect 3326 5216 3332 5228
rect 3191 5188 3332 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 4246 5176 4252 5228
rect 4304 5216 4310 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4304 5188 4997 5216
rect 4304 5176 4310 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 5810 5216 5816 5228
rect 5771 5188 5816 5216
rect 4985 5179 5043 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 6963 5188 7043 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5117 1639 5151
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1581 5111 1639 5117
rect 1596 5012 1624 5111
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 4062 5148 4068 5160
rect 4023 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 5074 5148 5080 5160
rect 5035 5120 5080 5148
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5626 5148 5632 5160
rect 5307 5120 5632 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5902 5148 5908 5160
rect 5863 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6730 5148 6736 5160
rect 6135 5120 6736 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 6178 5040 6184 5092
rect 6236 5040 6242 5092
rect 7015 5080 7043 5188
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7524 5188 7757 5216
rect 7524 5176 7530 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7852 5188 8064 5216
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7374 5148 7380 5160
rect 7156 5120 7380 5148
rect 7156 5108 7162 5120
rect 7374 5108 7380 5120
rect 7432 5108 7438 5160
rect 7190 5080 7196 5092
rect 7015 5052 7196 5080
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 6196 5012 6224 5040
rect 1596 4984 6224 5012
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6512 4984 6561 5012
rect 6512 4972 6518 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 7760 5012 7788 5179
rect 7852 5157 7880 5188
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 8036 5148 8064 5188
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8352 5188 8401 5216
rect 8352 5176 8358 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 9214 5216 9220 5228
rect 8389 5179 8447 5185
rect 8496 5188 9220 5216
rect 8496 5148 8524 5188
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5216 10287 5219
rect 11514 5216 11520 5228
rect 10275 5188 11520 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 13170 5216 13176 5228
rect 12483 5188 13176 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13872 5188 14105 5216
rect 13872 5176 13878 5188
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14139 5188 14749 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 8036 5120 8524 5148
rect 10321 5151 10379 5157
rect 7929 5111 7987 5117
rect 10321 5117 10333 5151
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 11974 5148 11980 5160
rect 11935 5120 11980 5148
rect 10413 5111 10471 5117
rect 7944 5080 7972 5111
rect 8110 5080 8116 5092
rect 7944 5052 8116 5080
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 9456 5052 10088 5080
rect 9456 5040 9462 5052
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7760 4984 8217 5012
rect 6549 4975 6607 4981
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10060 5012 10088 5052
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10336 5080 10364 5111
rect 10284 5052 10364 5080
rect 10284 5040 10290 5052
rect 10428 5012 10456 5111
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12526 5148 12532 5160
rect 12487 5120 12532 5148
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 12636 5080 12664 5111
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 14182 5148 14188 5160
rect 13504 5120 13549 5148
rect 14143 5120 14188 5148
rect 13504 5108 13510 5120
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 11296 5052 12664 5080
rect 11296 5040 11302 5052
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 14292 5080 14320 5111
rect 14642 5080 14648 5092
rect 13964 5052 14648 5080
rect 13964 5040 13970 5052
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 12066 5012 12072 5024
rect 9916 4984 9961 5012
rect 10060 4984 10456 5012
rect 12027 4984 12072 5012
rect 9916 4972 9922 4984
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12216 4984 12909 5012
rect 12216 4972 12222 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 13688 4984 13737 5012
rect 13688 4972 13694 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 13725 4975 13783 4981
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14550 5012 14556 5024
rect 14240 4984 14556 5012
rect 14240 4972 14246 4984
rect 14550 4972 14556 4984
rect 14608 5012 14614 5024
rect 14918 5012 14924 5024
rect 14608 4984 14924 5012
rect 14608 4972 14614 4984
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1857 4811 1915 4817
rect 1857 4808 1869 4811
rect 1820 4780 1869 4808
rect 1820 4768 1826 4780
rect 1857 4777 1869 4780
rect 1903 4777 1915 4811
rect 1857 4771 1915 4777
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3142 4808 3148 4820
rect 2915 4780 3148 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5258 4808 5264 4820
rect 4948 4780 5264 4808
rect 4948 4768 4954 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5718 4808 5724 4820
rect 5679 4780 5724 4808
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5960 4780 6193 4808
rect 5960 4768 5966 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 6420 4780 9137 4808
rect 6420 4768 6426 4780
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 2188 4712 3801 4740
rect 2188 4700 2194 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 3789 4703 3847 4709
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 5442 4740 5448 4752
rect 4304 4712 5448 4740
rect 4304 4700 4310 4712
rect 5442 4700 5448 4712
rect 5500 4740 5506 4752
rect 5813 4743 5871 4749
rect 5813 4740 5825 4743
rect 5500 4712 5825 4740
rect 5500 4700 5506 4712
rect 5813 4709 5825 4712
rect 5859 4709 5871 4743
rect 5813 4703 5871 4709
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6328 4712 6776 4740
rect 6328 4700 6334 4712
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2682 4672 2688 4684
rect 2547 4644 2688 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3694 4672 3700 4684
rect 3559 4644 3700 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 4338 4672 4344 4684
rect 4251 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4672 4402 4684
rect 4614 4672 4620 4684
rect 4396 4644 4620 4672
rect 4396 4632 4402 4644
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5902 4672 5908 4684
rect 5132 4644 5908 4672
rect 5132 4632 5138 4644
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6748 4681 6776 4712
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6733 4675 6791 4681
rect 6733 4641 6745 4675
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7300 4681 7328 4780
rect 9125 4777 9137 4780
rect 9171 4808 9183 4811
rect 9950 4808 9956 4820
rect 9171 4780 9956 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 10284 4780 10333 4808
rect 10284 4768 10290 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 10321 4771 10379 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 13170 4808 13176 4820
rect 13131 4780 13176 4808
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 15013 4811 15071 4817
rect 15013 4777 15025 4811
rect 15059 4808 15071 4811
rect 15102 4808 15108 4820
rect 15059 4780 15108 4808
rect 15059 4777 15071 4780
rect 15013 4771 15071 4777
rect 8573 4743 8631 4749
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 9398 4740 9404 4752
rect 8619 4712 9404 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 10870 4700 10876 4752
rect 10928 4740 10934 4752
rect 10928 4712 12434 4740
rect 10928 4700 10934 4712
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 7064 4644 7113 4672
rect 7064 4632 7070 4644
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8202 4672 8208 4684
rect 8067 4644 8208 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9214 4672 9220 4684
rect 8803 4644 9220 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4672 9830 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 9824 4644 12081 4672
rect 9824 4632 9830 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12406 4672 12434 4712
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 12676 4712 13768 4740
rect 12676 4700 12682 4712
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12406 4644 13001 4672
rect 12069 4635 12127 4641
rect 12989 4641 13001 4644
rect 13035 4672 13047 4675
rect 13446 4672 13452 4684
rect 13035 4644 13452 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13740 4681 13768 4712
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4641 13783 4675
rect 14642 4672 14648 4684
rect 14603 4644 14648 4672
rect 13725 4635 13783 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 4430 4604 4436 4616
rect 2271 4576 4436 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 7024 4576 7389 4604
rect 7024 4548 7052 4576
rect 7377 4573 7389 4576
rect 7423 4604 7435 4607
rect 7742 4604 7748 4616
rect 7423 4576 7748 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 7800 4576 8953 4604
rect 7800 4564 7806 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 11974 4564 11980 4616
rect 12032 4604 12038 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12032 4576 12725 4604
rect 12032 4564 12038 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 13354 4604 13360 4616
rect 12851 4576 13360 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15028 4604 15056 4771
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 14608 4576 15056 4604
rect 14608 4564 14614 4576
rect 3237 4539 3295 4545
rect 3237 4505 3249 4539
rect 3283 4536 3295 4539
rect 3786 4536 3792 4548
rect 3283 4508 3792 4536
rect 3283 4505 3295 4508
rect 3237 4499 3295 4505
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 4172 4508 4629 4536
rect 4172 4480 4200 4508
rect 4617 4505 4629 4508
rect 4663 4505 4675 4539
rect 4617 4499 4675 4505
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 4856 4508 6960 4536
rect 4856 4496 4862 4508
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 4154 4468 4160 4480
rect 3384 4440 3429 4468
rect 4115 4440 4160 4468
rect 3384 4428 3390 4440
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 4338 4468 4344 4480
rect 4295 4440 4344 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4338 4428 4344 4440
rect 4396 4468 4402 4480
rect 4890 4468 4896 4480
rect 4396 4440 4896 4468
rect 4396 4428 4402 4440
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5074 4468 5080 4480
rect 5035 4440 5080 4468
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5902 4468 5908 4480
rect 5583 4440 5908 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6512 4440 6561 4468
rect 6512 4428 6518 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6932 4468 6960 4508
rect 7006 4496 7012 4548
rect 7064 4496 7070 4548
rect 9582 4536 9588 4548
rect 7116 4508 9588 4536
rect 7116 4468 7144 4508
rect 9582 4496 9588 4508
rect 9640 4536 9646 4548
rect 11333 4539 11391 4545
rect 11333 4536 11345 4539
rect 9640 4508 11345 4536
rect 9640 4496 9646 4508
rect 11333 4505 11345 4508
rect 11379 4536 11391 4539
rect 11790 4536 11796 4548
rect 11379 4508 11796 4536
rect 11379 4505 11391 4508
rect 11333 4499 11391 4505
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 11885 4539 11943 4545
rect 11885 4505 11897 4539
rect 11931 4536 11943 4539
rect 13541 4539 13599 4545
rect 11931 4508 12388 4536
rect 11931 4505 11943 4508
rect 11885 4499 11943 4505
rect 7742 4468 7748 4480
rect 6932 4440 7144 4468
rect 7703 4440 7748 4468
rect 6549 4431 6607 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 8076 4440 8125 4468
rect 8076 4428 8082 4440
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8294 4468 8300 4480
rect 8251 4440 8300 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 9858 4468 9864 4480
rect 9819 4440 9864 4468
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 11057 4471 11115 4477
rect 10008 4440 10053 4468
rect 10008 4428 10014 4440
rect 11057 4437 11069 4471
rect 11103 4468 11115 4471
rect 11146 4468 11152 4480
rect 11103 4440 11152 4468
rect 11103 4437 11115 4440
rect 11057 4431 11115 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12158 4468 12164 4480
rect 12023 4440 12164 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12360 4477 12388 4508
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 13587 4508 14136 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 14108 4477 14136 4508
rect 12345 4471 12403 4477
rect 12345 4437 12357 4471
rect 12391 4437 12403 4471
rect 12345 4431 12403 4437
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1854 4264 1860 4276
rect 1719 4236 1860 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2041 4267 2099 4273
rect 2041 4233 2053 4267
rect 2087 4264 2099 4267
rect 2498 4264 2504 4276
rect 2087 4236 2504 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4264 3019 4267
rect 3326 4264 3332 4276
rect 3007 4236 3332 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3786 4224 3792 4276
rect 3844 4264 3850 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 3844 4236 4629 4264
rect 3844 4224 3850 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 4617 4227 4675 4233
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5074 4264 5080 4276
rect 5031 4236 5080 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5074 4224 5080 4236
rect 5132 4224 5138 4276
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 5316 4236 5457 4264
rect 5316 4224 5322 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5445 4227 5503 4233
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 5813 4267 5871 4273
rect 5813 4264 5825 4267
rect 5684 4236 5825 4264
rect 5684 4224 5690 4236
rect 5813 4233 5825 4236
rect 5859 4264 5871 4267
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 5859 4236 6469 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 6457 4233 6469 4236
rect 6503 4264 6515 4267
rect 7466 4264 7472 4276
rect 6503 4236 7472 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7800 4236 7941 4264
rect 7800 4224 7806 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4264 8079 4267
rect 8110 4264 8116 4276
rect 8067 4236 8116 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8389 4267 8447 4273
rect 8389 4264 8401 4267
rect 8352 4236 8401 4264
rect 8352 4224 8358 4236
rect 8389 4233 8401 4236
rect 8435 4233 8447 4267
rect 9398 4264 9404 4276
rect 9359 4236 9404 4264
rect 8389 4227 8447 4233
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 9858 4224 9864 4276
rect 9916 4264 9922 4276
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 9916 4236 10333 4264
rect 9916 4224 9922 4236
rect 10321 4233 10333 4236
rect 10367 4233 10379 4267
rect 10321 4227 10379 4233
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 10735 4236 11529 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11517 4227 11575 4233
rect 11790 4224 11796 4276
rect 11848 4264 11854 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11848 4236 11989 4264
rect 11848 4224 11854 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 12805 4267 12863 4273
rect 12805 4264 12817 4267
rect 12768 4236 12817 4264
rect 12768 4224 12774 4236
rect 12805 4233 12817 4236
rect 12851 4264 12863 4267
rect 13265 4267 13323 4273
rect 13265 4264 13277 4267
rect 12851 4236 13277 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 13265 4233 13277 4236
rect 13311 4264 13323 4267
rect 13354 4264 13360 4276
rect 13311 4236 13360 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 3970 4196 3976 4208
rect 3344 4168 3976 4196
rect 3344 4140 3372 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 5534 4196 5540 4208
rect 5092 4168 5540 4196
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2869 4131 2927 4137
rect 2188 4100 2233 4128
rect 2188 4088 2194 4100
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3326 4128 3332 4140
rect 2915 4100 3332 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3602 4128 3608 4140
rect 3467 4100 3608 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4982 4128 4988 4140
rect 4203 4100 4988 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2682 4060 2688 4072
rect 2363 4032 2688 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3970 4060 3976 4072
rect 3559 4032 3976 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 2222 3952 2228 4004
rect 2280 3992 2286 4004
rect 4172 3992 4200 4091
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5092 4137 5120 4168
rect 5534 4156 5540 4168
rect 5592 4196 5598 4208
rect 6086 4196 6092 4208
rect 5592 4168 6092 4196
rect 5592 4156 5598 4168
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 8128 4128 8156 4224
rect 9493 4199 9551 4205
rect 9493 4165 9505 4199
rect 9539 4196 9551 4199
rect 9766 4196 9772 4208
rect 9539 4168 9772 4196
rect 9539 4165 9551 4168
rect 9493 4159 9551 4165
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4196 11299 4199
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11287 4168 11897 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 11885 4165 11897 4168
rect 11931 4196 11943 4199
rect 13630 4196 13636 4208
rect 11931 4168 13636 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 5951 4100 6684 4128
rect 8128 4100 8493 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4522 4060 4528 4072
rect 4479 4032 4528 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 2280 3964 4200 3992
rect 2280 3952 2286 3964
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4264 3924 4292 4023
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4060 5227 4063
rect 5350 4060 5356 4072
rect 5215 4032 5356 4060
rect 5215 4029 5227 4032
rect 5169 4023 5227 4029
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 4540 3992 4568 4020
rect 6012 3992 6040 4023
rect 6656 4001 6684 4100
rect 8481 4097 8493 4100
rect 8527 4128 8539 4131
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8527 4100 8677 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8665 4097 8677 4100
rect 8711 4128 8723 4131
rect 8711 4100 11192 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 7190 4060 7196 4072
rect 7151 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 7926 4060 7932 4072
rect 7883 4032 7932 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9674 4060 9680 4072
rect 9355 4032 9680 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11164 4060 11192 4100
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12216 4100 12633 4128
rect 12216 4088 12222 4100
rect 12621 4097 12633 4100
rect 12667 4128 12679 4131
rect 12894 4128 12900 4140
rect 12667 4100 12900 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 13078 4128 13084 4140
rect 12952 4100 13084 4128
rect 12952 4088 12958 4100
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 11790 4060 11796 4072
rect 10928 4032 10973 4060
rect 11164 4032 11796 4060
rect 10928 4020 10934 4032
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 4540 3964 6040 3992
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 8386 3992 8392 4004
rect 6687 3964 8392 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 8386 3952 8392 3964
rect 8444 3992 8450 4004
rect 9214 3992 9220 4004
rect 8444 3964 9220 3992
rect 8444 3952 8450 3964
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9861 3995 9919 4001
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 10134 3992 10140 4004
rect 9907 3964 10140 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11882 3992 11888 4004
rect 11112 3964 11888 3992
rect 11112 3952 11118 3964
rect 11882 3952 11888 3964
rect 11940 3992 11946 4004
rect 12084 3992 12112 4023
rect 11940 3964 12112 3992
rect 11940 3952 11946 3964
rect 7098 3924 7104 3936
rect 4028 3896 7104 3924
rect 4028 3884 4034 3896
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11974 3924 11980 3936
rect 11204 3896 11980 3924
rect 11204 3884 11210 3896
rect 11974 3884 11980 3896
rect 12032 3924 12038 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12032 3896 12357 3924
rect 12032 3884 12038 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2372 3692 2697 3720
rect 2372 3680 2378 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 3234 3720 3240 3732
rect 2685 3683 2743 3689
rect 2976 3692 3240 3720
rect 2866 3652 2872 3664
rect 2056 3624 2872 3652
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1636 3556 1777 3584
rect 1636 3544 1642 3556
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2056 3525 2084 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3485 2099 3519
rect 2041 3479 2099 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2976 3516 3004 3692
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3602 3720 3608 3732
rect 3563 3692 3608 3720
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 3970 3720 3976 3732
rect 3931 3692 3976 3720
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 4430 3720 4436 3732
rect 4391 3692 4436 3720
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 5040 3692 5273 3720
rect 5040 3680 5046 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 5166 3652 5172 3664
rect 3160 3624 5172 3652
rect 3160 3593 3188 3624
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 5276 3652 5304 3683
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5868 3692 6009 3720
rect 5868 3680 5874 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 6512 3692 7849 3720
rect 6512 3680 6518 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 7837 3683 7895 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 10008 3692 10517 3720
rect 10008 3680 10014 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 10836 3692 11345 3720
rect 10836 3680 10842 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 12526 3720 12532 3732
rect 12207 3692 12532 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 7742 3652 7748 3664
rect 5276 3624 6868 3652
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3553 3203 3587
rect 3145 3547 3203 3553
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 4614 3584 4620 3596
rect 3375 3556 4620 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 4614 3544 4620 3556
rect 4672 3584 4678 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4672 3556 4997 3584
rect 4672 3544 4678 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 5626 3584 5632 3596
rect 4985 3547 5043 3553
rect 5092 3556 5632 3584
rect 5092 3528 5120 3556
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6270 3544 6276 3596
rect 6328 3584 6334 3596
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 6328 3556 6561 3584
rect 6328 3544 6334 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 2639 3488 3004 3516
rect 3053 3519 3111 3525
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3786 3516 3792 3528
rect 3099 3488 3792 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4847 3488 5028 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 2314 3448 2320 3460
rect 2275 3420 2320 3448
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 2608 3420 4200 3448
rect 2608 3392 2636 3420
rect 2590 3340 2596 3392
rect 2648 3340 2654 3392
rect 4172 3389 4200 3420
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3349 4215 3383
rect 4356 3380 4384 3479
rect 5000 3460 5028 3488
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3516 5595 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5583 3488 5917 3516
rect 5583 3485 5595 3488
rect 5537 3479 5595 3485
rect 5905 3485 5917 3488
rect 5951 3516 5963 3519
rect 5994 3516 6000 3528
rect 5951 3488 6000 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6840 3516 6868 3624
rect 7300 3624 7748 3652
rect 7300 3593 7328 3624
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 8294 3612 8300 3664
rect 8352 3652 8358 3664
rect 8352 3624 9168 3652
rect 8352 3612 8358 3624
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 9140 3593 9168 3624
rect 10870 3612 10876 3664
rect 10928 3612 10934 3664
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 11514 3652 11520 3664
rect 11020 3624 11520 3652
rect 11020 3612 11026 3624
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 11606 3612 11612 3664
rect 11664 3612 11670 3664
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 12342 3652 12348 3664
rect 11756 3624 12348 3652
rect 11756 3612 11762 3624
rect 12342 3612 12348 3624
rect 12400 3652 12406 3664
rect 13817 3655 13875 3661
rect 13817 3652 13829 3655
rect 12400 3624 13829 3652
rect 12400 3612 12406 3624
rect 13817 3621 13829 3624
rect 13863 3652 13875 3655
rect 13906 3652 13912 3664
rect 13863 3624 13912 3652
rect 13863 3621 13875 3624
rect 13817 3615 13875 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7432 3556 8401 3584
rect 7432 3544 7438 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3553 9183 3587
rect 10888 3584 10916 3612
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10888 3556 11069 3584
rect 9125 3547 9183 3553
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11057 3547 11115 3553
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 11624 3584 11652 3612
rect 11882 3584 11888 3596
rect 11204 3556 11652 3584
rect 11843 3556 11888 3584
rect 11204 3544 11210 3556
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12676 3556 12725 3584
rect 12676 3544 12682 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3584 13691 3587
rect 14090 3584 14096 3596
rect 13679 3556 14096 3584
rect 13679 3553 13691 3556
rect 13633 3547 13691 3553
rect 14090 3544 14096 3556
rect 14148 3584 14154 3596
rect 14642 3584 14648 3596
rect 14148 3556 14648 3584
rect 14148 3544 14154 3556
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 7190 3516 7196 3528
rect 6840 3488 6960 3516
rect 7151 3488 7196 3516
rect 4522 3408 4528 3460
rect 4580 3448 4586 3460
rect 4893 3451 4951 3457
rect 4893 3448 4905 3451
rect 4580 3420 4905 3448
rect 4580 3408 4586 3420
rect 4893 3417 4905 3420
rect 4939 3417 4951 3451
rect 4893 3411 4951 3417
rect 4982 3408 4988 3460
rect 5040 3408 5046 3460
rect 6365 3451 6423 3457
rect 6365 3417 6377 3451
rect 6411 3448 6423 3451
rect 6932 3448 6960 3488
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7926 3516 7932 3528
rect 7524 3488 7932 3516
rect 7524 3476 7530 3488
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 8168 3488 8217 3516
rect 8168 3476 8174 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3516 10931 3519
rect 11606 3516 11612 3528
rect 10919 3488 11612 3516
rect 10919 3485 10931 3488
rect 10873 3479 10931 3485
rect 11606 3476 11612 3488
rect 11664 3516 11670 3528
rect 15286 3516 15292 3528
rect 11664 3488 15292 3516
rect 11664 3476 11670 3488
rect 15286 3476 15292 3488
rect 15344 3476 15350 3528
rect 8297 3451 8355 3457
rect 8297 3448 8309 3451
rect 6411 3420 6868 3448
rect 6932 3420 8309 3448
rect 6411 3417 6423 3420
rect 6365 3411 6423 3417
rect 5166 3380 5172 3392
rect 4356 3352 5172 3380
rect 4157 3343 4215 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 5721 3383 5779 3389
rect 5721 3380 5733 3383
rect 5684 3352 5733 3380
rect 5684 3340 5690 3352
rect 5721 3349 5733 3352
rect 5767 3349 5779 3383
rect 6454 3380 6460 3392
rect 6415 3352 6460 3380
rect 5721 3343 5779 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6840 3389 6868 3420
rect 8297 3417 8309 3420
rect 8343 3448 8355 3451
rect 8665 3451 8723 3457
rect 8665 3448 8677 3451
rect 8343 3420 8677 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 8665 3417 8677 3420
rect 8711 3448 8723 3451
rect 8938 3448 8944 3460
rect 8711 3420 8944 3448
rect 8711 3417 8723 3420
rect 8665 3411 8723 3417
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 9766 3448 9772 3460
rect 9140 3420 9772 3448
rect 6825 3383 6883 3389
rect 6825 3349 6837 3383
rect 6871 3349 6883 3383
rect 6825 3343 6883 3349
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 9140 3380 9168 3420
rect 9766 3408 9772 3420
rect 9824 3448 9830 3460
rect 9824 3420 10916 3448
rect 9824 3408 9830 3420
rect 10888 3392 10916 3420
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11793 3451 11851 3457
rect 11793 3448 11805 3451
rect 11112 3420 11805 3448
rect 11112 3408 11118 3420
rect 11793 3417 11805 3420
rect 11839 3448 11851 3451
rect 12158 3448 12164 3460
rect 11839 3420 12164 3448
rect 11839 3417 11851 3420
rect 11793 3411 11851 3417
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 12529 3451 12587 3457
rect 12529 3417 12541 3451
rect 12575 3448 12587 3451
rect 13538 3448 13544 3460
rect 12575 3420 13544 3448
rect 12575 3417 12587 3420
rect 12529 3411 12587 3417
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 9306 3380 9312 3392
rect 7616 3352 9168 3380
rect 9267 3352 9312 3380
rect 7616 3340 7622 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10134 3380 10140 3392
rect 9456 3352 9501 3380
rect 10095 3352 10140 3380
rect 9456 3340 9462 3352
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10686 3380 10692 3392
rect 10284 3352 10692 3380
rect 10284 3340 10290 3352
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 10870 3340 10876 3392
rect 10928 3340 10934 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11701 3383 11759 3389
rect 11020 3352 11065 3380
rect 11020 3340 11026 3352
rect 11701 3349 11713 3383
rect 11747 3380 11759 3383
rect 11974 3380 11980 3392
rect 11747 3352 11980 3380
rect 11747 3349 11759 3352
rect 11701 3343 11759 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12621 3383 12679 3389
rect 12621 3349 12633 3383
rect 12667 3380 12679 3383
rect 12989 3383 13047 3389
rect 12989 3380 13001 3383
rect 12667 3352 13001 3380
rect 12667 3349 12679 3352
rect 12621 3343 12679 3349
rect 12989 3349 13001 3352
rect 13035 3349 13047 3383
rect 13354 3380 13360 3392
rect 13315 3352 13360 3380
rect 12989 3343 13047 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 13504 3352 13549 3380
rect 13504 3340 13510 3352
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 3145 3179 3203 3185
rect 3145 3176 3157 3179
rect 1636 3148 3157 3176
rect 1636 3136 1642 3148
rect 3145 3145 3157 3148
rect 3191 3145 3203 3179
rect 4522 3176 4528 3188
rect 4483 3148 4528 3176
rect 3145 3139 3203 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4856 3148 4905 3176
rect 4856 3136 4862 3148
rect 4893 3145 4905 3148
rect 4939 3176 4951 3179
rect 5166 3176 5172 3188
rect 4939 3148 5172 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5534 3176 5540 3188
rect 5399 3148 5540 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6365 3179 6423 3185
rect 5776 3148 5856 3176
rect 5776 3136 5782 3148
rect 4246 3108 4252 3120
rect 3344 3080 4252 3108
rect 2038 3040 2044 3052
rect 1951 3012 2044 3040
rect 2038 3000 2044 3012
rect 2096 3040 2102 3052
rect 2222 3040 2228 3052
rect 2096 3012 2228 3040
rect 2096 3000 2102 3012
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2556 3012 2789 3040
rect 2556 3000 2562 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3344 3049 3372 3080
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 5442 3108 5448 3120
rect 4448 3080 5448 3108
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3200 3012 3341 3040
rect 3200 3000 3206 3012
rect 3329 3009 3341 3012
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 3694 3040 3700 3052
rect 3568 3012 3700 3040
rect 3568 3000 3574 3012
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4338 3040 4344 3052
rect 3844 3012 4344 3040
rect 3844 3000 3850 3012
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4448 3049 4476 3080
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 4448 2972 4476 3003
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 5828 3049 5856 3148
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6454 3176 6460 3188
rect 6411 3148 6460 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 7285 3179 7343 3185
rect 7285 3176 7297 3179
rect 6871 3148 7297 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 7285 3145 7297 3148
rect 7331 3176 7343 3179
rect 7558 3176 7564 3188
rect 7331 3148 7564 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 6178 3068 6184 3120
rect 6236 3108 6242 3120
rect 6840 3108 6868 3139
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 9122 3176 9128 3188
rect 7892 3148 9128 3176
rect 7892 3136 7898 3148
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9364 3148 9413 3176
rect 9364 3136 9370 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9815 3148 10088 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 6236 3080 6868 3108
rect 6236 3068 6242 3080
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 9950 3108 9956 3120
rect 7524 3080 9956 3108
rect 7524 3068 7530 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4672 3012 4997 3040
rect 4672 3000 4678 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5825 3043 5883 3049
rect 5031 3012 5672 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 3007 2944 4476 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4580 2944 5089 2972
rect 4580 2932 4586 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5644 2972 5672 3012
rect 5825 3009 5837 3043
rect 5871 3009 5883 3043
rect 5825 3003 5883 3009
rect 5930 3043 5988 3049
rect 5930 3009 5942 3043
rect 5976 3040 5988 3043
rect 6086 3040 6092 3052
rect 5976 3012 6092 3040
rect 5976 3009 5988 3012
rect 5930 3003 5988 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7742 3040 7748 3052
rect 7423 3012 7748 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8110 3040 8116 3052
rect 7984 3012 8116 3040
rect 7984 3000 7990 3012
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3040 9002 3052
rect 9490 3040 9496 3052
rect 8996 3012 9496 3040
rect 8996 3000 9002 3012
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9824 3012 9873 3040
rect 9824 3000 9830 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 10060 3040 10088 3148
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10192 3148 10609 3176
rect 10192 3136 10198 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11020 3148 11529 3176
rect 11020 3136 11026 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 13081 3179 13139 3185
rect 13081 3176 13093 3179
rect 12032 3148 13093 3176
rect 12032 3136 12038 3148
rect 13081 3145 13093 3148
rect 13127 3145 13139 3179
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13081 3139 13139 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13906 3176 13912 3188
rect 13596 3148 13641 3176
rect 13867 3148 13912 3176
rect 13596 3136 13602 3148
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14918 3176 14924 3188
rect 14879 3148 14924 3176
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 11885 3111 11943 3117
rect 11885 3108 11897 3111
rect 11480 3080 11897 3108
rect 11480 3068 11486 3080
rect 11885 3077 11897 3080
rect 11931 3077 11943 3111
rect 11885 3071 11943 3077
rect 12066 3068 12072 3120
rect 12124 3108 12130 3120
rect 13722 3108 13728 3120
rect 12124 3080 13728 3108
rect 12124 3068 12130 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 14826 3108 14832 3120
rect 14787 3080 14832 3108
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 10226 3040 10232 3052
rect 10060 3012 10232 3040
rect 9861 3003 9919 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10962 3040 10968 3052
rect 10735 3012 10968 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 11330 3040 11336 3052
rect 11291 3012 11336 3040
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 12618 3000 12624 3052
rect 12676 3040 12682 3052
rect 14645 3043 14703 3049
rect 12676 3012 12721 3040
rect 12676 3000 12682 3012
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14844 3040 14872 3068
rect 14691 3012 14872 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15105 3043 15163 3049
rect 15105 3040 15117 3043
rect 14976 3012 15117 3040
rect 14976 3000 14982 3012
rect 15105 3009 15117 3012
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 6362 2972 6368 2984
rect 5644 2944 6368 2972
rect 5077 2935 5135 2941
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7282 2972 7288 2984
rect 7055 2944 7288 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7834 2972 7840 2984
rect 7795 2944 7840 2972
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 8294 2972 8300 2984
rect 8067 2944 8300 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8294 2932 8300 2944
rect 8352 2972 8358 2984
rect 8846 2972 8852 2984
rect 8352 2944 8852 2972
rect 8352 2932 8358 2944
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 1210 2864 1216 2916
rect 1268 2904 1274 2916
rect 2593 2907 2651 2913
rect 2593 2904 2605 2907
rect 1268 2876 2605 2904
rect 1268 2864 1274 2876
rect 2593 2873 2605 2876
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 4249 2907 4307 2913
rect 4249 2904 4261 2907
rect 3292 2876 4261 2904
rect 3292 2864 3298 2876
rect 4249 2873 4261 2876
rect 4295 2873 4307 2907
rect 4249 2867 4307 2873
rect 5258 2864 5264 2916
rect 5316 2904 5322 2916
rect 5629 2907 5687 2913
rect 5629 2904 5641 2907
rect 5316 2876 5641 2904
rect 5316 2864 5322 2876
rect 5629 2873 5641 2876
rect 5675 2873 5687 2907
rect 5629 2867 5687 2873
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 9048 2904 9076 2935
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 10042 2972 10048 2984
rect 9180 2944 9225 2972
rect 10003 2944 10048 2972
rect 9180 2932 9186 2944
rect 10042 2932 10048 2944
rect 10100 2972 10106 2984
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10100 2944 10793 2972
rect 10100 2932 10106 2944
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11572 2944 11989 2972
rect 11572 2932 11578 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 9306 2904 9312 2916
rect 6052 2876 8800 2904
rect 9048 2876 9312 2904
rect 6052 2864 6058 2876
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2836 1915 2839
rect 1946 2836 1952 2848
rect 1903 2808 1952 2836
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 1946 2796 1952 2808
rect 2004 2796 2010 2848
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2314 2836 2320 2848
rect 2271 2808 2320 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 3510 2836 3516 2848
rect 3471 2808 3516 2836
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4154 2836 4160 2848
rect 4019 2808 4160 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 5902 2836 5908 2848
rect 5592 2808 5908 2836
rect 5592 2796 5598 2808
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6089 2839 6147 2845
rect 6089 2805 6101 2839
rect 6135 2836 6147 2839
rect 6454 2836 6460 2848
rect 6135 2808 6460 2836
rect 6135 2805 6147 2808
rect 6089 2799 6147 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7561 2839 7619 2845
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 7834 2836 7840 2848
rect 7607 2808 7840 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8772 2836 8800 2876
rect 9306 2864 9312 2876
rect 9364 2864 9370 2916
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 9456 2876 10241 2904
rect 9456 2864 9462 2876
rect 10229 2873 10241 2876
rect 10275 2873 10287 2907
rect 10229 2867 10287 2873
rect 10318 2864 10324 2916
rect 10376 2904 10382 2916
rect 10376 2876 11284 2904
rect 10376 2864 10382 2876
rect 11149 2839 11207 2845
rect 11149 2836 11161 2839
rect 8628 2808 8673 2836
rect 8772 2808 11161 2836
rect 8628 2796 8634 2808
rect 11149 2805 11161 2808
rect 11195 2805 11207 2839
rect 11256 2836 11284 2876
rect 11882 2864 11888 2916
rect 11940 2904 11946 2916
rect 12084 2904 12112 2935
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12572 2972
rect 12492 2932 12498 2944
rect 11940 2876 12112 2904
rect 11940 2864 11946 2876
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 11256 2808 12449 2836
rect 11149 2799 11207 2805
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12544 2836 12572 2944
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 12989 2975 13047 2981
rect 12860 2944 12905 2972
rect 12860 2932 12866 2944
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13078 2972 13084 2984
rect 13035 2944 13084 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13872 2944 14013 2972
rect 13872 2932 13878 2944
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14001 2935 14059 2941
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 15381 2975 15439 2981
rect 14148 2944 14193 2972
rect 14148 2932 14154 2944
rect 15381 2941 15393 2975
rect 15427 2972 15439 2975
rect 15930 2972 15936 2984
rect 15427 2944 15936 2972
rect 15427 2941 15439 2944
rect 15381 2935 15439 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 14461 2907 14519 2913
rect 14461 2873 14473 2907
rect 14507 2873 14519 2907
rect 14461 2867 14519 2873
rect 14476 2836 14504 2867
rect 12544 2808 14504 2836
rect 12437 2799 12495 2805
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 2133 2635 2191 2641
rect 2133 2632 2145 2635
rect 2096 2604 2145 2632
rect 2096 2592 2102 2604
rect 2133 2601 2145 2604
rect 2179 2601 2191 2635
rect 2133 2595 2191 2601
rect 2406 2592 2412 2644
rect 2464 2632 2470 2644
rect 2501 2635 2559 2641
rect 2501 2632 2513 2635
rect 2464 2604 2513 2632
rect 2464 2592 2470 2604
rect 2501 2601 2513 2604
rect 2547 2601 2559 2635
rect 2501 2595 2559 2601
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 3142 2632 3148 2644
rect 3099 2604 3148 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3786 2632 3792 2644
rect 3651 2604 3792 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 14918 2632 14924 2644
rect 4028 2604 14924 2632
rect 4028 2592 4034 2604
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 3694 2564 3700 2576
rect 3283 2536 3700 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 4614 2564 4620 2576
rect 4575 2536 4620 2564
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 4798 2564 4804 2576
rect 4759 2536 4804 2564
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 5534 2564 5540 2576
rect 5495 2536 5540 2564
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 5810 2564 5816 2576
rect 5771 2536 5816 2564
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2533 6055 2567
rect 5997 2527 6055 2533
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4816 2496 4844 2524
rect 4111 2468 4844 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 5166 2456 5172 2508
rect 5224 2496 5230 2508
rect 6012 2496 6040 2527
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 6917 2567 6975 2573
rect 6917 2564 6929 2567
rect 6420 2536 6929 2564
rect 6420 2524 6426 2536
rect 6917 2533 6929 2536
rect 6963 2533 6975 2567
rect 6917 2527 6975 2533
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 7558 2564 7564 2576
rect 7331 2536 7564 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 7742 2564 7748 2576
rect 7703 2536 7748 2564
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 8018 2564 8024 2576
rect 7979 2536 8024 2564
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 8110 2524 8116 2576
rect 8168 2564 8174 2576
rect 8941 2567 8999 2573
rect 8941 2564 8953 2567
rect 8168 2536 8953 2564
rect 8168 2524 8174 2536
rect 8941 2533 8953 2536
rect 8987 2533 8999 2567
rect 10870 2564 10876 2576
rect 8941 2527 8999 2533
rect 10152 2536 10364 2564
rect 10831 2536 10876 2564
rect 5224 2468 6040 2496
rect 5224 2456 5230 2468
rect 6270 2456 6276 2508
rect 6328 2496 6334 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 6328 2468 7389 2496
rect 6328 2456 6334 2468
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 3602 2428 3608 2440
rect 3467 2400 3608 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 3602 2388 3608 2400
rect 3660 2428 3666 2440
rect 4433 2431 4491 2437
rect 4433 2428 4445 2431
rect 3660 2400 4445 2428
rect 3660 2388 3666 2400
rect 4433 2397 4445 2400
rect 4479 2397 4491 2431
rect 4433 2391 4491 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5031 2400 5304 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 2498 2320 2504 2372
rect 2556 2360 2562 2372
rect 2869 2363 2927 2369
rect 2869 2360 2881 2363
rect 2556 2332 2881 2360
rect 2556 2320 2562 2332
rect 2869 2329 2881 2332
rect 2915 2360 2927 2363
rect 5074 2360 5080 2372
rect 2915 2332 5080 2360
rect 2915 2329 2927 2332
rect 2869 2323 2927 2329
rect 5074 2320 5080 2332
rect 5132 2320 5138 2372
rect 5276 2360 5304 2400
rect 5350 2388 5356 2440
rect 5408 2428 5414 2440
rect 6178 2428 6184 2440
rect 5408 2400 5453 2428
rect 6091 2400 6184 2428
rect 5408 2388 5414 2400
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 7116 2437 7144 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 7377 2459 7435 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 10042 2496 10048 2508
rect 8711 2468 10048 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 10152 2428 10180 2536
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10336 2496 10364 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 11238 2524 11244 2576
rect 11296 2564 11302 2576
rect 11296 2536 13032 2564
rect 11296 2524 11302 2536
rect 10962 2496 10968 2508
rect 10336 2468 10968 2496
rect 10229 2459 10287 2465
rect 7699 2400 10180 2428
rect 10244 2428 10272 2459
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 11112 2468 11161 2496
rect 11112 2456 11118 2468
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 12437 2499 12495 2505
rect 12437 2496 12449 2499
rect 11388 2468 12449 2496
rect 11388 2456 11394 2468
rect 12437 2465 12449 2468
rect 12483 2465 12495 2499
rect 12437 2459 12495 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12860 2468 12909 2496
rect 12860 2456 12866 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 13004 2496 13032 2536
rect 13354 2524 13360 2576
rect 13412 2564 13418 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 13412 2536 13553 2564
rect 13412 2524 13418 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 13688 2536 13733 2564
rect 13688 2524 13694 2536
rect 13814 2496 13820 2508
rect 13004 2468 13820 2496
rect 12897 2459 12955 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 10244 2400 12434 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 6196 2360 6224 2388
rect 5276 2332 6224 2360
rect 6748 2360 6776 2391
rect 7668 2360 7696 2391
rect 6748 2332 7696 2360
rect 8389 2363 8447 2369
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 8570 2360 8576 2372
rect 8435 2332 8576 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8904 2332 9137 2360
rect 8904 2320 8910 2332
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 10686 2360 10692 2372
rect 9125 2323 9183 2329
rect 10336 2332 10692 2360
rect 10336 2304 10364 2332
rect 10686 2320 10692 2332
rect 10744 2320 10750 2372
rect 11238 2360 11244 2372
rect 10796 2332 11244 2360
rect 3786 2292 3792 2304
rect 3747 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 4120 2264 4261 2292
rect 4120 2252 4126 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 4580 2264 5181 2292
rect 4580 2252 4586 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 7098 2292 7104 2304
rect 6595 2264 7104 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9364 2264 9413 2292
rect 9364 2252 9370 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9401 2255 9459 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 10318 2292 10324 2304
rect 9732 2264 9777 2292
rect 10279 2264 10324 2292
rect 9732 2252 9738 2264
rect 10318 2252 10324 2264
rect 10376 2252 10382 2304
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 10796 2301 10824 2332
rect 11238 2320 11244 2332
rect 11296 2320 11302 2372
rect 11606 2360 11612 2372
rect 11567 2332 11612 2360
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 12158 2360 12164 2372
rect 11900 2332 12164 2360
rect 11900 2304 11928 2332
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 12406 2360 12434 2400
rect 12820 2360 12848 2456
rect 13078 2428 13084 2440
rect 13039 2400 13084 2428
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13630 2428 13636 2440
rect 13219 2400 13636 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 12406 2332 12848 2360
rect 13096 2360 13124 2388
rect 13817 2363 13875 2369
rect 13817 2360 13829 2363
rect 13096 2332 13829 2360
rect 13817 2329 13829 2332
rect 13863 2329 13875 2363
rect 13817 2323 13875 2329
rect 10781 2295 10839 2301
rect 10468 2264 10513 2292
rect 10468 2252 10474 2264
rect 10781 2261 10793 2295
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11020 2264 11713 2292
rect 11020 2252 11026 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11882 2292 11888 2304
rect 11843 2264 11888 2292
rect 11701 2255 11759 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12066 2292 12072 2304
rect 12027 2264 12072 2292
rect 12066 2252 12072 2264
rect 12124 2292 12130 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12124 2264 12265 2292
rect 12124 2252 12130 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12253 2255 12311 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 12400 2264 12633 2292
rect 12400 2252 12406 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 3786 2048 3792 2100
rect 3844 2088 3850 2100
rect 5350 2088 5356 2100
rect 3844 2060 5356 2088
rect 3844 2048 3850 2060
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 10410 2088 10416 2100
rect 5500 2060 10416 2088
rect 5500 2048 5506 2060
rect 10410 2048 10416 2060
rect 10468 2048 10474 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 12066 2088 12072 2100
rect 10744 2060 12072 2088
rect 10744 2048 10750 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 11054 2020 11060 2032
rect 9272 1992 11060 2020
rect 9272 1980 9278 1992
rect 11054 1980 11060 1992
rect 11112 1980 11118 2032
rect 11606 1980 11612 2032
rect 11664 2020 11670 2032
rect 12618 2020 12624 2032
rect 11664 1992 12624 2020
rect 11664 1980 11670 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 10502 1912 10508 1964
rect 10560 1952 10566 1964
rect 11422 1952 11428 1964
rect 10560 1924 11428 1952
rect 10560 1912 10566 1924
rect 11422 1912 11428 1924
rect 11480 1952 11486 1964
rect 11882 1952 11888 1964
rect 11480 1924 11888 1952
rect 11480 1912 11486 1924
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 9122 1844 9128 1896
rect 9180 1884 9186 1896
rect 12710 1884 12716 1896
rect 9180 1856 12716 1884
rect 9180 1844 9186 1856
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 5350 1776 5356 1828
rect 5408 1816 5414 1828
rect 15010 1816 15016 1828
rect 5408 1788 15016 1816
rect 5408 1776 5414 1788
rect 15010 1776 15016 1788
rect 15068 1776 15074 1828
rect 10226 1436 10232 1488
rect 10284 1476 10290 1488
rect 14458 1476 14464 1488
rect 10284 1448 14464 1476
rect 10284 1436 10290 1448
rect 14458 1436 14464 1448
rect 14516 1436 14522 1488
<< via1 >>
rect 4068 17960 4120 18012
rect 14464 17960 14516 18012
rect 6000 17824 6052 17876
rect 11244 17824 11296 17876
rect 4068 17756 4120 17808
rect 14556 17756 14608 17808
rect 1032 17484 1084 17536
rect 12900 17688 12952 17740
rect 6184 17620 6236 17672
rect 13360 17620 13412 17672
rect 10876 17552 10928 17604
rect 14648 17552 14700 17604
rect 8392 17484 8444 17536
rect 12992 17484 13044 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 6552 17212 6604 17264
rect 7288 17280 7340 17332
rect 9772 17280 9824 17332
rect 12716 17280 12768 17332
rect 12992 17323 13044 17332
rect 12992 17289 13001 17323
rect 13001 17289 13035 17323
rect 13035 17289 13044 17323
rect 12992 17280 13044 17289
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 7748 17212 7800 17264
rect 10876 17255 10928 17264
rect 10876 17221 10885 17255
rect 10885 17221 10919 17255
rect 10919 17221 10928 17255
rect 10876 17212 10928 17221
rect 5540 17144 5592 17196
rect 4252 17076 4304 17128
rect 8576 17144 8628 17196
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 10784 17144 10836 17196
rect 9772 17076 9824 17128
rect 10876 17076 10928 17128
rect 12532 17119 12584 17128
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 7656 17008 7708 17060
rect 11796 17008 11848 17060
rect 12808 17212 12860 17264
rect 13452 17212 13504 17264
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 13820 17076 13872 17128
rect 15384 17076 15436 17128
rect 4436 16983 4488 16992
rect 4436 16949 4445 16983
rect 4445 16949 4479 16983
rect 4479 16949 4488 16983
rect 4436 16940 4488 16949
rect 4712 16940 4764 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5724 16940 5776 16992
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 7932 16940 7984 16992
rect 9220 16940 9272 16992
rect 9588 16940 9640 16992
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 11980 16940 12032 16992
rect 12624 16940 12676 16992
rect 13176 16940 13228 16992
rect 13636 17008 13688 17060
rect 14924 16940 14976 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 2964 16736 3016 16788
rect 3700 16736 3752 16788
rect 4712 16736 4764 16788
rect 5172 16736 5224 16788
rect 7748 16736 7800 16788
rect 7932 16736 7984 16788
rect 11152 16736 11204 16788
rect 12532 16736 12584 16788
rect 1768 16575 1820 16584
rect 1768 16541 1777 16575
rect 1777 16541 1811 16575
rect 1811 16541 1820 16575
rect 1768 16532 1820 16541
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 3148 16532 3200 16584
rect 3332 16575 3384 16584
rect 3332 16541 3341 16575
rect 3341 16541 3375 16575
rect 3375 16541 3384 16575
rect 3332 16532 3384 16541
rect 3240 16464 3292 16516
rect 4436 16532 4488 16584
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 6276 16668 6328 16720
rect 5264 16532 5316 16584
rect 5724 16600 5776 16652
rect 7012 16600 7064 16652
rect 8208 16600 8260 16652
rect 6000 16532 6052 16584
rect 7564 16532 7616 16584
rect 9772 16668 9824 16720
rect 9404 16600 9456 16652
rect 11704 16668 11756 16720
rect 12624 16668 12676 16720
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 9588 16575 9640 16584
rect 9588 16541 9597 16575
rect 9597 16541 9631 16575
rect 9631 16541 9640 16575
rect 9588 16532 9640 16541
rect 9956 16532 10008 16584
rect 10876 16532 10928 16584
rect 11796 16600 11848 16652
rect 12532 16600 12584 16652
rect 13452 16600 13504 16652
rect 14464 16643 14516 16652
rect 14464 16609 14473 16643
rect 14473 16609 14507 16643
rect 14507 16609 14516 16643
rect 14464 16600 14516 16609
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 11152 16532 11204 16584
rect 12440 16532 12492 16584
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 13820 16532 13872 16584
rect 1860 16396 1912 16448
rect 3608 16396 3660 16448
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 4344 16396 4396 16448
rect 5080 16396 5132 16448
rect 5816 16396 5868 16448
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 8024 16464 8076 16516
rect 6368 16396 6420 16405
rect 7932 16396 7984 16448
rect 9772 16464 9824 16516
rect 9312 16396 9364 16448
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 11980 16396 12032 16448
rect 12808 16464 12860 16516
rect 13636 16396 13688 16448
rect 14832 16464 14884 16516
rect 14648 16396 14700 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 2504 16192 2556 16244
rect 3976 16192 4028 16244
rect 7472 16192 7524 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11152 16235 11204 16244
rect 11152 16201 11161 16235
rect 11161 16201 11195 16235
rect 11195 16201 11204 16235
rect 11152 16192 11204 16201
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 11980 16235 12032 16244
rect 11980 16201 11989 16235
rect 11989 16201 12023 16235
rect 12023 16201 12032 16235
rect 11980 16192 12032 16201
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 3332 16124 3384 16176
rect 3792 16124 3844 16176
rect 4620 16124 4672 16176
rect 9312 16124 9364 16176
rect 1584 15852 1636 15904
rect 3608 16056 3660 16108
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 5172 16031 5224 16040
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5908 15988 5960 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7380 16056 7432 16108
rect 7932 16056 7984 16108
rect 8944 16056 8996 16108
rect 11244 16056 11296 16108
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12532 16124 12584 16176
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 7656 15988 7708 16040
rect 8116 16031 8168 16040
rect 8116 15997 8125 16031
rect 8125 15997 8159 16031
rect 8159 15997 8168 16031
rect 8116 15988 8168 15997
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 8852 15988 8904 16040
rect 9404 15988 9456 16040
rect 10232 15988 10284 16040
rect 9220 15920 9272 15972
rect 10876 15988 10928 16040
rect 11428 15988 11480 16040
rect 13360 16056 13412 16108
rect 3424 15852 3476 15904
rect 3608 15852 3660 15904
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 6920 15852 6972 15904
rect 7196 15852 7248 15904
rect 7380 15895 7432 15904
rect 7380 15861 7389 15895
rect 7389 15861 7423 15895
rect 7423 15861 7432 15895
rect 7380 15852 7432 15861
rect 7472 15852 7524 15904
rect 7840 15852 7892 15904
rect 8392 15852 8444 15904
rect 9956 15852 10008 15904
rect 10048 15852 10100 15904
rect 12808 15920 12860 15972
rect 12900 15920 12952 15972
rect 14464 16192 14516 16244
rect 16120 16124 16172 16176
rect 15016 16056 15068 16108
rect 14832 15988 14884 16040
rect 15752 15920 15804 15972
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 15016 15895 15068 15904
rect 12440 15852 12492 15861
rect 15016 15861 15025 15895
rect 15025 15861 15059 15895
rect 15059 15861 15068 15895
rect 15016 15852 15068 15861
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 2136 15648 2188 15700
rect 1584 15580 1636 15632
rect 6184 15648 6236 15700
rect 6368 15691 6420 15700
rect 6368 15657 6377 15691
rect 6377 15657 6411 15691
rect 6411 15657 6420 15691
rect 6368 15648 6420 15657
rect 4068 15623 4120 15632
rect 4068 15589 4077 15623
rect 4077 15589 4111 15623
rect 4111 15589 4120 15623
rect 4068 15580 4120 15589
rect 7748 15648 7800 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 10968 15648 11020 15700
rect 11704 15648 11756 15700
rect 12900 15648 12952 15700
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 3884 15512 3936 15564
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 4528 15487 4580 15496
rect 1400 15376 1452 15428
rect 4068 15376 4120 15428
rect 2780 15308 2832 15360
rect 3884 15308 3936 15360
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 5632 15512 5684 15564
rect 5724 15512 5776 15564
rect 5264 15444 5316 15496
rect 6368 15444 6420 15496
rect 10692 15580 10744 15632
rect 11520 15580 11572 15632
rect 4436 15376 4488 15428
rect 5356 15376 5408 15428
rect 6276 15376 6328 15428
rect 7564 15512 7616 15564
rect 8208 15512 8260 15564
rect 9312 15512 9364 15564
rect 8024 15444 8076 15496
rect 8392 15444 8444 15496
rect 8944 15444 8996 15496
rect 9128 15444 9180 15496
rect 10692 15444 10744 15496
rect 10968 15444 11020 15496
rect 6920 15376 6972 15428
rect 7840 15376 7892 15428
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 5448 15308 5500 15360
rect 5632 15308 5684 15360
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 7656 15308 7708 15360
rect 9220 15376 9272 15428
rect 12808 15580 12860 15632
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 13084 15512 13136 15564
rect 12440 15444 12492 15496
rect 8300 15308 8352 15360
rect 9496 15308 9548 15360
rect 10600 15308 10652 15360
rect 11244 15308 11296 15360
rect 11888 15308 11940 15360
rect 12072 15376 12124 15428
rect 12624 15308 12676 15360
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 13544 15308 13596 15360
rect 14648 15308 14700 15360
rect 15200 15308 15252 15360
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 3976 15104 4028 15156
rect 4068 15104 4120 15156
rect 4620 15104 4672 15156
rect 5632 15147 5684 15156
rect 5632 15113 5641 15147
rect 5641 15113 5675 15147
rect 5675 15113 5684 15147
rect 5632 15104 5684 15113
rect 6828 15104 6880 15156
rect 8852 15104 8904 15156
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9036 15104 9088 15113
rect 9680 15104 9732 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 11336 15104 11388 15156
rect 12072 15104 12124 15156
rect 12624 15104 12676 15156
rect 14280 15104 14332 15156
rect 3516 15011 3568 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 5448 15036 5500 15088
rect 5816 15036 5868 15088
rect 8208 15036 8260 15088
rect 8392 15079 8444 15088
rect 8392 15045 8401 15079
rect 8401 15045 8435 15079
rect 8435 15045 8444 15079
rect 8392 15036 8444 15045
rect 11152 15036 11204 15088
rect 11612 15036 11664 15088
rect 5080 14968 5132 15020
rect 7288 14968 7340 15020
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 5172 14900 5224 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 7564 14900 7616 14952
rect 8024 14943 8076 14952
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 8852 14900 8904 14952
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 11612 14900 11664 14952
rect 12808 14968 12860 15020
rect 13360 14968 13412 15020
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14740 14968 14792 15020
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 13268 14943 13320 14952
rect 12900 14900 12952 14909
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 4988 14764 5040 14816
rect 7840 14764 7892 14816
rect 8852 14764 8904 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 13268 14764 13320 14816
rect 14924 14900 14976 14952
rect 15200 14832 15252 14884
rect 15476 14900 15528 14952
rect 14464 14764 14516 14816
rect 14556 14764 14608 14816
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 4896 14603 4948 14612
rect 4896 14569 4905 14603
rect 4905 14569 4939 14603
rect 4939 14569 4948 14603
rect 4896 14560 4948 14569
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 5724 14560 5776 14612
rect 7288 14603 7340 14612
rect 7288 14569 7297 14603
rect 7297 14569 7331 14603
rect 7331 14569 7340 14603
rect 7288 14560 7340 14569
rect 7840 14560 7892 14612
rect 9496 14560 9548 14612
rect 10876 14560 10928 14612
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 1676 14467 1728 14476
rect 1676 14433 1685 14467
rect 1685 14433 1719 14467
rect 1719 14433 1728 14467
rect 1676 14424 1728 14433
rect 2688 14424 2740 14476
rect 3148 14424 3200 14476
rect 3792 14424 3844 14476
rect 2596 14356 2648 14408
rect 5264 14492 5316 14544
rect 5540 14492 5592 14544
rect 5632 14492 5684 14544
rect 5908 14424 5960 14476
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 9128 14492 9180 14544
rect 8024 14424 8076 14476
rect 9036 14424 9088 14476
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 15476 14467 15528 14476
rect 5540 14356 5592 14408
rect 3240 14220 3292 14272
rect 5816 14288 5868 14340
rect 7840 14356 7892 14408
rect 8116 14356 8168 14408
rect 11336 14356 11388 14408
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 14464 14356 14516 14365
rect 4160 14220 4212 14272
rect 4896 14220 4948 14272
rect 4988 14220 5040 14272
rect 5632 14220 5684 14272
rect 6736 14220 6788 14272
rect 12992 14288 13044 14340
rect 13912 14288 13964 14340
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 8852 14220 8904 14272
rect 9588 14220 9640 14272
rect 9864 14220 9916 14272
rect 12072 14220 12124 14272
rect 13360 14220 13412 14272
rect 14464 14220 14516 14272
rect 14648 14220 14700 14272
rect 14832 14220 14884 14272
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 3516 14016 3568 14068
rect 5172 14016 5224 14068
rect 7748 14059 7800 14068
rect 2412 13812 2464 13864
rect 3332 13880 3384 13932
rect 3608 13880 3660 13932
rect 5540 13880 5592 13932
rect 5908 13948 5960 14000
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 8300 14016 8352 14068
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 6736 13948 6788 14000
rect 9128 14016 9180 14068
rect 9496 14016 9548 14068
rect 11244 14016 11296 14068
rect 11980 14016 12032 14068
rect 12992 14016 13044 14068
rect 10876 13991 10928 14000
rect 10876 13957 10885 13991
rect 10885 13957 10919 13991
rect 10919 13957 10928 13991
rect 10876 13948 10928 13957
rect 11060 13948 11112 14000
rect 12808 13948 12860 14000
rect 13268 13948 13320 14000
rect 14556 13991 14608 14000
rect 14556 13957 14565 13991
rect 14565 13957 14599 13991
rect 14599 13957 14608 13991
rect 14556 13948 14608 13957
rect 15476 13991 15528 14000
rect 15476 13957 15485 13991
rect 15485 13957 15519 13991
rect 15519 13957 15528 13991
rect 15476 13948 15528 13957
rect 15568 13991 15620 14000
rect 15568 13957 15577 13991
rect 15577 13957 15611 13991
rect 15611 13957 15620 13991
rect 15568 13948 15620 13957
rect 9588 13880 9640 13932
rect 9956 13880 10008 13932
rect 11152 13880 11204 13932
rect 3792 13812 3844 13864
rect 3608 13744 3660 13796
rect 4160 13812 4212 13864
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 2504 13676 2556 13728
rect 5080 13676 5132 13728
rect 7380 13744 7432 13796
rect 8852 13812 8904 13864
rect 9956 13744 10008 13796
rect 10048 13744 10100 13796
rect 11336 13812 11388 13864
rect 14648 13812 14700 13864
rect 10232 13676 10284 13728
rect 13820 13676 13872 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 2688 13472 2740 13524
rect 5080 13472 5132 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 6092 13472 6144 13524
rect 7380 13472 7432 13524
rect 5908 13404 5960 13456
rect 2688 13336 2740 13388
rect 3516 13379 3568 13388
rect 3516 13345 3525 13379
rect 3525 13345 3559 13379
rect 3559 13345 3568 13379
rect 3516 13336 3568 13345
rect 2320 13268 2372 13320
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 5540 13268 5592 13320
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 3792 13200 3844 13252
rect 6460 13200 6512 13252
rect 7748 13200 7800 13252
rect 3240 13132 3292 13184
rect 10232 13472 10284 13524
rect 11612 13472 11664 13524
rect 12072 13472 12124 13524
rect 8852 13336 8904 13388
rect 9128 13336 9180 13388
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 13176 13472 13228 13524
rect 13360 13472 13412 13524
rect 14004 13472 14056 13524
rect 14832 13472 14884 13524
rect 15476 13472 15528 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 14464 13268 14516 13320
rect 14924 13268 14976 13320
rect 10140 13243 10192 13252
rect 8484 13132 8536 13184
rect 10140 13209 10174 13243
rect 10174 13209 10192 13243
rect 10140 13200 10192 13209
rect 12900 13200 12952 13252
rect 13360 13200 13412 13252
rect 13728 13200 13780 13252
rect 12532 13132 12584 13184
rect 13268 13132 13320 13184
rect 14188 13132 14240 13184
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 2320 12928 2372 12980
rect 3516 12928 3568 12980
rect 3148 12792 3200 12844
rect 3332 12860 3384 12912
rect 3792 12860 3844 12912
rect 3424 12792 3476 12844
rect 3976 12792 4028 12844
rect 4160 12792 4212 12844
rect 4620 12792 4672 12844
rect 5540 12860 5592 12912
rect 5080 12835 5132 12844
rect 5080 12801 5114 12835
rect 5114 12801 5132 12835
rect 5080 12792 5132 12801
rect 3332 12724 3384 12776
rect 7380 12928 7432 12980
rect 2596 12588 2648 12640
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 13268 12928 13320 12980
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 15016 12928 15068 12980
rect 8760 12860 8812 12912
rect 11336 12903 11388 12912
rect 9312 12792 9364 12844
rect 11336 12869 11345 12903
rect 11345 12869 11379 12903
rect 11379 12869 11388 12903
rect 11336 12860 11388 12869
rect 11612 12860 11664 12912
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 13912 12724 13964 12776
rect 14464 12724 14516 12776
rect 14740 12724 14792 12776
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 8944 12656 8996 12708
rect 12808 12656 12860 12708
rect 14188 12699 14240 12708
rect 9772 12588 9824 12640
rect 10232 12588 10284 12640
rect 11796 12588 11848 12640
rect 12164 12588 12216 12640
rect 14188 12665 14197 12699
rect 14197 12665 14231 12699
rect 14231 12665 14240 12699
rect 14188 12656 14240 12665
rect 14832 12588 14884 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 3148 12384 3200 12436
rect 3424 12384 3476 12436
rect 3976 12384 4028 12436
rect 6460 12384 6512 12436
rect 5172 12316 5224 12368
rect 5448 12316 5500 12368
rect 9128 12384 9180 12436
rect 9312 12384 9364 12436
rect 8116 12316 8168 12368
rect 10692 12384 10744 12436
rect 11612 12384 11664 12436
rect 11980 12384 12032 12436
rect 11336 12316 11388 12368
rect 4160 12248 4212 12300
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 7288 12180 7340 12232
rect 4252 12112 4304 12164
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 8760 12180 8812 12189
rect 1492 12044 1544 12096
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 3700 12044 3752 12096
rect 3976 12044 4028 12096
rect 8116 12044 8168 12096
rect 8300 12044 8352 12096
rect 9036 12044 9088 12096
rect 10876 12180 10928 12232
rect 13820 12384 13872 12436
rect 15108 12384 15160 12436
rect 14648 12248 14700 12300
rect 14832 12248 14884 12300
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 15108 12180 15160 12232
rect 9496 12112 9548 12164
rect 11428 12112 11480 12164
rect 12532 12112 12584 12164
rect 11796 12044 11848 12096
rect 11888 12044 11940 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 12992 12044 13044 12096
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 2780 11840 2832 11892
rect 3884 11840 3936 11892
rect 4160 11840 4212 11892
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 4252 11772 4304 11824
rect 9220 11840 9272 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 5172 11815 5224 11824
rect 5172 11781 5190 11815
rect 5190 11781 5224 11815
rect 5172 11772 5224 11781
rect 5540 11772 5592 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 2504 11704 2556 11756
rect 3148 11704 3200 11756
rect 4344 11704 4396 11756
rect 9036 11772 9088 11824
rect 12716 11772 12768 11824
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 2596 11500 2648 11552
rect 3884 11636 3936 11688
rect 3516 11500 3568 11552
rect 3700 11500 3752 11552
rect 5080 11500 5132 11552
rect 5264 11500 5316 11552
rect 5540 11500 5592 11552
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 7840 11500 7892 11552
rect 9864 11704 9916 11756
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 12532 11704 12584 11756
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 11612 11636 11664 11688
rect 12072 11636 12124 11688
rect 13176 11636 13228 11688
rect 10968 11568 11020 11620
rect 14648 11636 14700 11688
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13728 11500 13780 11552
rect 15568 11500 15620 11552
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 1952 11296 2004 11348
rect 5816 11339 5868 11348
rect 2504 11160 2556 11212
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 7104 11296 7156 11348
rect 7656 11296 7708 11348
rect 9404 11296 9456 11348
rect 10140 11296 10192 11348
rect 3976 11228 4028 11280
rect 4344 11271 4396 11280
rect 4344 11237 4353 11271
rect 4353 11237 4387 11271
rect 4387 11237 4396 11271
rect 4344 11228 4396 11237
rect 9036 11271 9088 11280
rect 9036 11237 9045 11271
rect 9045 11237 9079 11271
rect 9079 11237 9088 11271
rect 9036 11228 9088 11237
rect 3516 11203 3568 11212
rect 3516 11169 3525 11203
rect 3525 11169 3559 11203
rect 3559 11169 3568 11203
rect 3516 11160 3568 11169
rect 10508 11160 10560 11212
rect 10876 11296 10928 11348
rect 15292 11296 15344 11348
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 14648 11160 14700 11169
rect 3332 11135 3384 11144
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 9404 11135 9456 11144
rect 9404 11101 9438 11135
rect 9438 11101 9456 11135
rect 9404 11092 9456 11101
rect 12624 11092 12676 11144
rect 6276 11024 6328 11076
rect 2596 10956 2648 11008
rect 7840 11024 7892 11076
rect 8944 11024 8996 11076
rect 9956 11024 10008 11076
rect 10968 11024 11020 11076
rect 11888 10956 11940 11008
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 14096 10999 14148 11008
rect 12072 10956 12124 10965
rect 14096 10965 14105 10999
rect 14105 10965 14139 10999
rect 14139 10965 14148 10999
rect 14096 10956 14148 10965
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 2044 10752 2096 10804
rect 2136 10752 2188 10804
rect 5172 10752 5224 10804
rect 6276 10752 6328 10804
rect 4344 10684 4396 10736
rect 5448 10684 5500 10736
rect 5632 10684 5684 10736
rect 5816 10727 5868 10736
rect 5816 10693 5834 10727
rect 5834 10693 5868 10727
rect 5816 10684 5868 10693
rect 3424 10616 3476 10668
rect 3792 10616 3844 10668
rect 4068 10616 4120 10668
rect 7564 10659 7616 10668
rect 7564 10625 7582 10659
rect 7582 10625 7616 10659
rect 7564 10616 7616 10625
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 9036 10752 9088 10804
rect 9956 10752 10008 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 11244 10752 11296 10804
rect 12624 10795 12676 10804
rect 12624 10761 12633 10795
rect 12633 10761 12667 10795
rect 12667 10761 12676 10795
rect 12624 10752 12676 10761
rect 13360 10752 13412 10804
rect 10048 10684 10100 10736
rect 10140 10684 10192 10736
rect 12808 10684 12860 10736
rect 14096 10684 14148 10736
rect 7840 10616 7892 10625
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 3516 10548 3568 10600
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 11888 10591 11940 10600
rect 5724 10412 5776 10464
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 12532 10412 12584 10464
rect 12716 10412 12768 10464
rect 13360 10412 13412 10464
rect 14556 10412 14608 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3516 10208 3568 10260
rect 8760 10251 8812 10260
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 3884 10004 3936 10056
rect 4160 10004 4212 10056
rect 2780 9868 2832 9920
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4344 9868 4396 9920
rect 5724 10004 5776 10056
rect 8116 10004 8168 10056
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 9036 10208 9088 10260
rect 10140 10208 10192 10260
rect 11428 10208 11480 10260
rect 13820 10208 13872 10260
rect 11152 10072 11204 10124
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 7656 9979 7708 9988
rect 7656 9945 7690 9979
rect 7690 9945 7708 9979
rect 7656 9936 7708 9945
rect 9588 9936 9640 9988
rect 12072 9936 12124 9988
rect 11612 9868 11664 9920
rect 14280 9936 14332 9988
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 13636 9868 13688 9920
rect 15476 9936 15528 9988
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 8300 9664 8352 9716
rect 9588 9707 9640 9716
rect 9588 9673 9597 9707
rect 9597 9673 9631 9707
rect 9631 9673 9640 9707
rect 9588 9664 9640 9673
rect 11152 9664 11204 9716
rect 13084 9664 13136 9716
rect 14280 9707 14332 9716
rect 14280 9673 14289 9707
rect 14289 9673 14323 9707
rect 14323 9673 14332 9707
rect 14280 9664 14332 9673
rect 14556 9664 14608 9716
rect 2412 9596 2464 9648
rect 2044 9528 2096 9580
rect 2596 9528 2648 9580
rect 1400 9460 1452 9512
rect 3884 9528 3936 9580
rect 10140 9596 10192 9648
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 8208 9528 8260 9580
rect 12808 9528 12860 9580
rect 13820 9528 13872 9580
rect 14924 9528 14976 9580
rect 13636 9503 13688 9512
rect 2688 9392 2740 9444
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 15292 9503 15344 9512
rect 2504 9324 2556 9376
rect 7564 9324 7616 9376
rect 9588 9324 9640 9376
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2136 9120 2188 9172
rect 3240 9120 3292 9172
rect 4068 9120 4120 9172
rect 4344 9120 4396 9172
rect 8116 9120 8168 9172
rect 8944 9120 8996 9172
rect 10140 9120 10192 9172
rect 10692 9120 10744 9172
rect 10048 9095 10100 9104
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 10048 9061 10057 9095
rect 10057 9061 10091 9095
rect 10091 9061 10100 9095
rect 10048 9052 10100 9061
rect 4160 8984 4212 9036
rect 5724 8984 5776 9036
rect 13636 9120 13688 9172
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 12808 9052 12860 9104
rect 13912 9052 13964 9104
rect 3056 8848 3108 8900
rect 4068 8848 4120 8900
rect 6000 8916 6052 8968
rect 11336 8916 11388 8968
rect 11612 8916 11664 8968
rect 15108 8984 15160 9036
rect 14924 8916 14976 8968
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 15752 8916 15804 8968
rect 5540 8848 5592 8900
rect 3148 8780 3200 8832
rect 5632 8780 5684 8832
rect 12072 8848 12124 8900
rect 12716 8848 12768 8900
rect 14648 8848 14700 8900
rect 7288 8823 7340 8832
rect 7288 8789 7297 8823
rect 7297 8789 7331 8823
rect 7331 8789 7340 8823
rect 7288 8780 7340 8789
rect 12808 8780 12860 8832
rect 13728 8823 13780 8832
rect 13728 8789 13737 8823
rect 13737 8789 13771 8823
rect 13771 8789 13780 8823
rect 13728 8780 13780 8789
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 2320 8576 2372 8628
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 3148 8619 3200 8628
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 3240 8576 3292 8628
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 12716 8619 12768 8628
rect 12716 8585 12725 8619
rect 12725 8585 12759 8619
rect 12759 8585 12768 8619
rect 12716 8576 12768 8585
rect 13728 8576 13780 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14004 8576 14056 8628
rect 2136 8551 2188 8560
rect 2136 8517 2145 8551
rect 2145 8517 2179 8551
rect 2179 8517 2188 8551
rect 2136 8508 2188 8517
rect 3424 8508 3476 8560
rect 3792 8508 3844 8560
rect 3884 8440 3936 8492
rect 7196 8551 7248 8560
rect 7196 8517 7205 8551
rect 7205 8517 7239 8551
rect 7239 8517 7248 8551
rect 7196 8508 7248 8517
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 7472 8440 7524 8492
rect 13268 8508 13320 8560
rect 13544 8508 13596 8560
rect 14556 8576 14608 8628
rect 14832 8619 14884 8628
rect 14832 8585 14841 8619
rect 14841 8585 14875 8619
rect 14875 8585 14884 8619
rect 14832 8576 14884 8585
rect 15752 8576 15804 8628
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 9220 8483 9272 8492
rect 9220 8449 9254 8483
rect 9254 8449 9272 8483
rect 9220 8440 9272 8449
rect 2412 8304 2464 8356
rect 13912 8372 13964 8424
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 7104 8304 7156 8356
rect 11796 8304 11848 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 2504 8236 2556 8288
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 5356 8236 5408 8288
rect 10968 8236 11020 8288
rect 11060 8236 11112 8288
rect 11612 8236 11664 8288
rect 13820 8236 13872 8288
rect 14372 8236 14424 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 3148 8032 3200 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 2412 7896 2464 7948
rect 3424 7896 3476 7948
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 12072 8032 12124 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 15752 8032 15804 8084
rect 12624 7964 12676 8016
rect 14280 8007 14332 8016
rect 14280 7973 14289 8007
rect 14289 7973 14323 8007
rect 14323 7973 14332 8007
rect 14280 7964 14332 7973
rect 14740 7964 14792 8016
rect 5172 7828 5224 7880
rect 7288 7828 7340 7880
rect 14924 7896 14976 7948
rect 9864 7828 9916 7880
rect 11336 7828 11388 7880
rect 13820 7828 13872 7880
rect 14556 7828 14608 7880
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 3976 7760 4028 7812
rect 4160 7760 4212 7812
rect 2412 7692 2464 7701
rect 4252 7692 4304 7744
rect 5448 7692 5500 7744
rect 5724 7760 5776 7812
rect 9588 7803 9640 7812
rect 7012 7692 7064 7744
rect 9588 7769 9622 7803
rect 9622 7769 9640 7803
rect 9588 7760 9640 7769
rect 12624 7760 12676 7812
rect 13084 7760 13136 7812
rect 15108 7760 15160 7812
rect 15016 7692 15068 7744
rect 15200 7692 15252 7744
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 2412 7488 2464 7540
rect 3516 7488 3568 7540
rect 3700 7488 3752 7540
rect 5724 7488 5776 7540
rect 1584 7420 1636 7472
rect 3332 7352 3384 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4160 7352 4212 7404
rect 5448 7395 5500 7404
rect 5448 7361 5466 7395
rect 5466 7361 5500 7395
rect 5448 7352 5500 7361
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3884 7284 3936 7336
rect 6920 7488 6972 7540
rect 7012 7488 7064 7540
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 7012 7395 7064 7404
rect 7012 7361 7046 7395
rect 7046 7361 7064 7395
rect 7012 7352 7064 7361
rect 9312 7395 9364 7404
rect 9312 7361 9330 7395
rect 9330 7361 9364 7395
rect 9312 7352 9364 7361
rect 13912 7488 13964 7540
rect 14280 7531 14332 7540
rect 14280 7497 14289 7531
rect 14289 7497 14323 7531
rect 14323 7497 14332 7531
rect 14280 7488 14332 7497
rect 14832 7488 14884 7540
rect 15752 7488 15804 7540
rect 11796 7463 11848 7472
rect 11796 7429 11830 7463
rect 11830 7429 11848 7463
rect 11796 7420 11848 7429
rect 12808 7420 12860 7472
rect 11060 7395 11112 7404
rect 11060 7361 11078 7395
rect 11078 7361 11112 7395
rect 11060 7352 11112 7361
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 12072 7352 12124 7404
rect 4252 7216 4304 7268
rect 9588 7216 9640 7268
rect 12900 7259 12952 7268
rect 4436 7148 4488 7200
rect 5816 7148 5868 7200
rect 7012 7148 7064 7200
rect 7840 7148 7892 7200
rect 8208 7148 8260 7200
rect 9956 7191 10008 7200
rect 9956 7157 9965 7191
rect 9965 7157 9999 7191
rect 9999 7157 10008 7191
rect 9956 7148 10008 7157
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 13728 7352 13780 7404
rect 15384 7352 15436 7404
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 15108 7216 15160 7268
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15292 7148 15344 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 3516 6876 3568 6928
rect 3976 6876 4028 6928
rect 4160 6876 4212 6928
rect 8852 6808 8904 6860
rect 9864 6944 9916 6996
rect 13084 6944 13136 6996
rect 9956 6808 10008 6860
rect 10876 6808 10928 6860
rect 14096 6944 14148 6996
rect 14556 6944 14608 6996
rect 14004 6876 14056 6928
rect 14464 6876 14516 6928
rect 15108 6876 15160 6928
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 3148 6647 3200 6656
rect 2780 6604 2832 6613
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 3424 6604 3476 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4344 6672 4396 6724
rect 9404 6740 9456 6792
rect 11336 6740 11388 6792
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 6460 6604 6512 6656
rect 7472 6604 7524 6656
rect 8116 6604 8168 6656
rect 11244 6672 11296 6724
rect 9772 6604 9824 6656
rect 10876 6604 10928 6656
rect 11888 6604 11940 6656
rect 12532 6604 12584 6656
rect 12900 6672 12952 6724
rect 13912 6740 13964 6792
rect 14740 6740 14792 6792
rect 13728 6672 13780 6724
rect 13544 6604 13596 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 14740 6604 14792 6656
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 2688 6400 2740 6452
rect 3884 6400 3936 6452
rect 6092 6400 6144 6452
rect 6184 6443 6236 6452
rect 6184 6409 6193 6443
rect 6193 6409 6227 6443
rect 6227 6409 6236 6443
rect 6184 6400 6236 6409
rect 9128 6400 9180 6452
rect 11336 6400 11388 6452
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 13820 6400 13872 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 2780 6264 2832 6316
rect 3884 6264 3936 6316
rect 4436 6307 4488 6316
rect 4436 6273 4454 6307
rect 4454 6273 4488 6307
rect 4436 6264 4488 6273
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 5540 6264 5592 6316
rect 6460 6307 6512 6316
rect 6460 6273 6469 6307
rect 6469 6273 6503 6307
rect 6503 6273 6512 6307
rect 6460 6264 6512 6273
rect 7932 6264 7984 6316
rect 8852 6332 8904 6384
rect 14740 6332 14792 6384
rect 8944 6307 8996 6316
rect 8944 6273 8978 6307
rect 8978 6273 8996 6307
rect 8944 6264 8996 6273
rect 13820 6264 13872 6316
rect 15016 6332 15068 6384
rect 15476 6264 15528 6316
rect 13084 6239 13136 6248
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 13452 6128 13504 6180
rect 13728 6128 13780 6180
rect 14096 6128 14148 6180
rect 14648 6196 14700 6248
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 4344 6060 4396 6112
rect 8208 6060 8260 6112
rect 8944 6060 8996 6112
rect 9680 6060 9732 6112
rect 12900 6060 12952 6112
rect 14004 6060 14056 6112
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 5816 5899 5868 5908
rect 5816 5865 5825 5899
rect 5825 5865 5859 5899
rect 5859 5865 5868 5899
rect 5816 5856 5868 5865
rect 6276 5856 6328 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 8852 5856 8904 5908
rect 11244 5899 11296 5908
rect 2228 5720 2280 5772
rect 3700 5720 3752 5772
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 8300 5720 8352 5772
rect 11244 5865 11253 5899
rect 11253 5865 11287 5899
rect 11287 5865 11296 5899
rect 11244 5856 11296 5865
rect 11060 5788 11112 5840
rect 4068 5652 4120 5704
rect 5724 5652 5776 5704
rect 6460 5652 6512 5704
rect 7104 5652 7156 5704
rect 7656 5652 7708 5704
rect 13636 5856 13688 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 14740 5856 14792 5908
rect 14924 5856 14976 5908
rect 15476 5899 15528 5908
rect 15476 5865 15485 5899
rect 15485 5865 15519 5899
rect 15519 5865 15528 5899
rect 15476 5856 15528 5865
rect 14648 5788 14700 5840
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 11796 5652 11848 5704
rect 14464 5652 14516 5704
rect 2412 5516 2464 5568
rect 2964 5559 3016 5568
rect 2964 5525 2973 5559
rect 2973 5525 3007 5559
rect 3007 5525 3016 5559
rect 2964 5516 3016 5525
rect 3424 5516 3476 5568
rect 5356 5584 5408 5636
rect 7288 5584 7340 5636
rect 4068 5516 4120 5568
rect 7012 5516 7064 5568
rect 7196 5516 7248 5568
rect 9128 5584 9180 5636
rect 9680 5584 9732 5636
rect 12532 5584 12584 5636
rect 7932 5516 7984 5568
rect 9864 5516 9916 5568
rect 10140 5516 10192 5568
rect 13084 5516 13136 5568
rect 13820 5516 13872 5568
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2320 5312 2372 5364
rect 2964 5312 3016 5364
rect 5172 5312 5224 5364
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 6920 5312 6972 5364
rect 9864 5312 9916 5364
rect 10232 5312 10284 5364
rect 10692 5312 10744 5364
rect 11796 5312 11848 5364
rect 14188 5312 14240 5364
rect 2596 5287 2648 5296
rect 2596 5253 2605 5287
rect 2605 5253 2639 5287
rect 2639 5253 2648 5287
rect 2596 5244 2648 5253
rect 3240 5244 3292 5296
rect 4804 5244 4856 5296
rect 7840 5244 7892 5296
rect 13636 5244 13688 5296
rect 2412 5176 2464 5228
rect 3332 5176 3384 5228
rect 4252 5176 4304 5228
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 5632 5108 5684 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 6736 5108 6788 5160
rect 6184 5040 6236 5092
rect 7472 5176 7524 5228
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7380 5108 7432 5160
rect 7196 5040 7248 5092
rect 6460 4972 6512 5024
rect 8300 5176 8352 5228
rect 9220 5176 9272 5228
rect 11520 5176 11572 5228
rect 13176 5176 13228 5228
rect 13820 5176 13872 5228
rect 11980 5151 12032 5160
rect 8116 5040 8168 5092
rect 9404 5040 9456 5092
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 10232 5040 10284 5092
rect 11980 5117 11989 5151
rect 11989 5117 12023 5151
rect 12023 5117 12032 5151
rect 11980 5108 12032 5117
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 11244 5040 11296 5092
rect 13452 5151 13504 5160
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 14188 5151 14240 5160
rect 13452 5108 13504 5117
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 13912 5040 13964 5092
rect 14648 5040 14700 5092
rect 12072 5015 12124 5024
rect 9864 4972 9916 4981
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 12164 4972 12216 5024
rect 13636 4972 13688 5024
rect 14188 4972 14240 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 14924 4972 14976 5024
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 1768 4768 1820 4820
rect 3148 4768 3200 4820
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 5264 4768 5316 4820
rect 5724 4811 5776 4820
rect 5724 4777 5733 4811
rect 5733 4777 5767 4811
rect 5767 4777 5776 4811
rect 5724 4768 5776 4777
rect 5908 4768 5960 4820
rect 6368 4768 6420 4820
rect 2136 4700 2188 4752
rect 4252 4700 4304 4752
rect 5448 4700 5500 4752
rect 6276 4700 6328 4752
rect 2688 4632 2740 4684
rect 3700 4632 3752 4684
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 4620 4632 4672 4684
rect 5080 4632 5132 4684
rect 5908 4632 5960 4684
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6460 4632 6512 4684
rect 7012 4632 7064 4684
rect 9956 4768 10008 4820
rect 10232 4768 10284 4820
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 13176 4811 13228 4820
rect 13176 4777 13185 4811
rect 13185 4777 13219 4811
rect 13219 4777 13228 4811
rect 13176 4768 13228 4777
rect 9404 4700 9456 4752
rect 10876 4700 10928 4752
rect 8208 4632 8260 4684
rect 9220 4632 9272 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 12624 4700 12676 4752
rect 13452 4632 13504 4684
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 4436 4564 4488 4616
rect 7748 4564 7800 4616
rect 11980 4564 12032 4616
rect 13360 4564 13412 4616
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 15108 4768 15160 4820
rect 14556 4564 14608 4573
rect 3792 4496 3844 4548
rect 4804 4496 4856 4548
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 3332 4471 3384 4480
rect 3332 4437 3341 4471
rect 3341 4437 3375 4471
rect 3375 4437 3384 4471
rect 4160 4471 4212 4480
rect 3332 4428 3384 4437
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 4344 4428 4396 4480
rect 4896 4428 4948 4480
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 5908 4428 5960 4480
rect 6460 4428 6512 4480
rect 7012 4496 7064 4548
rect 9588 4496 9640 4548
rect 11796 4496 11848 4548
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 8024 4428 8076 4480
rect 8300 4428 8352 4480
rect 9864 4471 9916 4480
rect 9864 4437 9873 4471
rect 9873 4437 9907 4471
rect 9907 4437 9916 4471
rect 9864 4428 9916 4437
rect 9956 4471 10008 4480
rect 9956 4437 9965 4471
rect 9965 4437 9999 4471
rect 9999 4437 10008 4471
rect 9956 4428 10008 4437
rect 11152 4428 11204 4480
rect 12164 4428 12216 4480
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 1860 4224 1912 4276
rect 2504 4224 2556 4276
rect 3332 4224 3384 4276
rect 3792 4224 3844 4276
rect 5080 4224 5132 4276
rect 5264 4224 5316 4276
rect 5632 4224 5684 4276
rect 7472 4224 7524 4276
rect 7748 4224 7800 4276
rect 8116 4224 8168 4276
rect 8300 4224 8352 4276
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 9864 4224 9916 4276
rect 11796 4224 11848 4276
rect 12716 4224 12768 4276
rect 13360 4224 13412 4276
rect 3976 4156 4028 4208
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3608 4088 3660 4140
rect 2688 4020 2740 4072
rect 3976 4020 4028 4072
rect 2228 3952 2280 4004
rect 4988 4088 5040 4140
rect 5540 4156 5592 4208
rect 6092 4156 6144 4208
rect 9772 4156 9824 4208
rect 13636 4156 13688 4208
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 3976 3884 4028 3936
rect 4528 4020 4580 4072
rect 5356 4020 5408 4072
rect 7196 4063 7248 4072
rect 7196 4029 7205 4063
rect 7205 4029 7239 4063
rect 7239 4029 7248 4063
rect 7196 4020 7248 4029
rect 7932 4020 7984 4072
rect 9680 4020 9732 4072
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 12164 4088 12216 4140
rect 12900 4088 12952 4140
rect 13084 4088 13136 4140
rect 10876 4020 10928 4029
rect 11796 4020 11848 4072
rect 8392 3952 8444 4004
rect 9220 3952 9272 4004
rect 10140 3952 10192 4004
rect 11060 3952 11112 4004
rect 11888 3952 11940 4004
rect 7104 3884 7156 3936
rect 11152 3884 11204 3936
rect 11980 3884 12032 3936
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 2320 3680 2372 3732
rect 1584 3544 1636 3596
rect 2872 3612 2924 3664
rect 3240 3680 3292 3732
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 4988 3680 5040 3732
rect 5172 3612 5224 3664
rect 5816 3680 5868 3732
rect 6460 3680 6512 3732
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 9956 3680 10008 3732
rect 10784 3680 10836 3732
rect 12532 3680 12584 3732
rect 7748 3655 7800 3664
rect 4620 3544 4672 3596
rect 5632 3544 5684 3596
rect 6276 3544 6328 3596
rect 3792 3476 3844 3528
rect 2320 3451 2372 3460
rect 2320 3417 2329 3451
rect 2329 3417 2363 3451
rect 2363 3417 2372 3451
rect 2320 3408 2372 3417
rect 2596 3340 2648 3392
rect 5080 3476 5132 3528
rect 6000 3476 6052 3528
rect 7748 3621 7757 3655
rect 7757 3621 7791 3655
rect 7791 3621 7800 3655
rect 7748 3612 7800 3621
rect 8300 3612 8352 3664
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 10876 3612 10928 3664
rect 10968 3612 11020 3664
rect 11520 3612 11572 3664
rect 11612 3612 11664 3664
rect 11704 3612 11756 3664
rect 12348 3612 12400 3664
rect 13912 3612 13964 3664
rect 7380 3544 7432 3553
rect 11152 3544 11204 3596
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 12624 3544 12676 3596
rect 14096 3544 14148 3596
rect 14648 3544 14700 3596
rect 7196 3519 7248 3528
rect 4528 3408 4580 3460
rect 4988 3408 5040 3460
rect 7196 3485 7205 3519
rect 7205 3485 7239 3519
rect 7239 3485 7248 3519
rect 7196 3476 7248 3485
rect 7472 3476 7524 3528
rect 7932 3476 7984 3528
rect 8116 3476 8168 3528
rect 11612 3476 11664 3528
rect 15292 3476 15344 3528
rect 5172 3340 5224 3392
rect 5632 3340 5684 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 8944 3408 8996 3460
rect 7564 3340 7616 3392
rect 9772 3408 9824 3460
rect 11060 3408 11112 3460
rect 12164 3408 12216 3460
rect 13544 3408 13596 3460
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 10140 3383 10192 3392
rect 9404 3340 9456 3349
rect 10140 3349 10149 3383
rect 10149 3349 10183 3383
rect 10183 3349 10192 3383
rect 10140 3340 10192 3349
rect 10232 3383 10284 3392
rect 10232 3349 10241 3383
rect 10241 3349 10275 3383
rect 10275 3349 10284 3383
rect 10232 3340 10284 3349
rect 10692 3340 10744 3392
rect 10876 3340 10928 3392
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 11980 3340 12032 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 13452 3383 13504 3392
rect 13452 3349 13461 3383
rect 13461 3349 13495 3383
rect 13495 3349 13504 3383
rect 13452 3340 13504 3349
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 1584 3136 1636 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 4804 3136 4856 3188
rect 5172 3136 5224 3188
rect 5540 3136 5592 3188
rect 5724 3136 5776 3188
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2228 3000 2280 3052
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2504 3000 2556 3052
rect 3148 3000 3200 3052
rect 4252 3068 4304 3120
rect 3516 3000 3568 3052
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4344 3000 4396 3052
rect 5448 3068 5500 3120
rect 4620 3000 4672 3052
rect 6460 3136 6512 3188
rect 6184 3068 6236 3120
rect 7564 3136 7616 3188
rect 7840 3136 7892 3188
rect 9128 3136 9180 3188
rect 9312 3136 9364 3188
rect 7472 3068 7524 3120
rect 9956 3068 10008 3120
rect 4528 2932 4580 2984
rect 6092 3000 6144 3052
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 7748 3000 7800 3052
rect 7932 3000 7984 3052
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9496 3000 9548 3052
rect 9772 3000 9824 3052
rect 10140 3136 10192 3188
rect 10968 3136 11020 3188
rect 11980 3136 12032 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13544 3179 13596 3188
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13912 3179 13964 3188
rect 13544 3136 13596 3145
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 11428 3068 11480 3120
rect 12072 3068 12124 3120
rect 13728 3068 13780 3120
rect 14832 3111 14884 3120
rect 14832 3077 14841 3111
rect 14841 3077 14875 3111
rect 14875 3077 14884 3111
rect 14832 3068 14884 3077
rect 10232 3000 10284 3052
rect 10968 3000 11020 3052
rect 11336 3043 11388 3052
rect 11336 3009 11345 3043
rect 11345 3009 11379 3043
rect 11379 3009 11388 3043
rect 11336 3000 11388 3009
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 14924 3000 14976 3052
rect 6368 2932 6420 2984
rect 7288 2932 7340 2984
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 8300 2932 8352 2984
rect 8852 2932 8904 2984
rect 1216 2864 1268 2916
rect 3240 2864 3292 2916
rect 5264 2864 5316 2916
rect 6000 2864 6052 2916
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 10048 2975 10100 2984
rect 9128 2932 9180 2941
rect 10048 2941 10057 2975
rect 10057 2941 10091 2975
rect 10091 2941 10100 2975
rect 10048 2932 10100 2941
rect 11520 2932 11572 2984
rect 1952 2796 2004 2848
rect 2320 2796 2372 2848
rect 3516 2839 3568 2848
rect 3516 2805 3525 2839
rect 3525 2805 3559 2839
rect 3559 2805 3568 2839
rect 3516 2796 3568 2805
rect 4160 2796 4212 2848
rect 5540 2796 5592 2848
rect 5908 2796 5960 2848
rect 6460 2796 6512 2848
rect 7840 2796 7892 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 9312 2864 9364 2916
rect 9404 2864 9456 2916
rect 10324 2864 10376 2916
rect 8576 2796 8628 2805
rect 11888 2864 11940 2916
rect 12440 2932 12492 2984
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 13084 2932 13136 2984
rect 13820 2932 13872 2984
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 15936 2932 15988 2984
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 2044 2592 2096 2644
rect 2412 2592 2464 2644
rect 3148 2592 3200 2644
rect 3792 2592 3844 2644
rect 3976 2592 4028 2644
rect 14924 2592 14976 2644
rect 3700 2524 3752 2576
rect 4620 2567 4672 2576
rect 4620 2533 4629 2567
rect 4629 2533 4663 2567
rect 4663 2533 4672 2567
rect 4620 2524 4672 2533
rect 4804 2567 4856 2576
rect 4804 2533 4813 2567
rect 4813 2533 4847 2567
rect 4847 2533 4856 2567
rect 4804 2524 4856 2533
rect 5540 2567 5592 2576
rect 5540 2533 5549 2567
rect 5549 2533 5583 2567
rect 5583 2533 5592 2567
rect 5540 2524 5592 2533
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 5172 2456 5224 2508
rect 6368 2524 6420 2576
rect 7564 2524 7616 2576
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 8116 2524 8168 2576
rect 10876 2567 10928 2576
rect 6276 2456 6328 2508
rect 3608 2388 3660 2440
rect 2504 2320 2556 2372
rect 5080 2320 5132 2372
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 6184 2431 6236 2440
rect 5356 2388 5408 2397
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 10048 2456 10100 2508
rect 10876 2533 10885 2567
rect 10885 2533 10919 2567
rect 10919 2533 10928 2567
rect 10876 2524 10928 2533
rect 11244 2524 11296 2576
rect 10968 2456 11020 2508
rect 11060 2456 11112 2508
rect 11336 2456 11388 2508
rect 12808 2456 12860 2508
rect 13360 2524 13412 2576
rect 13636 2567 13688 2576
rect 13636 2533 13645 2567
rect 13645 2533 13679 2567
rect 13679 2533 13688 2567
rect 13636 2524 13688 2533
rect 13820 2456 13872 2508
rect 8576 2320 8628 2372
rect 8852 2320 8904 2372
rect 10692 2320 10744 2372
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 4068 2252 4120 2304
rect 4528 2252 4580 2304
rect 7104 2252 7156 2304
rect 9312 2252 9364 2304
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 10324 2295 10376 2304
rect 9680 2252 9732 2261
rect 10324 2261 10333 2295
rect 10333 2261 10367 2295
rect 10367 2261 10376 2295
rect 10324 2252 10376 2261
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 11244 2320 11296 2372
rect 11612 2363 11664 2372
rect 11612 2329 11621 2363
rect 11621 2329 11655 2363
rect 11655 2329 11664 2363
rect 11612 2320 11664 2329
rect 12164 2320 12216 2372
rect 13084 2431 13136 2440
rect 13084 2397 13093 2431
rect 13093 2397 13127 2431
rect 13127 2397 13136 2431
rect 13084 2388 13136 2397
rect 13636 2388 13688 2440
rect 10416 2252 10468 2261
rect 10968 2252 11020 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 12348 2252 12400 2304
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 3792 2048 3844 2100
rect 5356 2048 5408 2100
rect 5448 2048 5500 2100
rect 10416 2048 10468 2100
rect 10692 2048 10744 2100
rect 12072 2048 12124 2100
rect 9220 1980 9272 2032
rect 11060 1980 11112 2032
rect 11612 1980 11664 2032
rect 12624 1980 12676 2032
rect 10508 1912 10560 1964
rect 11428 1912 11480 1964
rect 11888 1912 11940 1964
rect 9128 1844 9180 1896
rect 12716 1844 12768 1896
rect 5356 1776 5408 1828
rect 15016 1776 15068 1828
rect 10232 1436 10284 1488
rect 14464 1436 14516 1488
<< metal2 >>
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 2976 19230 3188 19258
rect 1044 17542 1072 19200
rect 1032 17536 1084 17542
rect 1032 17478 1084 17484
rect 1412 15434 1440 19200
rect 1674 19136 1730 19145
rect 1674 19071 1730 19080
rect 1688 16250 1716 19071
rect 1780 17898 1808 19200
rect 1780 17870 1900 17898
rect 1766 16688 1822 16697
rect 1766 16623 1822 16632
rect 1780 16590 1808 16623
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1872 16454 1900 17870
rect 2044 16584 2096 16590
rect 2042 16552 2044 16561
rect 2096 16552 2098 16561
rect 2042 16487 2098 16496
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15638 1624 15846
rect 2148 15706 2176 19200
rect 2318 17640 2374 17649
rect 2318 17575 2374 17584
rect 2332 16590 2360 17575
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2516 16250 2544 19200
rect 2884 19122 2912 19200
rect 2976 19122 3004 19230
rect 2884 19094 3004 19122
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2976 16590 3004 16730
rect 3160 16590 3188 19230
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 8864 19230 9076 19258
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3252 16522 3280 19200
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3240 16516 3292 16522
rect 3240 16458 3292 16464
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 3344 16182 3372 16526
rect 3620 16454 3648 19200
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3332 16176 3384 16182
rect 3252 16136 3332 16164
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11762 1532 12038
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 4321 1440 9454
rect 1596 9160 1624 15574
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 15366 2820 15438
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1674 14784 1730 14793
rect 1674 14719 1730 14728
rect 1688 14482 1716 14719
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1780 13841 1808 14894
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 3160 14482 3188 14758
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2412 13864 2464 13870
rect 1766 13832 1822 13841
rect 2412 13806 2464 13812
rect 1766 13767 1822 13776
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13326 2360 13670
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 12889 1716 13194
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12986 2360 13126
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 1674 12880 1730 12889
rect 2424 12866 2452 13806
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 1674 12815 1730 12824
rect 2332 12838 2452 12866
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1766 11928 1822 11937
rect 1766 11863 1822 11872
rect 1780 11830 1808 11863
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1964 11354 1992 12038
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1688 10130 1716 10911
rect 2056 10810 2084 12038
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 10810 2176 11494
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 2228 10056 2280 10062
rect 2226 10024 2228 10033
rect 2280 10024 2282 10033
rect 2226 9959 2282 9968
rect 2332 9874 2360 12838
rect 2516 11762 2544 13670
rect 2608 12646 2636 14350
rect 2700 13530 2728 14418
rect 3252 14362 3280 16136
rect 3332 16118 3384 16124
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3620 15910 3648 16050
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3330 15600 3386 15609
rect 3330 15535 3332 15544
rect 3384 15535 3386 15544
rect 3332 15506 3384 15512
rect 3160 14334 3280 14362
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2700 13394 2728 13466
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 3160 12968 3188 14334
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3252 13326 3280 14214
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3344 13841 3372 13874
rect 3330 13832 3386 13841
rect 3330 13767 3386 13776
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 2884 12940 3188 12968
rect 2884 12730 2912 12940
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2700 12702 2912 12730
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2700 12322 2728 12702
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 3160 12442 3188 12786
rect 3148 12436 3200 12442
rect 3252 12434 3280 13126
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3344 12782 3372 12854
rect 3436 12850 3464 15846
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3528 14074 3556 14962
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3620 13938 3648 15846
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 12986 3556 13330
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3344 12646 3372 12718
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3424 12436 3476 12442
rect 3252 12406 3372 12434
rect 3148 12378 3200 12384
rect 2700 12294 2820 12322
rect 2792 11898 2820 12294
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2792 11642 2820 11834
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2700 11614 2820 11642
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2516 10606 2544 11154
rect 2608 11014 2636 11494
rect 2700 11336 2728 11614
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 2700 11308 2820 11336
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2792 10452 2820 11308
rect 2746 10424 2820 10452
rect 2746 10146 2774 10424
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 3160 10266 3188 11698
rect 3344 11150 3372 12406
rect 3424 12378 3476 12384
rect 3332 11144 3384 11150
rect 3330 11112 3332 11121
rect 3384 11112 3386 11121
rect 3330 11047 3386 11056
rect 3436 10792 3464 12378
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11218 3556 11494
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3344 10764 3464 10792
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2746 10118 2820 10146
rect 2792 9926 2820 10118
rect 2240 9846 2360 9874
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9178 2084 9522
rect 1504 9132 1624 9160
rect 2044 9172 2096 9178
rect 1398 4312 1454 4321
rect 1398 4247 1454 4256
rect 1216 2916 1268 2922
rect 1216 2858 1268 2864
rect 1228 800 1256 2858
rect 1504 921 1532 9132
rect 2044 9114 2096 9120
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 1596 7478 1624 9007
rect 2148 8566 2176 9114
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 1674 8120 1730 8129
rect 1674 8055 1730 8064
rect 1688 7954 1716 8055
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1582 7168 1638 7177
rect 1582 7103 1638 7112
rect 1596 3602 1624 7103
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1688 5273 1716 6190
rect 1674 5264 1730 5273
rect 1674 5199 1730 5208
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4826 1808 5102
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1872 4282 1900 5170
rect 2148 4842 2176 8502
rect 2240 5778 2268 9846
rect 2332 9710 2544 9738
rect 2332 8634 2360 9710
rect 2516 9674 2544 9710
rect 2792 9674 2820 9862
rect 2412 9648 2464 9654
rect 2516 9646 2820 9674
rect 3160 9674 3188 10202
rect 3160 9646 3280 9674
rect 2412 9590 2464 9596
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2424 8362 2452 9590
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9042 2544 9318
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2608 8634 2636 9522
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2700 8378 2728 9386
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 3252 9178 3280 9646
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2516 8350 2728 8378
rect 2424 7954 2452 8298
rect 2516 8294 2544 8350
rect 2504 8288 2556 8294
rect 3068 8276 3096 8842
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8634 3188 8774
rect 3252 8634 3280 9114
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3344 8344 3372 10764
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 9926 3464 10610
rect 3528 10606 3556 11154
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10266 3556 10542
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 8566 3464 9862
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3252 8316 3372 8344
rect 3068 8248 3188 8276
rect 2504 8230 2556 8236
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 3160 8090 3188 8248
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7546 2452 7686
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2594 6216 2650 6225
rect 2594 6151 2650 6160
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2240 5352 2268 5714
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 5364 2372 5370
rect 2240 5324 2320 5352
rect 2320 5306 2372 5312
rect 2332 5114 2360 5306
rect 2424 5234 2452 5510
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2332 5086 2452 5114
rect 2148 4814 2268 4842
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 2148 4146 2176 4694
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2240 4010 2268 4814
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1490 912 1546 921
rect 1490 847 1546 856
rect 1596 800 1624 3130
rect 2240 3058 2268 3946
rect 2332 3738 2360 4422
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2332 3369 2360 3402
rect 2318 3360 2374 3369
rect 2318 3295 2374 3304
rect 2424 3058 2452 5086
rect 2516 4282 2544 6054
rect 2608 5302 2636 6151
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2700 4690 2728 6394
rect 2792 6322 2820 6598
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2976 5370 3004 5510
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 3160 4826 3188 6598
rect 3252 5302 3280 8316
rect 3330 8256 3386 8265
rect 3330 8191 3386 8200
rect 3344 7410 3372 8191
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3436 7342 3464 7890
rect 3528 7546 3556 8366
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5914 3464 6598
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3330 5264 3386 5273
rect 3330 5199 3332 5208
rect 3384 5199 3386 5208
rect 3332 5170 3384 5176
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2700 4078 2728 4626
rect 3238 4584 3294 4593
rect 3238 4519 3294 4528
rect 3146 4176 3202 4185
rect 3146 4111 3202 4120
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 2872 3664 2924 3670
rect 3160 3618 3188 4111
rect 3252 3738 3280 4519
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4282 3372 4422
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3344 3641 3372 4082
rect 2924 3612 3188 3618
rect 2872 3606 3188 3612
rect 2884 3590 3188 3606
rect 3330 3632 3386 3641
rect 3330 3567 3386 3576
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1964 800 1992 2790
rect 2056 2650 2084 2994
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2332 800 2360 2790
rect 2424 2650 2452 2994
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2516 2378 2544 2994
rect 2608 2774 2636 3334
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2608 2746 2728 2774
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 2700 800 2728 2746
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 3160 2650 3188 2994
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3252 1442 3280 2858
rect 3436 2774 3464 5510
rect 3528 3058 3556 6870
rect 3620 4146 3648 13738
rect 3712 12102 3740 16730
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16182 3832 16390
rect 3988 16250 4016 19200
rect 4066 18592 4122 18601
rect 4066 18527 4122 18536
rect 4080 18018 4108 18527
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3804 15473 3832 16118
rect 4080 15638 4108 17750
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4068 15632 4120 15638
rect 3988 15592 4068 15620
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3790 15464 3846 15473
rect 3790 15399 3846 15408
rect 3896 15366 3924 15506
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14482 3832 14894
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3804 13870 3832 14418
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13258 3832 13806
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3804 12918 3832 13194
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3896 12434 3924 15302
rect 3988 15162 4016 15592
rect 4068 15574 4120 15580
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4080 15162 4108 15370
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13870 4200 14214
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4264 13240 4292 17070
rect 4356 16454 4384 19200
rect 4724 17626 4752 19200
rect 4632 17598 4752 17626
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16590 4476 16934
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4448 15434 4476 16526
rect 4632 16182 4660 17598
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16794 4752 16934
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4724 16590 4752 16730
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 5092 16454 5120 19200
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 4620 16176 4672 16182
rect 5184 16130 5212 16730
rect 5276 16590 5304 16934
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 4620 16118 4672 16124
rect 5092 16102 5212 16130
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15502 4568 15846
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4436 15428 4488 15434
rect 4436 15370 4488 15376
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 15162 4660 15302
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 5092 15201 5120 16102
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 5078 15192 5134 15201
rect 4620 15156 4672 15162
rect 5078 15127 5134 15136
rect 4620 15098 4672 15104
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 4894 14920 4950 14929
rect 4894 14855 4950 14864
rect 4908 14618 4936 14855
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4908 14278 4936 14554
rect 5000 14278 5028 14758
rect 5092 14618 5120 14962
rect 5184 14958 5212 15982
rect 5276 15502 5304 16526
rect 5460 16153 5488 19200
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5446 16144 5502 16153
rect 5446 16079 5502 16088
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4988 14272 5040 14278
rect 5040 14232 5120 14260
rect 4988 14214 5040 14220
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 5092 13734 5120 14232
rect 5184 14074 5212 14894
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 4264 13212 4384 13240
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3988 12442 4016 12786
rect 3804 12406 3924 12434
rect 3976 12436 4028 12442
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3712 11558 3740 12038
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3804 10674 3832 12406
rect 3976 12378 4028 12384
rect 4172 12306 4200 12786
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3884 12232 3936 12238
rect 3882 12200 3884 12209
rect 3936 12200 3938 12209
rect 3882 12135 3938 12144
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11914 4016 12038
rect 3896 11898 4016 11914
rect 4172 11898 4200 12242
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 3884 11892 4016 11898
rect 3936 11886 4016 11892
rect 3884 11834 3936 11840
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3896 10062 3924 11630
rect 3988 11286 4016 11886
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4264 11830 4292 12106
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4356 11762 4384 13212
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 5092 12850 5120 13466
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4632 12238 4660 12786
rect 5276 12434 5304 14486
rect 5092 12406 5304 12434
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 5092 12084 5120 12406
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4632 12056 5120 12084
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4356 11286 4384 11698
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4344 11280 4396 11286
rect 4396 11240 4476 11268
rect 4344 11222 4396 11228
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3804 8294 3832 8502
rect 3896 8498 3924 9522
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3712 5778 3740 7482
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3712 4690 3740 5714
rect 3804 5352 3832 8230
rect 3896 8090 3924 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7818 4016 11222
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4080 9178 4108 10610
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4172 10062 4200 10542
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4356 9926 4384 10678
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 9178 4384 9862
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4080 8906 4108 9114
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4172 7818 4200 8978
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 3988 7410 4016 7754
rect 4252 7744 4304 7750
rect 4448 7732 4476 11240
rect 4304 7704 4476 7732
rect 4252 7686 4304 7692
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 6662 3924 7278
rect 3988 6934 4016 7346
rect 4172 6934 4200 7346
rect 4264 7274 4292 7686
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4264 6746 4292 7210
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4172 6718 4292 6746
rect 4344 6724 4396 6730
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6458 3924 6598
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3896 5778 3924 6258
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 4068 5704 4120 5710
rect 3974 5672 4030 5681
rect 4068 5646 4120 5652
rect 3974 5607 4030 5616
rect 3804 5324 3924 5352
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3804 4282 3832 4490
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 3738 3648 4082
rect 3792 3936 3844 3942
rect 3896 3924 3924 5324
rect 3988 4214 4016 5607
rect 4080 5574 4108 5646
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5166 4108 5510
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3976 4072 4028 4078
rect 4080 4060 4108 5102
rect 4172 4486 4200 6718
rect 4344 6666 4396 6672
rect 4356 6118 4384 6666
rect 4448 6322 4476 7142
rect 4436 6316 4488 6322
rect 4488 6276 4568 6304
rect 4436 6258 4488 6264
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 4758 4292 5170
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4028 4032 4108 4060
rect 3976 4014 4028 4020
rect 3976 3936 4028 3942
rect 3896 3896 3976 3924
rect 3792 3878 3844 3884
rect 3976 3878 4028 3884
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3344 2746 3464 2774
rect 3344 1465 3372 2746
rect 3068 1414 3280 1442
rect 3330 1456 3386 1465
rect 3068 800 3096 1414
rect 3330 1391 3386 1400
rect 3528 1034 3556 2790
rect 3620 2446 3648 3674
rect 3804 3534 3832 3878
rect 3988 3738 4016 3878
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4172 3097 4200 4422
rect 4264 3126 4292 4694
rect 4356 4690 4384 6054
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4252 3120 4304 3126
rect 4158 3088 4214 3097
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3792 3052 3844 3058
rect 4252 3062 4304 3068
rect 4356 3058 4384 4422
rect 4448 3738 4476 4558
rect 4540 4078 4568 6276
rect 4632 5681 4660 12056
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 5184 11830 5212 12310
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 4618 5672 4674 5681
rect 4618 5607 4674 5616
rect 4698 5468 5006 5477
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4540 3584 4568 4014
rect 4632 3602 4660 4626
rect 4816 4554 4844 5238
rect 5092 5166 5120 11494
rect 5184 10810 5212 11766
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 5370 5212 7822
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4908 4486 4936 4762
rect 5092 4690 5120 5102
rect 5276 4826 5304 11494
rect 5368 8294 5396 15370
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15094 5488 15302
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5460 14396 5488 15030
rect 5552 14550 5580 17138
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16658 5764 16934
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5736 16266 5764 16594
rect 5828 16454 5856 19200
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 6012 16998 6040 17818
rect 6196 17678 6224 19200
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6564 17270 6592 19200
rect 6932 17338 6960 19200
rect 7300 17338 7328 19200
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 7668 17066 7696 19200
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 6012 16590 6040 16934
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5736 16238 5856 16266
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15570 5764 16050
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5644 15366 5672 15506
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5644 15162 5672 15302
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5644 14550 5672 15098
rect 5828 15094 5856 16238
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5736 14618 5764 14894
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5632 14544 5684 14550
rect 5632 14486 5684 14492
rect 5540 14408 5592 14414
rect 5460 14368 5540 14396
rect 5540 14350 5592 14356
rect 5828 14346 5856 15030
rect 5920 14958 5948 15982
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5920 14482 5948 14894
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5816 14340 5868 14346
rect 5816 14282 5868 14288
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5552 13530 5580 13874
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5552 13326 5580 13466
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12918 5580 13262
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5460 10742 5488 12310
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5552 11558 5580 11766
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5644 10742 5672 14214
rect 5920 14006 5948 14418
rect 5908 14000 5960 14006
rect 6196 13977 6224 15642
rect 6288 15434 6316 16662
rect 7012 16652 7064 16658
rect 7064 16612 7144 16640
rect 7012 16594 7064 16600
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15706 6408 16390
rect 6828 16040 6880 16046
rect 6880 15988 6960 15994
rect 6828 15982 6960 15988
rect 6840 15966 6960 15982
rect 6932 15910 6960 15966
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6380 15502 6408 15533
rect 6368 15496 6420 15502
rect 6420 15444 6960 15450
rect 6368 15438 6960 15444
rect 6380 15434 6960 15438
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6380 15428 6972 15434
rect 6380 15422 6920 15428
rect 5908 13942 5960 13948
rect 6182 13968 6238 13977
rect 5920 13462 5948 13942
rect 6182 13903 6238 13912
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13530 6132 13806
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10742 5856 11290
rect 6288 11082 6316 15370
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5644 9674 5672 10678
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10062 5764 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5736 9722 5764 9998
rect 5460 9646 5672 9674
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5460 7834 5488 9646
rect 5736 9042 5764 9658
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8634 5580 8842
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5368 7806 5488 7834
rect 5368 5760 5396 7806
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7410 5488 7686
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5368 5732 5580 5760
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 5092 4282 5120 4422
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 3738 5028 4082
rect 5276 4060 5304 4218
rect 5368 4078 5396 5578
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5184 4032 5304 4060
rect 5356 4072 5408 4078
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5184 3670 5212 4032
rect 5460 4049 5488 4694
rect 5552 4298 5580 5732
rect 5644 5166 5672 8774
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5828 5914 5856 7142
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5736 4826 5764 5646
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5552 4282 5672 4298
rect 5552 4276 5684 4282
rect 5552 4270 5632 4276
rect 5632 4218 5684 4224
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5356 4014 5408 4020
rect 5446 4040 5502 4049
rect 5446 3975 5502 3984
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 4448 3556 4568 3584
rect 4620 3596 4672 3602
rect 4158 3023 4214 3032
rect 4344 3052 4396 3058
rect 3792 2994 3844 3000
rect 4344 2994 4396 3000
rect 3712 2582 3740 2994
rect 3804 2650 3832 2994
rect 4448 2972 4476 3556
rect 4620 3538 4672 3544
rect 5080 3528 5132 3534
rect 4986 3496 5042 3505
rect 4528 3460 4580 3466
rect 5080 3470 5132 3476
rect 4986 3431 4988 3440
rect 4528 3402 4580 3408
rect 5040 3431 5042 3440
rect 4988 3402 5040 3408
rect 4540 3194 4568 3402
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4528 2984 4580 2990
rect 4448 2944 4528 2972
rect 4528 2926 4580 2932
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3974 2680 4030 2689
rect 3792 2644 3844 2650
rect 3974 2615 3976 2624
rect 3792 2586 3844 2592
rect 4028 2615 4030 2624
rect 3976 2586 4028 2592
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3804 2106 3832 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3436 1006 3556 1034
rect 3436 800 3464 1006
rect 3804 870 3924 898
rect 3804 800 3832 870
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 3896 762 3924 870
rect 4080 762 4108 2246
rect 4172 800 4200 2790
rect 4632 2582 4660 2994
rect 4816 2582 4844 3130
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 5092 2378 5120 3470
rect 5184 3398 5212 3429
rect 5172 3392 5224 3398
rect 5170 3360 5172 3369
rect 5224 3360 5226 3369
rect 5170 3295 5226 3304
rect 5184 3194 5212 3295
rect 5552 3194 5580 4150
rect 5644 3602 5672 4218
rect 5828 3738 5856 5170
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5920 4486 5948 4626
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5920 3618 5948 4422
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5828 3590 5948 3618
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 800 4568 2246
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 4908 870 5028 898
rect 4908 800 4936 870
rect 3896 734 4108 762
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5000 762 5028 870
rect 5184 762 5212 2450
rect 5276 800 5304 2858
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5368 2106 5396 2382
rect 5460 2106 5488 3062
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2582 5580 2790
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 5368 1834 5396 2042
rect 5356 1828 5408 1834
rect 5356 1770 5408 1776
rect 5644 800 5672 3334
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2564 5764 3130
rect 5828 3097 5856 3590
rect 6012 3534 6040 8910
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6104 4978 6132 6394
rect 6196 5098 6224 6394
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6104 4950 6224 4978
rect 6090 4720 6146 4729
rect 6090 4655 6092 4664
rect 6144 4655 6146 4664
rect 6092 4626 6144 4632
rect 6104 4214 6132 4626
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 6000 3528 6052 3534
rect 5906 3496 5962 3505
rect 6000 3470 6052 3476
rect 5906 3431 5962 3440
rect 5814 3088 5870 3097
rect 5814 3023 5870 3032
rect 5920 2854 5948 3431
rect 6104 3058 6132 4150
rect 6196 3482 6224 4950
rect 6288 4758 6316 5850
rect 6380 4826 6408 15422
rect 6920 15370 6972 15376
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15162 6868 15302
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 13258 6500 14418
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14006 6776 14214
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6472 12442 6500 13194
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 7116 11354 7144 16612
rect 7576 16590 7604 16934
rect 7760 16794 7788 17206
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7944 16794 7972 16934
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7944 16454 7972 16730
rect 8036 16522 8064 19200
rect 8404 17542 8432 19200
rect 8772 19122 8800 19200
rect 8864 19122 8892 19230
rect 8772 19094 8892 19122
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16658 8248 17070
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7392 15910 7420 16050
rect 7484 15910 7512 16186
rect 7944 16114 7972 16390
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 7656 16040 7708 16046
rect 8116 16040 8168 16046
rect 7656 15982 7708 15988
rect 8114 16008 8116 16017
rect 8168 16008 8170 16017
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7208 12434 7236 15846
rect 7484 15609 7512 15846
rect 7470 15600 7526 15609
rect 7470 15535 7526 15544
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14618 7328 14962
rect 7576 14958 7604 15506
rect 7668 15366 7696 15982
rect 8114 15943 8170 15952
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13530 7420 13738
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7392 12986 7420 13466
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7208 12406 7420 12434
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 7300 11558 7328 12174
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7546 6960 7890
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7546 7052 7686
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7024 7206 7052 7346
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6322 6500 6598
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6472 5710 6500 6258
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6734 5808 6790 5817
rect 6734 5743 6790 5752
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5370 6500 5646
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6748 5166 6776 5743
rect 7116 5710 7144 8298
rect 7208 8090 7236 8502
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7300 7886 7328 8774
rect 7392 8616 7420 12406
rect 7576 10674 7604 14894
rect 7668 12434 7696 15302
rect 7760 14074 7788 15642
rect 7852 15434 7880 15846
rect 8220 15570 8248 16594
rect 8588 16590 8616 17138
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8404 15910 8432 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8404 15502 8432 15846
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 8036 14958 8064 15438
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15178 8340 15302
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8220 15150 8340 15178
rect 8864 15162 8892 15982
rect 8956 15706 8984 16050
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8852 15156 8904 15162
rect 8220 15094 8248 15150
rect 8852 15098 8904 15104
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7852 14618 7880 14758
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 14414 7880 14554
rect 8036 14482 8064 14894
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 8116 14408 8168 14414
rect 8220 14396 8248 15030
rect 8168 14368 8248 14396
rect 8404 14362 8432 15030
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8864 14822 8892 14894
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8116 14350 8168 14356
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7760 13258 7788 14010
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 8128 12434 8156 14350
rect 8312 14334 8432 14362
rect 8312 14074 8340 14334
rect 8864 14278 8892 14758
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8496 13190 8524 14010
rect 8864 13870 8892 14214
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13394 8892 13806
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 7668 12406 7788 12434
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 9382 7604 10610
rect 7668 9994 7696 11290
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7392 8588 7604 8616
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5364 6972 5370
rect 7024 5352 7052 5510
rect 6972 5324 7052 5352
rect 6920 5306 6972 5312
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6288 3602 6316 4694
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6196 3454 6316 3482
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5816 2576 5868 2582
rect 5736 2544 5816 2564
rect 5868 2544 5870 2553
rect 5736 2536 5814 2544
rect 5814 2479 5870 2488
rect 6012 800 6040 2858
rect 6196 2446 6224 3062
rect 6288 2514 6316 3454
rect 6380 2990 6408 4762
rect 6472 4690 6500 4966
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 7024 4690 7052 5324
rect 7116 5166 7144 5646
rect 7300 5642 7328 7822
rect 7484 6662 7512 8434
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7288 5636 7340 5642
rect 7288 5578 7340 5584
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7208 5098 7236 5510
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 3738 6500 4422
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6460 3392 6512 3398
rect 7024 3369 7052 4490
rect 7208 4162 7236 5034
rect 7116 4134 7236 4162
rect 7116 3942 7144 4134
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7208 3534 7236 4014
rect 7392 3602 7420 5102
rect 7484 4282 7512 5170
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 3596 7432 3602
rect 7300 3556 7380 3584
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6460 3334 6512 3340
rect 7010 3360 7066 3369
rect 6472 3194 6500 3334
rect 7010 3295 7066 3304
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6368 2984 6420 2990
rect 6748 2961 6776 2994
rect 7300 2990 7328 3556
rect 7380 3538 7432 3544
rect 7484 3534 7512 4218
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7576 3398 7604 8588
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 3194 7604 3334
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7288 2984 7340 2990
rect 6368 2926 6420 2932
rect 6734 2952 6790 2961
rect 7288 2926 7340 2932
rect 6734 2887 6790 2896
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6380 800 6408 2518
rect 5000 734 5212 762
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6472 762 6500 2790
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 6656 870 6776 898
rect 6656 762 6684 870
rect 6748 800 6776 870
rect 7116 800 7144 2246
rect 7484 800 7512 3062
rect 7562 2816 7618 2825
rect 7562 2751 7618 2760
rect 7576 2582 7604 2751
rect 7564 2576 7616 2582
rect 7668 2553 7696 5646
rect 7760 4622 7788 12406
rect 8036 12406 8156 12434
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11082 7880 11494
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7852 10674 7880 11018
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7852 5817 7880 7142
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7838 5808 7894 5817
rect 7838 5743 7894 5752
rect 7944 5574 7972 6258
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7760 4282 7788 4422
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7746 3768 7802 3777
rect 7746 3703 7802 3712
rect 7760 3670 7788 3703
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7760 3058 7788 3606
rect 7852 3194 7880 5238
rect 7944 4078 7972 5510
rect 8036 4740 8064 12406
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8128 12102 8156 12310
rect 8772 12238 8800 12854
rect 8956 12714 8984 15438
rect 9048 15162 9076 19230
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11702 19200 11758 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14384 19230 14596 19258
rect 9140 15722 9168 19200
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 16590 9260 16934
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9232 16289 9260 16526
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9218 16280 9274 16289
rect 9218 16215 9274 16224
rect 9232 15978 9260 16215
rect 9324 16182 9352 16390
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9416 16046 9444 16594
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9140 15694 9260 15722
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9140 14550 9168 15438
rect 9232 15434 9260 15694
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9586 8156 9998
rect 8312 9722 8340 12038
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 8956 11082 8984 12650
rect 9048 12102 9076 14418
rect 9140 14074 9168 14486
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9140 12442 9168 13330
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9232 11898 9260 15370
rect 9324 14958 9352 15506
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 12850 9352 14894
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9048 11286 9076 11766
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 9048 10810 9076 11222
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8758 10568 8814 10577
rect 8758 10503 8814 10512
rect 8772 10266 8800 10503
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8128 9178 8156 9522
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8220 7206 8248 9522
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8956 8498 8984 9114
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8090 8984 8434
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 5098 8156 6598
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8864 6390 8892 6802
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8036 4712 8156 4740
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7760 2582 7788 2994
rect 7852 2990 7880 3130
rect 7944 3058 7972 3470
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7748 2576 7800 2582
rect 7564 2518 7616 2524
rect 7654 2544 7710 2553
rect 7748 2518 7800 2524
rect 7654 2479 7710 2488
rect 7852 800 7880 2790
rect 8036 2582 8064 4422
rect 8128 4282 8156 4712
rect 8220 4690 8248 6054
rect 8864 5914 8892 6326
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 6118 8984 6258
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8312 5778 8340 5850
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5234 8340 5714
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8128 3534 8156 4218
rect 8220 4162 8248 4626
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4282 8340 4422
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8220 4134 8340 4162
rect 8206 3768 8262 3777
rect 8206 3703 8262 3712
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8220 3233 8248 3703
rect 8312 3670 8340 4134
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 8404 3380 8432 3946
rect 8850 3632 8906 3641
rect 8850 3567 8906 3576
rect 8312 3352 8432 3380
rect 8864 3369 8892 3567
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 8850 3360 8906 3369
rect 8206 3224 8262 3233
rect 8206 3159 8262 3168
rect 8206 3088 8262 3097
rect 8116 3052 8168 3058
rect 8206 3023 8262 3032
rect 8116 2994 8168 3000
rect 8128 2582 8156 2994
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8220 800 8248 3023
rect 8312 2990 8340 3352
rect 8446 3292 8754 3301
rect 8850 3295 8906 3304
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8956 3058 8984 3402
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8496 2514 8524 2790
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8588 2378 8616 2790
rect 8864 2378 8892 2926
rect 9048 2774 9076 10202
rect 9220 8492 9272 8498
rect 9140 8452 9220 8480
rect 9140 6458 9168 8452
rect 9220 8434 9272 8440
rect 9324 7528 9352 12378
rect 9416 11354 9444 15982
rect 9508 15366 9536 19200
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9784 17134 9812 17274
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9600 16590 9628 16934
rect 9784 16726 9812 17070
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9588 16584 9640 16590
rect 9586 16552 9588 16561
rect 9640 16552 9642 16561
rect 9784 16522 9812 16662
rect 9586 16487 9642 16496
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 14618 9536 15302
rect 9692 15162 9720 16390
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9508 14074 9536 14554
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9600 13938 9628 14214
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9784 12646 9812 16458
rect 9876 15994 9904 19200
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9968 16590 9996 16934
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10244 16130 10272 19200
rect 10612 16980 10640 19200
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17270 10916 17546
rect 10876 17264 10928 17270
rect 10874 17232 10876 17241
rect 10928 17232 10930 17241
rect 10784 17196 10836 17202
rect 10874 17167 10930 17176
rect 10784 17138 10836 17144
rect 10612 16952 10732 16980
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10152 16102 10272 16130
rect 10152 16017 10180 16102
rect 10232 16040 10284 16046
rect 10138 16008 10194 16017
rect 9876 15966 10088 15994
rect 9876 14278 9904 15966
rect 10060 15910 10088 15966
rect 10232 15982 10284 15988
rect 10138 15943 10194 15952
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9968 15162 9996 15846
rect 10244 15706 10272 15982
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10704 15638 10732 16952
rect 10796 16250 10824 17138
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16590 10916 17070
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10888 16046 10916 16526
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10980 15706 11008 19200
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11164 16590 11192 16730
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 16153 11192 16186
rect 11150 16144 11206 16153
rect 11256 16114 11284 17818
rect 11150 16079 11206 16088
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10980 15502 11008 15642
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10600 15360 10652 15366
rect 10598 15328 10600 15337
rect 10652 15328 10654 15337
rect 10598 15263 10654 15272
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9996 13954
rect 9876 13932 10008 13938
rect 9876 13926 9956 13932
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9876 11762 9904 13926
rect 9956 13874 10008 13880
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9416 11150 9444 11290
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9968 11082 9996 13738
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9968 10810 9996 11018
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10060 10742 10088 13738
rect 10152 13258 10180 14894
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13530 10272 13670
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 11354 10180 13194
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9722 9628 9930
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 7818 9628 9318
rect 10060 9110 10088 10678
rect 10152 10266 10180 10678
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10152 9654 10180 10202
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 9178 10180 9590
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9232 7500 9352 7528
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9140 3890 9168 5578
rect 9232 5234 9260 7500
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 7290 9352 7346
rect 9324 7262 9444 7290
rect 9600 7274 9628 7754
rect 9876 7546 9904 7822
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9416 6798 9444 7262
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9876 7002 9904 7482
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9968 6866 9996 7142
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 4690 9260 5170
rect 9416 5098 9444 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5642 9720 6054
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9232 4010 9260 4626
rect 9416 4282 9444 4694
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9600 3890 9628 4490
rect 9692 4078 9720 5578
rect 9784 4690 9812 6598
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 9876 5370 9904 5510
rect 9864 5364 9916 5370
rect 9916 5324 10088 5352
rect 9864 5306 9916 5312
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9876 4593 9904 4966
rect 9954 4856 10010 4865
rect 9954 4791 9956 4800
rect 10008 4791 10010 4800
rect 9956 4762 10008 4768
rect 9862 4584 9918 4593
rect 9862 4519 9918 4528
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9876 4282 9904 4422
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9140 3862 9260 3890
rect 9600 3862 9720 3890
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9140 2990 9168 3130
rect 9232 3074 9260 3862
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9324 3194 9352 3334
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9232 3046 9352 3074
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9218 2952 9274 2961
rect 9324 2922 9352 3046
rect 9416 2922 9444 3334
rect 9692 3210 9720 3862
rect 9784 3738 9812 4150
rect 9968 3738 9996 4422
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9600 3182 9720 3210
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9218 2887 9274 2896
rect 9312 2916 9364 2922
rect 9048 2746 9168 2774
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8588 870 8708 898
rect 8588 800 8616 870
rect 6472 734 6684 762
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8680 762 8708 870
rect 8864 762 8892 2314
rect 9140 1902 9168 2746
rect 9232 2038 9260 2887
rect 9312 2858 9364 2864
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 9324 2310 9352 2858
rect 9508 2774 9536 2994
rect 9600 2836 9628 3182
rect 9784 3058 9812 3402
rect 9956 3120 10008 3126
rect 9954 3088 9956 3097
rect 10008 3088 10010 3097
rect 9772 3052 9824 3058
rect 9954 3023 10010 3032
rect 9772 2994 9824 3000
rect 10060 2990 10088 5324
rect 10152 4010 10180 5510
rect 10244 5370 10272 12582
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10704 12442 10732 15438
rect 11256 15366 11284 16050
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11348 15162 11376 19200
rect 11716 17082 11744 19200
rect 11624 17054 11744 17082
rect 11796 17060 11848 17066
rect 11518 16416 11574 16425
rect 11518 16351 11574 16360
rect 11532 16250 11560 16351
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11152 15088 11204 15094
rect 10874 15056 10930 15065
rect 11152 15030 11204 15036
rect 10874 14991 10930 15000
rect 10888 14618 10916 14991
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10888 14006 10916 14554
rect 11072 14090 11100 14758
rect 10980 14062 11100 14090
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10980 13841 11008 14062
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10966 13832 11022 13841
rect 11072 13818 11100 13942
rect 11164 13938 11192 15030
rect 11348 14929 11376 15098
rect 11334 14920 11390 14929
rect 11334 14855 11390 14864
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11072 13790 11192 13818
rect 10966 13767 11022 13776
rect 10980 13716 11008 13767
rect 10980 13688 11100 13716
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11762 10916 12174
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10888 11354 10916 11698
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10810 10548 11154
rect 10980 11082 11008 11562
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10704 8634 10732 9114
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11072 8294 11100 13688
rect 11164 10282 11192 13790
rect 11256 10810 11284 14010
rect 11348 13870 11376 14350
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11348 13394 11376 13806
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11348 12918 11376 13330
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12374 11376 12854
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11440 12170 11468 15982
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11164 10254 11284 10282
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9722 11192 10066
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10888 6662 10916 6802
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4826 10272 5034
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10704 3398 10732 5306
rect 10888 4758 10916 6598
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10888 4078 10916 4694
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10796 3738 10824 4014
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10888 3670 10916 4014
rect 10980 3670 11008 8230
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 5846 11100 7346
rect 11256 6882 11284 10254
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11334 9072 11390 9081
rect 11334 9007 11390 9016
rect 11348 8974 11376 9007
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11348 7410 11376 7822
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11164 6854 11284 6882
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 4010 11100 5782
rect 11164 4570 11192 6854
rect 11348 6798 11376 7346
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 5914 11284 6666
rect 11348 6458 11376 6734
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 6202 11468 10202
rect 11348 6174 11468 6202
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11256 5098 11284 5850
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11164 4542 11284 4570
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4049 11192 4422
rect 11150 4040 11206 4049
rect 11060 4004 11112 4010
rect 11150 3975 11206 3984
rect 11060 3946 11112 3952
rect 11164 3942 11192 3975
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10980 3482 11008 3606
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 10796 3454 11008 3482
rect 11060 3460 11112 3466
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10152 3194 10180 3334
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 3058 10272 3334
rect 10322 3088 10378 3097
rect 10232 3052 10284 3058
rect 10796 3040 10824 3454
rect 11060 3402 11112 3408
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10322 3023 10378 3032
rect 10232 2994 10284 3000
rect 10048 2984 10100 2990
rect 10100 2944 10180 2972
rect 10048 2926 10100 2932
rect 9600 2808 9904 2836
rect 9508 2746 9674 2774
rect 9646 2496 9674 2746
rect 9646 2468 9720 2496
rect 9692 2310 9720 2468
rect 9876 2417 9904 2808
rect 10152 2774 10180 2944
rect 10060 2746 10180 2774
rect 10060 2514 10088 2746
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9862 2408 9918 2417
rect 9862 2343 9918 2352
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 8956 870 9076 898
rect 8956 800 8984 870
rect 8680 734 8892 762
rect 8942 0 8998 800
rect 9048 762 9076 870
rect 9232 762 9260 1974
rect 9324 800 9352 2246
rect 9876 2122 9904 2343
rect 10046 2272 10102 2281
rect 10046 2207 10102 2216
rect 9692 2094 9904 2122
rect 9692 800 9720 2094
rect 10060 800 10088 2207
rect 10244 1494 10272 2994
rect 10336 2922 10364 3023
rect 10520 3012 10824 3040
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10520 2836 10548 3012
rect 10612 2961 10824 2972
rect 10598 2952 10824 2961
rect 10654 2944 10824 2952
rect 10598 2887 10654 2896
rect 10520 2808 10732 2836
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10704 2378 10732 2808
rect 10692 2372 10744 2378
rect 10692 2314 10744 2320
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10336 1986 10364 2246
rect 10428 2122 10456 2246
rect 10428 2106 10548 2122
rect 10704 2106 10732 2314
rect 10416 2100 10548 2106
rect 10468 2094 10548 2100
rect 10416 2042 10468 2048
rect 10336 1958 10456 1986
rect 10520 1970 10548 2094
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10232 1488 10284 1494
rect 10232 1430 10284 1436
rect 10428 800 10456 1958
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 10796 800 10824 2944
rect 10888 2582 10916 3334
rect 10980 3194 11008 3334
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10966 3088 11022 3097
rect 10966 3023 10968 3032
rect 11020 3023 11022 3032
rect 10968 2994 11020 3000
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10980 2514 11008 2994
rect 11072 2514 11100 3402
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10980 2310 11008 2450
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11072 2038 11100 2450
rect 11060 2032 11112 2038
rect 11060 1974 11112 1980
rect 11164 800 11192 3538
rect 11256 3505 11284 4542
rect 11242 3496 11298 3505
rect 11242 3431 11298 3440
rect 11256 2825 11284 3431
rect 11348 3058 11376 6174
rect 11532 6066 11560 15574
rect 11624 15094 11652 17054
rect 11796 17002 11848 17008
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11716 16726 11744 16934
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11808 16658 11836 17002
rect 11980 16992 12032 16998
rect 11900 16952 11980 16980
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 15706 11744 16390
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11624 13530 11652 14894
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 12918 11652 13466
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11808 12730 11836 16594
rect 11900 16114 11928 16952
rect 11980 16934 12032 16940
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 16250 12020 16390
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 12084 15881 12112 19200
rect 12452 17626 12480 19200
rect 12452 17598 12572 17626
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12544 17218 12572 17598
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12452 17190 12572 17218
rect 12452 16590 12480 17190
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12544 16794 12572 17070
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12636 16726 12664 16934
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12544 16182 12572 16594
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12440 15904 12492 15910
rect 12070 15872 12126 15881
rect 12440 15846 12492 15852
rect 12070 15807 12126 15816
rect 12452 15502 12480 15846
rect 12544 15570 12572 16118
rect 12636 16114 12664 16526
rect 12728 16250 12756 17274
rect 12820 17270 12848 19200
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12820 15978 12848 16458
rect 12912 15978 12940 17682
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17338 13032 17478
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13188 16998 13216 19200
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17338 13400 17614
rect 13556 17354 13584 19200
rect 13360 17332 13412 17338
rect 13556 17326 13768 17354
rect 13360 17274 13412 17280
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12912 15706 12940 15914
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11624 12702 11836 12730
rect 11624 12442 11652 12702
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 11694 11652 12378
rect 11808 12102 11836 12582
rect 11900 12102 11928 15302
rect 12084 15162 12112 15370
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11992 12442 12020 14010
rect 12084 13530 12112 14214
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12084 12628 12112 13466
rect 12544 13190 12572 15506
rect 12820 15366 12848 15574
rect 13096 15570 13124 16050
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13188 15450 13216 16934
rect 13464 16658 13492 17206
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13372 15994 13400 16050
rect 13096 15422 13216 15450
rect 13280 15966 13400 15994
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12636 15162 12664 15302
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12820 15026 12848 15302
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12164 12640 12216 12646
rect 12084 12600 12164 12628
rect 12164 12582 12216 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12544 12170 12572 13126
rect 12820 12714 12848 13942
rect 12912 13258 12940 14894
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 14074 13032 14282
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 13096 12434 13124 15422
rect 13280 15366 13308 15966
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15065 13308 15302
rect 13266 15056 13322 15065
rect 13266 14991 13322 15000
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14822 13308 14894
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13188 13530 13216 14350
rect 13280 14006 13308 14758
rect 13372 14278 13400 14962
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13372 13530 13400 14214
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12986 13308 13126
rect 13372 12986 13400 13194
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13096 12406 13216 12434
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11014 12112 11630
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11900 10606 11928 10950
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 12084 9994 12112 10950
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12544 10470 12572 11698
rect 12636 11150 12664 12174
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10810 12664 11086
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12728 10470 12756 11766
rect 12820 10742 12848 12038
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12714 10024 12770 10033
rect 12072 9988 12124 9994
rect 12714 9959 12770 9968
rect 12072 9930 12124 9936
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11624 8974 11652 9862
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 12728 8906 12756 9959
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9110 12848 9522
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11440 6038 11560 6066
rect 11440 3126 11468 6038
rect 11624 5273 11652 8230
rect 11808 7478 11836 8298
rect 12084 8090 12112 8842
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 12728 8634 12756 8842
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12820 8401 12848 8774
rect 12806 8392 12862 8401
rect 12806 8327 12808 8336
rect 12860 8327 12862 8336
rect 12808 8298 12860 8304
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 12084 7410 12112 8026
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7818 12664 7958
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11808 5710 11836 6394
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 5370 11836 5646
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11610 5264 11666 5273
rect 11520 5228 11572 5234
rect 11610 5199 11666 5208
rect 11520 5170 11572 5176
rect 11532 4826 11560 5170
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11624 3670 11652 5199
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 4282 11836 4490
rect 11900 4468 11928 6598
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12544 5642 12572 6598
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12544 5250 12572 5578
rect 12544 5222 12664 5250
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 11992 4622 12020 5102
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11900 4440 12020 4468
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11242 2816 11298 2825
rect 11242 2751 11298 2760
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 11256 2378 11284 2518
rect 11348 2514 11376 2994
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11440 1970 11468 3062
rect 11532 2990 11560 3606
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11532 800 11560 2751
rect 11624 2378 11652 3470
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11624 2038 11652 2314
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11716 1034 11744 3606
rect 11808 1442 11836 4014
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 3602 11928 3946
rect 11992 3942 12020 4440
rect 12084 4185 12112 4966
rect 12176 4486 12204 4966
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12070 4176 12126 4185
rect 12070 4111 12126 4120
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12070 4040 12126 4049
rect 12070 3975 12126 3984
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 2922 11928 3538
rect 11992 3398 12020 3878
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3194 12020 3334
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12084 3126 12112 3975
rect 12176 3466 12204 4082
rect 12346 3768 12402 3777
rect 12544 3738 12572 5102
rect 12636 4758 12664 5222
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12346 3703 12402 3712
rect 12532 3732 12584 3738
rect 12360 3670 12388 3703
rect 12532 3674 12584 3680
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12636 3602 12664 4694
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12346 3088 12402 3097
rect 12346 3023 12402 3032
rect 12624 3052 12676 3058
rect 12360 2938 12388 3023
rect 12728 3040 12756 4218
rect 12676 3012 12756 3040
rect 12624 2994 12676 3000
rect 12820 2990 12848 7414
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 6730 12940 7210
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 4146 12940 6054
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12440 2984 12492 2990
rect 12360 2932 12440 2938
rect 12360 2926 12492 2932
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 11888 2916 11940 2922
rect 12360 2910 12480 2926
rect 11888 2858 11940 2864
rect 12820 2514 12848 2926
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12176 2378 12388 2394
rect 12164 2372 12388 2378
rect 12216 2366 12388 2372
rect 12164 2314 12216 2320
rect 12360 2310 12388 2366
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 11900 1970 11928 2246
rect 12084 2106 12112 2246
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12714 2136 12770 2145
rect 12072 2100 12124 2106
rect 12714 2071 12770 2080
rect 12072 2042 12124 2048
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11808 1414 12020 1442
rect 11716 1006 11928 1034
rect 11900 800 11928 1006
rect 9048 734 9260 762
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 11992 762 12020 1414
rect 12176 870 12296 898
rect 12176 762 12204 870
rect 12268 800 12296 870
rect 12636 800 12664 1974
rect 12728 1902 12756 2071
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 13004 800 13032 12038
rect 13188 11694 13216 12406
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13188 11558 13216 11630
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9081 13216 11494
rect 13372 10810 13400 11494
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13174 9072 13230 9081
rect 13174 9007 13230 9016
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7002 13124 7754
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 6254 13124 6938
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 4706 13124 5510
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13188 4826 13216 5170
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13096 4678 13216 4706
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 2990 13124 4082
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13188 2836 13216 4678
rect 13096 2808 13216 2836
rect 13096 2446 13124 2808
rect 13084 2440 13136 2446
rect 13082 2408 13084 2417
rect 13136 2408 13138 2417
rect 13280 2394 13308 8502
rect 13372 4622 13400 10406
rect 13464 7426 13492 16594
rect 13556 15366 13584 17138
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13648 16454 13676 17002
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 15026 13584 15302
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 8566 13584 14962
rect 13648 9926 13676 16390
rect 13740 13258 13768 17326
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16590 13860 17070
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13924 14498 13952 19200
rect 14292 19122 14320 19200
rect 14384 19122 14412 19230
rect 14292 19094 14412 19122
rect 14464 18012 14516 18018
rect 14464 17954 14516 17960
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14476 16658 14504 17954
rect 14568 17814 14596 19230
rect 14646 19200 14702 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14476 16250 14504 16594
rect 14568 16561 14596 17750
rect 14660 17610 14688 19200
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14554 16552 14610 16561
rect 14554 16487 14610 16496
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 14660 15366 14688 16390
rect 14844 16046 14872 16458
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14648 15360 14700 15366
rect 14700 15308 14780 15314
rect 14648 15302 14780 15308
rect 14660 15286 14780 15302
rect 14280 15156 14332 15162
rect 14332 15116 14688 15144
rect 14280 15098 14332 15104
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 13832 14470 13952 14498
rect 13832 13734 13860 14470
rect 14476 14414 14504 14758
rect 14568 14482 14596 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 12322 13768 13194
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12442 13860 12786
rect 13924 12782 13952 14282
rect 14660 14278 14688 15116
rect 14752 15026 14780 15286
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14016 12628 14044 13466
rect 14476 13326 14504 14214
rect 14556 14000 14608 14006
rect 14554 13968 14556 13977
rect 14608 13968 14610 13977
rect 14554 13903 14610 13912
rect 14660 13870 14688 14214
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12714 14228 13126
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 13924 12600 14044 12628
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13740 12294 13860 12322
rect 13726 12200 13782 12209
rect 13726 12135 13782 12144
rect 13740 11762 13768 12135
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11558 13768 11698
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13832 10266 13860 12294
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9178 13676 9454
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 8634 13768 8774
rect 13832 8634 13860 9522
rect 13924 9194 13952 12600
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10742 14136 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10299 14376 10308
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9722 14320 9930
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 13924 9166 14044 9194
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13924 8430 13952 9046
rect 14016 8634 14044 9166
rect 14476 8922 14504 12718
rect 14660 12434 14688 13806
rect 14752 12782 14780 14962
rect 14844 14498 14872 15982
rect 14936 15042 14964 16934
rect 15028 16232 15056 19200
rect 15396 17218 15424 19200
rect 15474 17912 15530 17921
rect 15474 17847 15530 17856
rect 15304 17190 15424 17218
rect 15028 16204 15148 16232
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15028 15910 15056 16050
rect 15016 15904 15068 15910
rect 15014 15872 15016 15881
rect 15068 15872 15070 15881
rect 15014 15807 15070 15816
rect 14936 15014 15056 15042
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 14618 14964 14894
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14844 14470 14964 14498
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 13530 14872 14214
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14936 13326 14964 14470
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14844 12646 14872 12718
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14660 12406 14780 12434
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14568 10470 14596 12174
rect 14660 11694 14688 12242
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14660 11218 14688 11630
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9722 14596 9862
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14384 8894 14504 8922
rect 14648 8900 14700 8906
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8288 13872 8294
rect 14016 8242 14044 8570
rect 14384 8294 14412 8894
rect 14648 8842 14700 8848
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13924 8214 14044 8242
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13832 7886 13860 8026
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13924 7546 13952 8214
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14476 8090 14504 8774
rect 14568 8634 14596 8774
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14292 7546 14320 7958
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 13464 7398 13676 7426
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 6186 13492 7278
rect 13542 6896 13598 6905
rect 13542 6831 13598 6840
rect 13556 6798 13584 6831
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13556 6662 13584 6734
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13648 5914 13676 7398
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 6730 13768 7346
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13832 6458 13860 7142
rect 13924 6905 13952 7482
rect 14292 7290 14320 7482
rect 14292 7262 14504 7290
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14004 6928 14056 6934
rect 13910 6896 13966 6905
rect 14004 6870 14056 6876
rect 13910 6831 13966 6840
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13648 5302 13676 5850
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 4690 13492 5102
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4690 13676 4966
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13360 4616 13412 4622
rect 13740 4570 13768 6122
rect 13832 5574 13860 6258
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13360 4558 13412 4564
rect 13372 4282 13400 4558
rect 13648 4542 13768 4570
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13648 4214 13676 4542
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13372 2582 13400 3334
rect 13464 3194 13492 3334
rect 13556 3194 13584 3402
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13648 2582 13676 4150
rect 13832 4049 13860 5170
rect 13924 5098 13952 6734
rect 14016 6118 14044 6870
rect 14108 6186 14136 6938
rect 14476 6934 14504 7262
rect 14568 7002 14596 7822
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14464 6928 14516 6934
rect 14464 6870 14516 6876
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6338 14688 8842
rect 14752 8650 14780 12406
rect 14844 12306 14872 12582
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14936 10033 14964 13262
rect 15028 12986 15056 15014
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14922 10024 14978 10033
rect 14922 9959 14978 9968
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 9178 14964 9522
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14752 8634 14872 8650
rect 14752 8628 14884 8634
rect 14752 8622 14832 8628
rect 14752 8022 14780 8622
rect 14832 8570 14884 8576
rect 14936 8430 14964 8910
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14936 7954 14964 8366
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15028 7834 15056 12922
rect 15120 12442 15148 16204
rect 15304 15609 15332 17190
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15290 15600 15346 15609
rect 15290 15535 15346 15544
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15212 14890 15240 15302
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15120 12238 15148 12378
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 9042 15148 10066
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14936 7806 15056 7834
rect 15108 7812 15160 7818
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6798 14780 7142
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6390 14780 6598
rect 14568 6310 14688 6338
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14200 5370 14228 5850
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 14200 5030 14228 5102
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 14476 4622 14504 5646
rect 14568 5030 14596 6310
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14660 5846 14688 6190
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14660 4690 14688 5034
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14464 4616 14516 4622
rect 14556 4616 14608 4622
rect 14464 4558 14516 4564
rect 14554 4584 14556 4593
rect 14608 4584 14610 4593
rect 14554 4519 14610 4528
rect 13818 4040 13874 4049
rect 13818 3975 13874 3984
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13832 3074 13860 3975
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13924 3194 13952 3606
rect 14660 3602 14688 4626
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13648 2446 13676 2518
rect 13636 2440 13688 2446
rect 13280 2366 13400 2394
rect 13636 2382 13688 2388
rect 13082 2343 13138 2352
rect 13372 800 13400 2366
rect 13740 800 13768 3062
rect 13832 3046 13952 3074
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13832 2514 13860 2926
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13924 2394 13952 3046
rect 14108 2990 14136 3538
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14752 2774 14780 5850
rect 14844 3126 14872 7482
rect 14936 5914 14964 7806
rect 15108 7754 15160 7760
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 6390 15056 7686
rect 15120 7274 15148 7754
rect 15212 7750 15240 14826
rect 15304 11354 15332 15535
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 8974 15332 9454
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15396 7562 15424 17070
rect 15488 16658 15516 17847
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15764 15978 15792 19200
rect 16132 16182 16160 19200
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14482 15516 14894
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15476 14000 15528 14006
rect 15568 14000 15620 14006
rect 15476 13942 15528 13948
rect 15566 13968 15568 13977
rect 15620 13968 15622 13977
rect 15488 13530 15516 13942
rect 15566 13903 15622 13912
rect 15580 13530 15608 13903
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15304 7534 15424 7562
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15120 6934 15148 7210
rect 15304 7206 15332 7534
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 15120 6254 15148 6870
rect 15304 6662 15332 7142
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15212 5778 15240 6015
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14936 4468 14964 4966
rect 15106 4856 15162 4865
rect 15106 4791 15108 4800
rect 15160 4791 15162 4800
rect 15108 4762 15160 4768
rect 14936 4440 15056 4468
rect 14922 4040 14978 4049
rect 14922 3975 14978 3984
rect 14936 3194 14964 3975
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14936 3058 14964 3130
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14752 2746 14872 2774
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 13924 2366 14136 2394
rect 14108 800 14136 2366
rect 14464 1488 14516 1494
rect 14464 1430 14516 1436
rect 14476 800 14504 1430
rect 14844 800 14872 2746
rect 14936 2650 14964 2994
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15028 1834 15056 4440
rect 15304 3534 15332 6598
rect 15396 6458 15424 7346
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6322 15516 9930
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 5914 15516 6258
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15198 2952 15254 2961
rect 15198 2887 15254 2896
rect 15016 1828 15068 1834
rect 15016 1770 15068 1776
rect 15212 800 15240 2887
rect 15488 2774 15516 5850
rect 15580 2961 15608 11494
rect 15764 8974 15792 15914
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8634 15792 8910
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15764 8090 15792 8570
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15764 7546 15792 8026
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15936 2984 15988 2990
rect 15566 2952 15622 2961
rect 15936 2926 15988 2932
rect 15566 2887 15622 2896
rect 15488 2746 15608 2774
rect 15580 800 15608 2746
rect 15948 800 15976 2926
rect 11992 734 12204 762
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
<< via2 >>
rect 1674 19080 1730 19136
rect 1766 16632 1822 16688
rect 2042 16532 2044 16552
rect 2044 16532 2096 16552
rect 2096 16532 2098 16552
rect 2042 16496 2098 16532
rect 2318 17584 2374 17640
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 1674 14728 1730 14784
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 1766 13776 1822 13832
rect 1674 12824 1730 12880
rect 1766 11872 1822 11928
rect 1674 10920 1730 10976
rect 2226 10004 2228 10024
rect 2228 10004 2280 10024
rect 2280 10004 2282 10024
rect 2226 9968 2282 10004
rect 3330 15564 3386 15600
rect 3330 15544 3332 15564
rect 3332 15544 3384 15564
rect 3384 15544 3386 15564
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 3330 13776 3386 13832
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 3330 11092 3332 11112
rect 3332 11092 3384 11112
rect 3384 11092 3386 11112
rect 3330 11056 3386 11092
rect 1398 4256 1454 4312
rect 1582 9016 1638 9072
rect 1674 8064 1730 8120
rect 1582 7112 1638 7168
rect 1674 5208 1730 5264
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2594 6160 2650 6216
rect 1490 856 1546 912
rect 2318 3304 2374 3360
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 3330 8200 3386 8256
rect 3330 5228 3386 5264
rect 3330 5208 3332 5228
rect 3332 5208 3384 5228
rect 3384 5208 3386 5228
rect 3238 4528 3294 4584
rect 3146 4120 3202 4176
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 3330 3576 3386 3632
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 4066 18536 4122 18592
rect 3790 15408 3846 15464
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 5078 15136 5134 15192
rect 4894 14864 4950 14920
rect 5446 16088 5502 16144
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 3882 12180 3884 12200
rect 3884 12180 3936 12200
rect 3936 12180 3938 12200
rect 3882 12144 3938 12180
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 3974 5616 4030 5672
rect 3330 1400 3386 1456
rect 4158 3032 4214 3088
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4618 5616 4674 5672
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6182 13912 6238 13968
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 5446 3984 5502 4040
rect 4986 3460 5042 3496
rect 4986 3440 4988 3460
rect 4988 3440 5040 3460
rect 5040 3440 5042 3460
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 3974 2644 4030 2680
rect 3974 2624 3976 2644
rect 3976 2624 4028 2644
rect 4028 2624 4030 2644
rect 5170 3340 5172 3360
rect 5172 3340 5224 3360
rect 5224 3340 5226 3360
rect 5170 3304 5226 3340
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 6090 4684 6146 4720
rect 6090 4664 6092 4684
rect 6092 4664 6144 4684
rect 6144 4664 6146 4684
rect 5906 3440 5962 3496
rect 5814 3032 5870 3088
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8114 15988 8116 16008
rect 8116 15988 8168 16008
rect 8168 15988 8170 16008
rect 7470 15544 7526 15600
rect 8114 15952 8170 15988
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6734 5752 6790 5808
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 5814 2524 5816 2544
rect 5816 2524 5868 2544
rect 5868 2524 5870 2544
rect 5814 2488 5870 2524
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 7010 3304 7066 3360
rect 6734 2896 6790 2952
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7562 2760 7618 2816
rect 7838 5752 7894 5808
rect 7746 3712 7802 3768
rect 9218 16224 9274 16280
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8758 10512 8814 10568
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 7654 2488 7710 2544
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8206 3712 8262 3768
rect 8850 3576 8906 3632
rect 8206 3168 8262 3224
rect 8206 3032 8262 3088
rect 8850 3304 8906 3360
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 9586 16532 9588 16552
rect 9588 16532 9640 16552
rect 9640 16532 9642 16552
rect 9586 16496 9642 16532
rect 10874 17212 10876 17232
rect 10876 17212 10928 17232
rect 10928 17212 10930 17232
rect 10874 17176 10930 17212
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10138 15952 10194 16008
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 11150 16088 11206 16144
rect 10598 15308 10600 15328
rect 10600 15308 10652 15328
rect 10652 15308 10654 15328
rect 10598 15272 10654 15308
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 9954 4820 10010 4856
rect 9954 4800 9956 4820
rect 9956 4800 10008 4820
rect 10008 4800 10010 4820
rect 9862 4528 9918 4584
rect 9218 2896 9274 2952
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9954 3068 9956 3088
rect 9956 3068 10008 3088
rect 10008 3068 10010 3088
rect 9954 3032 10010 3068
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 11518 16360 11574 16416
rect 10874 15000 10930 15056
rect 10966 13776 11022 13832
rect 11334 14864 11390 14920
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 11334 9016 11390 9072
rect 11150 3984 11206 4040
rect 10322 3032 10378 3088
rect 9862 2352 9918 2408
rect 10046 2216 10102 2272
rect 10598 2896 10654 2952
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 10966 3052 11022 3088
rect 10966 3032 10968 3052
rect 10968 3032 11020 3052
rect 11020 3032 11022 3052
rect 11242 3440 11298 3496
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12070 15816 12126 15872
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 13266 15000 13322 15056
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12714 9968 12770 10024
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12806 8356 12862 8392
rect 12806 8336 12808 8356
rect 12808 8336 12860 8356
rect 12860 8336 12862 8356
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 11610 5208 11666 5264
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 11242 2760 11298 2816
rect 11518 2760 11574 2816
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12070 4120 12126 4176
rect 12070 3984 12126 4040
rect 12346 3712 12402 3768
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12346 3032 12402 3088
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12714 2080 12770 2136
rect 13174 9016 13230 9072
rect 13082 2388 13084 2408
rect 13084 2388 13136 2408
rect 13136 2388 13138 2408
rect 13082 2352 13138 2388
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14554 16496 14610 16552
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14554 13948 14556 13968
rect 14556 13948 14608 13968
rect 14608 13948 14610 13968
rect 14554 13912 14610 13948
rect 13726 12144 13782 12200
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 15474 17856 15530 17912
rect 15014 15852 15016 15872
rect 15016 15852 15068 15872
rect 15068 15852 15070 15872
rect 15014 15816 15070 15852
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 13542 6840 13598 6896
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 13910 6840 13966 6896
rect 14922 9968 14978 10024
rect 15290 15544 15346 15600
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14554 4564 14556 4584
rect 14556 4564 14608 4584
rect 14608 4564 14610 4584
rect 14554 4528 14610 4564
rect 13818 3984 13874 4040
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 15566 13948 15568 13968
rect 15568 13948 15620 13968
rect 15620 13948 15622 13968
rect 15566 13912 15622 13948
rect 15198 6024 15254 6080
rect 15106 4820 15162 4856
rect 15106 4800 15108 4820
rect 15108 4800 15160 4820
rect 15160 4800 15162 4820
rect 14922 3984 14978 4040
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 15198 2896 15254 2952
rect 15566 2896 15622 2952
<< metal3 >>
rect 0 19546 800 19576
rect 0 19486 1042 19546
rect 0 19456 800 19486
rect 982 19138 1042 19486
rect 1669 19138 1735 19141
rect 982 19136 1735 19138
rect 982 19080 1674 19136
rect 1730 19080 1735 19136
rect 982 19078 1735 19080
rect 1669 19075 1735 19078
rect 0 18594 800 18624
rect 4061 18594 4127 18597
rect 0 18592 4127 18594
rect 0 18536 4066 18592
rect 4122 18536 4127 18592
rect 0 18534 4127 18536
rect 0 18504 800 18534
rect 4061 18531 4127 18534
rect 15469 17914 15535 17917
rect 16400 17914 17200 17944
rect 15469 17912 17200 17914
rect 15469 17856 15474 17912
rect 15530 17856 17200 17912
rect 15469 17854 17200 17856
rect 15469 17851 15535 17854
rect 16400 17824 17200 17854
rect 0 17642 800 17672
rect 2313 17642 2379 17645
rect 0 17640 2379 17642
rect 0 17584 2318 17640
rect 2374 17584 2379 17640
rect 0 17582 2379 17584
rect 0 17552 800 17582
rect 2313 17579 2379 17582
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 10726 17172 10732 17236
rect 10796 17234 10802 17236
rect 10869 17234 10935 17237
rect 10796 17232 10935 17234
rect 10796 17176 10874 17232
rect 10930 17176 10935 17232
rect 10796 17174 10935 17176
rect 10796 17172 10802 17174
rect 10869 17171 10935 17174
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 0 16690 800 16720
rect 1761 16690 1827 16693
rect 0 16688 1827 16690
rect 0 16632 1766 16688
rect 1822 16632 1827 16688
rect 0 16630 1827 16632
rect 0 16600 800 16630
rect 1761 16627 1827 16630
rect 2037 16554 2103 16557
rect 2037 16552 9322 16554
rect 2037 16496 2042 16552
rect 2098 16496 9322 16552
rect 2037 16494 9322 16496
rect 2037 16491 2103 16494
rect 9262 16418 9322 16494
rect 9438 16492 9444 16556
rect 9508 16554 9514 16556
rect 9581 16554 9647 16557
rect 9508 16552 9647 16554
rect 9508 16496 9586 16552
rect 9642 16496 9647 16552
rect 9508 16494 9647 16496
rect 9508 16492 9514 16494
rect 9581 16491 9647 16494
rect 14549 16554 14615 16557
rect 14774 16554 14780 16556
rect 14549 16552 14780 16554
rect 14549 16496 14554 16552
rect 14610 16496 14780 16552
rect 14549 16494 14780 16496
rect 14549 16491 14615 16494
rect 14774 16492 14780 16494
rect 14844 16492 14850 16556
rect 11513 16418 11579 16421
rect 9262 16416 11579 16418
rect 9262 16360 11518 16416
rect 11574 16360 11579 16416
rect 9262 16358 11579 16360
rect 11513 16355 11579 16358
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 9213 16284 9279 16285
rect 9213 16282 9260 16284
rect 9168 16280 9260 16282
rect 9168 16224 9218 16280
rect 9168 16222 9260 16224
rect 9213 16220 9260 16222
rect 9324 16220 9330 16284
rect 9213 16219 9279 16220
rect 5441 16146 5507 16149
rect 11145 16146 11211 16149
rect 5441 16144 11211 16146
rect 5441 16088 5446 16144
rect 5502 16088 11150 16144
rect 11206 16088 11211 16144
rect 5441 16086 11211 16088
rect 5441 16083 5507 16086
rect 11145 16083 11211 16086
rect 8109 16010 8175 16013
rect 10133 16010 10199 16013
rect 8109 16008 10199 16010
rect 8109 15952 8114 16008
rect 8170 15952 10138 16008
rect 10194 15952 10199 16008
rect 8109 15950 10199 15952
rect 8109 15947 8175 15950
rect 10133 15947 10199 15950
rect 12065 15876 12131 15877
rect 15009 15876 15075 15877
rect 12014 15874 12020 15876
rect 11974 15814 12020 15874
rect 12084 15872 12131 15876
rect 12126 15816 12131 15872
rect 12014 15812 12020 15814
rect 12084 15812 12131 15816
rect 14958 15812 14964 15876
rect 15028 15874 15075 15876
rect 15028 15872 15120 15874
rect 15070 15816 15120 15872
rect 15028 15814 15120 15816
rect 15028 15812 15075 15814
rect 12065 15811 12131 15812
rect 15009 15811 15075 15812
rect 2820 15808 3136 15809
rect 0 15738 800 15768
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 0 15678 2698 15738
rect 0 15648 800 15678
rect 2638 15602 2698 15678
rect 3325 15602 3391 15605
rect 2638 15600 3391 15602
rect 2638 15544 3330 15600
rect 3386 15544 3391 15600
rect 2638 15542 3391 15544
rect 3325 15539 3391 15542
rect 7465 15602 7531 15605
rect 7782 15602 7788 15604
rect 7465 15600 7788 15602
rect 7465 15544 7470 15600
rect 7526 15544 7788 15600
rect 7465 15542 7788 15544
rect 7465 15539 7531 15542
rect 7782 15540 7788 15542
rect 7852 15602 7858 15604
rect 15285 15602 15351 15605
rect 7852 15600 15351 15602
rect 7852 15544 15290 15600
rect 15346 15544 15351 15600
rect 7852 15542 15351 15544
rect 7852 15540 7858 15542
rect 15285 15539 15351 15542
rect 3785 15466 3851 15469
rect 3785 15464 10242 15466
rect 3785 15408 3790 15464
rect 3846 15408 10242 15464
rect 3785 15406 10242 15408
rect 3785 15403 3851 15406
rect 10182 15332 10242 15406
rect 10174 15268 10180 15332
rect 10244 15330 10250 15332
rect 10593 15330 10659 15333
rect 10244 15328 10659 15330
rect 10244 15272 10598 15328
rect 10654 15272 10659 15328
rect 10244 15270 10659 15272
rect 10244 15268 10250 15270
rect 10593 15267 10659 15270
rect 4694 15264 5010 15265
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 5073 15194 5139 15197
rect 5073 15192 8218 15194
rect 5073 15136 5078 15192
rect 5134 15136 8218 15192
rect 5073 15134 8218 15136
rect 5073 15131 5139 15134
rect 8158 15058 8218 15134
rect 10869 15058 10935 15061
rect 8158 15056 10935 15058
rect 8158 15000 10874 15056
rect 10930 15000 10935 15056
rect 8158 14998 10935 15000
rect 10869 14995 10935 14998
rect 11094 14996 11100 15060
rect 11164 15058 11170 15060
rect 13261 15058 13327 15061
rect 11164 15056 13327 15058
rect 11164 15000 13266 15056
rect 13322 15000 13327 15056
rect 11164 14998 13327 15000
rect 11164 14996 11170 14998
rect 13261 14995 13327 14998
rect 4889 14922 4955 14925
rect 11329 14922 11395 14925
rect 4889 14920 11395 14922
rect 4889 14864 4894 14920
rect 4950 14864 11334 14920
rect 11390 14864 11395 14920
rect 4889 14862 11395 14864
rect 4889 14859 4955 14862
rect 11329 14859 11395 14862
rect 0 14786 800 14816
rect 1669 14786 1735 14789
rect 0 14784 1735 14786
rect 0 14728 1674 14784
rect 1730 14728 1735 14784
rect 0 14726 1735 14728
rect 0 14696 800 14726
rect 1669 14723 1735 14726
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 6177 13970 6243 13973
rect 14549 13970 14615 13973
rect 6177 13968 14615 13970
rect 6177 13912 6182 13968
rect 6238 13912 14554 13968
rect 14610 13912 14615 13968
rect 6177 13910 14615 13912
rect 6177 13907 6243 13910
rect 14549 13907 14615 13910
rect 15561 13970 15627 13973
rect 16400 13970 17200 14000
rect 15561 13968 17200 13970
rect 15561 13912 15566 13968
rect 15622 13912 17200 13968
rect 15561 13910 17200 13912
rect 15561 13907 15627 13910
rect 16400 13880 17200 13910
rect 0 13834 800 13864
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 3325 13834 3391 13837
rect 10961 13834 11027 13837
rect 3325 13832 11027 13834
rect 3325 13776 3330 13832
rect 3386 13776 10966 13832
rect 11022 13776 11027 13832
rect 3325 13774 11027 13776
rect 3325 13771 3391 13774
rect 10961 13771 11027 13774
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 0 12882 800 12912
rect 1669 12882 1735 12885
rect 0 12880 1735 12882
rect 0 12824 1674 12880
rect 1730 12824 1735 12880
rect 0 12822 1735 12824
rect 0 12792 800 12822
rect 1669 12819 1735 12822
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 3877 12204 3943 12205
rect 3877 12202 3924 12204
rect 3832 12200 3924 12202
rect 3832 12144 3882 12200
rect 3832 12142 3924 12144
rect 3877 12140 3924 12142
rect 3988 12140 3994 12204
rect 9254 12140 9260 12204
rect 9324 12202 9330 12204
rect 13721 12202 13787 12205
rect 9324 12200 13787 12202
rect 9324 12144 13726 12200
rect 13782 12144 13787 12200
rect 9324 12142 13787 12144
rect 9324 12140 9330 12142
rect 3877 12139 3943 12140
rect 13721 12139 13787 12142
rect 4694 12000 5010 12001
rect 0 11930 800 11960
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 1761 11930 1827 11933
rect 0 11928 1827 11930
rect 0 11872 1766 11928
rect 1822 11872 1827 11928
rect 0 11870 1827 11872
rect 0 11840 800 11870
rect 1761 11867 1827 11870
rect 2820 11456 3136 11457
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 3325 11116 3391 11117
rect 3325 11114 3372 11116
rect 3280 11112 3372 11114
rect 3280 11056 3330 11112
rect 3280 11054 3372 11056
rect 3325 11052 3372 11054
rect 3436 11052 3442 11116
rect 3325 11051 3391 11052
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 8753 10570 8819 10573
rect 11094 10570 11100 10572
rect 8753 10568 11100 10570
rect 8753 10512 8758 10568
rect 8814 10512 11100 10568
rect 8753 10510 11100 10512
rect 8753 10507 8819 10510
rect 11094 10508 11100 10510
rect 11164 10508 11170 10572
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 0 10026 800 10056
rect 2221 10026 2287 10029
rect 0 10024 2287 10026
rect 0 9968 2226 10024
rect 2282 9968 2287 10024
rect 0 9966 2287 9968
rect 0 9936 800 9966
rect 2221 9963 2287 9966
rect 12014 9964 12020 10028
rect 12084 10026 12090 10028
rect 12709 10026 12775 10029
rect 12084 10024 12775 10026
rect 12084 9968 12714 10024
rect 12770 9968 12775 10024
rect 12084 9966 12775 9968
rect 12084 9964 12090 9966
rect 12709 9963 12775 9966
rect 14917 10026 14983 10029
rect 16400 10026 17200 10056
rect 14917 10024 17200 10026
rect 14917 9968 14922 10024
rect 14978 9968 17200 10024
rect 14917 9966 17200 9968
rect 14917 9963 14983 9966
rect 16400 9936 17200 9966
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 9438 9556 9444 9620
rect 9508 9618 9514 9620
rect 12566 9618 12572 9620
rect 9508 9558 12572 9618
rect 9508 9556 9514 9558
rect 12566 9556 12572 9558
rect 12636 9556 12642 9620
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 0 9074 800 9104
rect 1577 9074 1643 9077
rect 0 9072 1643 9074
rect 0 9016 1582 9072
rect 1638 9016 1643 9072
rect 0 9014 1643 9016
rect 0 8984 800 9014
rect 1577 9011 1643 9014
rect 11329 9074 11395 9077
rect 13169 9074 13235 9077
rect 11329 9072 13235 9074
rect 11329 9016 11334 9072
rect 11390 9016 13174 9072
rect 13230 9016 13235 9072
rect 11329 9014 13235 9016
rect 11329 9011 11395 9014
rect 13169 9011 13235 9014
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 12566 8332 12572 8396
rect 12636 8394 12642 8396
rect 12801 8394 12867 8397
rect 12636 8392 12867 8394
rect 12636 8336 12806 8392
rect 12862 8336 12867 8392
rect 12636 8334 12867 8336
rect 12636 8332 12642 8334
rect 12801 8331 12867 8334
rect 3325 8260 3391 8261
rect 3325 8256 3372 8260
rect 3436 8258 3442 8260
rect 3325 8200 3330 8256
rect 3325 8196 3372 8200
rect 3436 8198 3482 8258
rect 3436 8196 3442 8198
rect 3325 8195 3391 8196
rect 2820 8192 3136 8193
rect 0 8122 800 8152
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 1669 8122 1735 8125
rect 0 8120 1735 8122
rect 0 8064 1674 8120
rect 1730 8064 1735 8120
rect 0 8062 1735 8064
rect 0 8032 800 8062
rect 1669 8059 1735 8062
rect 4694 7648 5010 7649
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 0 7170 800 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 800 7110
rect 1577 7107 1643 7110
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 13537 6898 13603 6901
rect 13905 6898 13971 6901
rect 13537 6896 13971 6898
rect 13537 6840 13542 6896
rect 13598 6840 13910 6896
rect 13966 6840 13971 6896
rect 13537 6838 13971 6840
rect 13537 6835 13603 6838
rect 13905 6835 13971 6838
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 0 6218 800 6248
rect 2589 6218 2655 6221
rect 0 6216 2655 6218
rect 0 6160 2594 6216
rect 2650 6160 2655 6216
rect 0 6158 2655 6160
rect 0 6128 800 6158
rect 2589 6155 2655 6158
rect 15193 6082 15259 6085
rect 16400 6082 17200 6112
rect 15193 6080 17200 6082
rect 15193 6024 15198 6080
rect 15254 6024 17200 6080
rect 15193 6022 17200 6024
rect 15193 6019 15259 6022
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 16400 5992 17200 6022
rect 14064 5951 14380 5952
rect 6729 5810 6795 5813
rect 7833 5810 7899 5813
rect 6729 5808 7899 5810
rect 6729 5752 6734 5808
rect 6790 5752 7838 5808
rect 7894 5752 7899 5808
rect 6729 5750 7899 5752
rect 6729 5747 6795 5750
rect 7833 5747 7899 5750
rect 3969 5674 4035 5677
rect 4613 5674 4679 5677
rect 3969 5672 4679 5674
rect 3969 5616 3974 5672
rect 4030 5616 4618 5672
rect 4674 5616 4679 5672
rect 3969 5614 4679 5616
rect 3969 5611 4035 5614
rect 4613 5611 4679 5614
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 0 5266 800 5296
rect 1669 5266 1735 5269
rect 0 5264 1735 5266
rect 0 5208 1674 5264
rect 1730 5208 1735 5264
rect 0 5206 1735 5208
rect 0 5176 800 5206
rect 1669 5203 1735 5206
rect 3325 5266 3391 5269
rect 11605 5266 11671 5269
rect 3325 5264 11671 5266
rect 3325 5208 3330 5264
rect 3386 5208 11610 5264
rect 11666 5208 11671 5264
rect 3325 5206 11671 5208
rect 3325 5203 3391 5206
rect 11605 5203 11671 5206
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 9949 4860 10015 4861
rect 9949 4856 9996 4860
rect 10060 4858 10066 4860
rect 9949 4800 9954 4856
rect 9949 4796 9996 4800
rect 10060 4798 10106 4858
rect 10060 4796 10066 4798
rect 14774 4796 14780 4860
rect 14844 4858 14850 4860
rect 15101 4858 15167 4861
rect 14844 4856 15167 4858
rect 14844 4800 15106 4856
rect 15162 4800 15167 4856
rect 14844 4798 15167 4800
rect 14844 4796 14850 4798
rect 9949 4795 10015 4796
rect 15101 4795 15167 4798
rect 6085 4722 6151 4725
rect 6085 4720 12450 4722
rect 6085 4664 6090 4720
rect 6146 4664 12450 4720
rect 6085 4662 12450 4664
rect 6085 4659 6151 4662
rect 3233 4586 3299 4589
rect 9857 4586 9923 4589
rect 3233 4584 9923 4586
rect 3233 4528 3238 4584
rect 3294 4528 9862 4584
rect 9918 4528 9923 4584
rect 3233 4526 9923 4528
rect 12390 4586 12450 4662
rect 14549 4586 14615 4589
rect 12390 4584 14615 4586
rect 12390 4528 14554 4584
rect 14610 4528 14615 4584
rect 12390 4526 14615 4528
rect 3233 4523 3299 4526
rect 9857 4523 9923 4526
rect 14549 4523 14615 4526
rect 4694 4384 5010 4385
rect 0 4314 800 4344
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 1393 4314 1459 4317
rect 0 4312 1459 4314
rect 0 4256 1398 4312
rect 1454 4256 1459 4312
rect 0 4254 1459 4256
rect 0 4224 800 4254
rect 1393 4251 1459 4254
rect 3141 4178 3207 4181
rect 12065 4178 12131 4181
rect 3141 4176 12131 4178
rect 3141 4120 3146 4176
rect 3202 4120 12070 4176
rect 12126 4120 12131 4176
rect 3141 4118 12131 4120
rect 3141 4115 3207 4118
rect 12065 4115 12131 4118
rect 5441 4042 5507 4045
rect 11145 4042 11211 4045
rect 12065 4042 12131 4045
rect 13813 4042 13879 4045
rect 14917 4044 14983 4045
rect 14917 4042 14964 4044
rect 5441 4040 11211 4042
rect 5441 3984 5446 4040
rect 5502 3984 11150 4040
rect 11206 3984 11211 4040
rect 5441 3982 11211 3984
rect 5441 3979 5507 3982
rect 11145 3979 11211 3982
rect 11286 4040 12131 4042
rect 11286 3984 12070 4040
rect 12126 3984 12131 4040
rect 11286 3982 12131 3984
rect 2820 3840 3136 3841
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 7741 3772 7807 3773
rect 7741 3770 7788 3772
rect 7696 3768 7788 3770
rect 7696 3712 7746 3768
rect 7696 3710 7788 3712
rect 7741 3708 7788 3710
rect 7852 3708 7858 3772
rect 8201 3770 8267 3773
rect 8201 3768 9138 3770
rect 8201 3712 8206 3768
rect 8262 3712 9138 3768
rect 8201 3710 9138 3712
rect 7741 3707 7807 3708
rect 8201 3707 8267 3710
rect 3325 3634 3391 3637
rect 8845 3634 8911 3637
rect 3325 3632 8911 3634
rect 3325 3576 3330 3632
rect 3386 3576 8850 3632
rect 8906 3576 8911 3632
rect 3325 3574 8911 3576
rect 9078 3634 9138 3710
rect 11286 3634 11346 3982
rect 12065 3979 12131 3982
rect 12390 4040 13879 4042
rect 12390 3984 13818 4040
rect 13874 3984 13879 4040
rect 12390 3982 13879 3984
rect 14872 4040 14964 4042
rect 14872 3984 14922 4040
rect 14872 3982 14964 3984
rect 12390 3906 12450 3982
rect 13813 3979 13879 3982
rect 14917 3980 14964 3982
rect 15028 3980 15034 4044
rect 14917 3979 14983 3980
rect 9078 3574 11346 3634
rect 11470 3846 12450 3906
rect 3325 3571 3391 3574
rect 8845 3571 8911 3574
rect 4981 3498 5047 3501
rect 5901 3498 5967 3501
rect 11237 3498 11303 3501
rect 4981 3496 11303 3498
rect 4981 3440 4986 3496
rect 5042 3440 5906 3496
rect 5962 3440 11242 3496
rect 11298 3440 11303 3496
rect 4981 3438 11303 3440
rect 4981 3435 5047 3438
rect 5901 3435 5967 3438
rect 11237 3435 11303 3438
rect 0 3362 800 3392
rect 2313 3362 2379 3365
rect 0 3360 2379 3362
rect 0 3304 2318 3360
rect 2374 3304 2379 3360
rect 0 3302 2379 3304
rect 0 3272 800 3302
rect 2313 3299 2379 3302
rect 5165 3362 5231 3365
rect 7005 3362 7071 3365
rect 5165 3360 7071 3362
rect 5165 3304 5170 3360
rect 5226 3304 7010 3360
rect 7066 3304 7071 3360
rect 5165 3302 7071 3304
rect 5165 3299 5231 3302
rect 7005 3299 7071 3302
rect 8845 3362 8911 3365
rect 11470 3362 11530 3846
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 12341 3770 12407 3773
rect 12566 3770 12572 3772
rect 12341 3768 12572 3770
rect 12341 3712 12346 3768
rect 12402 3712 12572 3768
rect 12341 3710 12572 3712
rect 12341 3707 12407 3710
rect 12566 3708 12572 3710
rect 12636 3708 12642 3772
rect 8845 3360 11530 3362
rect 8845 3304 8850 3360
rect 8906 3304 11530 3360
rect 8845 3302 11530 3304
rect 8845 3299 8911 3302
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 12190 3231 12506 3232
rect 8201 3226 8267 3229
rect 5214 3224 8267 3226
rect 5214 3168 8206 3224
rect 8262 3168 8267 3224
rect 5214 3166 8267 3168
rect 4153 3090 4219 3093
rect 5214 3090 5274 3166
rect 8201 3163 8267 3166
rect 8894 3166 11162 3226
rect 4153 3088 5274 3090
rect 4153 3032 4158 3088
rect 4214 3032 5274 3088
rect 4153 3030 5274 3032
rect 5809 3090 5875 3093
rect 8201 3090 8267 3093
rect 8894 3090 8954 3166
rect 5809 3088 7482 3090
rect 5809 3032 5814 3088
rect 5870 3032 7482 3088
rect 5809 3030 7482 3032
rect 4153 3027 4219 3030
rect 5809 3027 5875 3030
rect 6729 2954 6795 2957
rect 7422 2954 7482 3030
rect 8201 3088 8954 3090
rect 8201 3032 8206 3088
rect 8262 3032 8954 3088
rect 8201 3030 8954 3032
rect 9949 3090 10015 3093
rect 10317 3090 10383 3093
rect 9949 3088 10383 3090
rect 9949 3032 9954 3088
rect 10010 3032 10322 3088
rect 10378 3032 10383 3088
rect 9949 3030 10383 3032
rect 8201 3027 8267 3030
rect 9949 3027 10015 3030
rect 10317 3027 10383 3030
rect 10726 3028 10732 3092
rect 10796 3090 10802 3092
rect 10961 3090 11027 3093
rect 10796 3088 11027 3090
rect 10796 3032 10966 3088
rect 11022 3032 11027 3088
rect 10796 3030 11027 3032
rect 11102 3090 11162 3166
rect 12341 3090 12407 3093
rect 11102 3088 12407 3090
rect 11102 3032 12346 3088
rect 12402 3032 12407 3088
rect 11102 3030 12407 3032
rect 10796 3028 10802 3030
rect 10961 3027 11027 3030
rect 12341 3027 12407 3030
rect 9213 2954 9279 2957
rect 6729 2952 7114 2954
rect 6729 2896 6734 2952
rect 6790 2896 7114 2952
rect 6729 2894 7114 2896
rect 7422 2952 9279 2954
rect 7422 2896 9218 2952
rect 9274 2896 9279 2952
rect 7422 2894 9279 2896
rect 6729 2891 6795 2894
rect 7054 2818 7114 2894
rect 9213 2891 9279 2894
rect 10174 2892 10180 2956
rect 10244 2954 10250 2956
rect 10593 2954 10659 2957
rect 15193 2954 15259 2957
rect 15561 2954 15627 2957
rect 10244 2952 10659 2954
rect 10244 2896 10598 2952
rect 10654 2896 10659 2952
rect 10244 2894 10659 2896
rect 10244 2892 10250 2894
rect 10593 2891 10659 2894
rect 10734 2952 15627 2954
rect 10734 2896 15198 2952
rect 15254 2896 15566 2952
rect 15622 2896 15627 2952
rect 10734 2894 15627 2896
rect 7557 2818 7623 2821
rect 7054 2816 10242 2818
rect 7054 2760 7562 2816
rect 7618 2760 10242 2816
rect 7054 2758 10242 2760
rect 7557 2755 7623 2758
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 3969 2684 4035 2685
rect 3918 2682 3924 2684
rect 3878 2622 3924 2682
rect 3988 2680 4035 2684
rect 4030 2624 4035 2680
rect 3918 2620 3924 2622
rect 3988 2620 4035 2624
rect 3926 2619 4035 2620
rect 0 2410 800 2440
rect 3926 2410 3986 2619
rect 5809 2546 5875 2549
rect 7649 2546 7715 2549
rect 5809 2544 7715 2546
rect 5809 2488 5814 2544
rect 5870 2488 7654 2544
rect 7710 2488 7715 2544
rect 5809 2486 7715 2488
rect 10182 2546 10242 2758
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 10734 2546 10794 2894
rect 15193 2891 15259 2894
rect 15561 2891 15627 2894
rect 11237 2818 11303 2821
rect 11513 2818 11579 2821
rect 11237 2816 11579 2818
rect 11237 2760 11242 2816
rect 11298 2760 11518 2816
rect 11574 2760 11579 2816
rect 11237 2758 11579 2760
rect 11237 2755 11303 2758
rect 11513 2755 11579 2758
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 10182 2486 10794 2546
rect 5809 2483 5875 2486
rect 7649 2483 7715 2486
rect 0 2350 3986 2410
rect 9857 2410 9923 2413
rect 13077 2410 13143 2413
rect 9857 2408 13143 2410
rect 9857 2352 9862 2408
rect 9918 2352 13082 2408
rect 13138 2352 13143 2408
rect 9857 2350 13143 2352
rect 0 2320 800 2350
rect 9857 2347 9923 2350
rect 13077 2347 13143 2350
rect 10041 2276 10107 2277
rect 9990 2212 9996 2276
rect 10060 2274 10107 2276
rect 10060 2272 10152 2274
rect 10102 2216 10152 2272
rect 10060 2214 10152 2216
rect 10060 2212 10107 2214
rect 10041 2211 10107 2212
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 12709 2138 12775 2141
rect 16400 2138 17200 2168
rect 12709 2136 17200 2138
rect 12709 2080 12714 2136
rect 12770 2080 17200 2136
rect 12709 2078 17200 2080
rect 12709 2075 12775 2078
rect 16400 2048 17200 2078
rect 0 1458 800 1488
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1368 800 1398
rect 3325 1395 3391 1398
rect 1485 914 1551 917
rect 982 912 1551 914
rect 982 856 1490 912
rect 1546 856 1551 912
rect 982 854 1551 856
rect 0 506 800 536
rect 982 506 1042 854
rect 1485 851 1551 854
rect 0 446 1042 506
rect 0 416 800 446
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 10732 17172 10796 17236
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 9444 16492 9508 16556
rect 14780 16492 14844 16556
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 9260 16280 9324 16284
rect 9260 16224 9274 16280
rect 9274 16224 9324 16280
rect 9260 16220 9324 16224
rect 12020 15872 12084 15876
rect 12020 15816 12070 15872
rect 12070 15816 12084 15872
rect 12020 15812 12084 15816
rect 14964 15872 15028 15876
rect 14964 15816 15014 15872
rect 15014 15816 15028 15872
rect 14964 15812 15028 15816
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 7788 15540 7852 15604
rect 10180 15268 10244 15332
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 11100 14996 11164 15060
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 3924 12200 3988 12204
rect 3924 12144 3938 12200
rect 3938 12144 3988 12200
rect 3924 12140 3988 12144
rect 9260 12140 9324 12204
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 3372 11112 3436 11116
rect 3372 11056 3386 11112
rect 3386 11056 3436 11112
rect 3372 11052 3436 11056
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 11100 10508 11164 10572
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 12020 9964 12084 10028
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 9444 9556 9508 9620
rect 12572 9556 12636 9620
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 12572 8332 12636 8396
rect 3372 8256 3436 8260
rect 3372 8200 3386 8256
rect 3386 8200 3436 8256
rect 3372 8196 3436 8200
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 9996 4856 10060 4860
rect 9996 4800 10010 4856
rect 10010 4800 10060 4856
rect 9996 4796 10060 4800
rect 14780 4796 14844 4860
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 7788 3768 7852 3772
rect 7788 3712 7802 3768
rect 7802 3712 7852 3768
rect 7788 3708 7852 3712
rect 14964 4040 15028 4044
rect 14964 3984 14978 4040
rect 14978 3984 15028 4040
rect 14964 3980 15028 3984
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 12572 3708 12636 3772
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 10732 3028 10796 3092
rect 10180 2892 10244 2956
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 3924 2680 3988 2684
rect 3924 2624 3974 2680
rect 3974 2624 3988 2680
rect 3924 2620 3988 2624
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 9996 2272 10060 2276
rect 9996 2216 10046 2272
rect 10046 2216 10060 2272
rect 9996 2212 10060 2216
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 3923 12204 3989 12205
rect 3923 12140 3924 12204
rect 3988 12140 3989 12204
rect 3923 12139 3989 12140
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 3374 8261 3434 11051
rect 3371 8260 3437 8261
rect 3371 8196 3372 8260
rect 3436 8196 3437 8260
rect 3371 8195 3437 8196
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 3926 2685 3986 12139
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 3923 2684 3989 2685
rect 3923 2620 3924 2684
rect 3988 2620 3989 2684
rect 3923 2619 3989 2620
rect 4692 2208 5012 3232
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 10314 16896 10634 17456
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 10731 17236 10797 17237
rect 10731 17172 10732 17236
rect 10796 17172 10797 17236
rect 10731 17171 10797 17172
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 9443 16556 9509 16557
rect 9443 16492 9444 16556
rect 9508 16492 9509 16556
rect 9443 16491 9509 16492
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 7787 15604 7853 15605
rect 7787 15540 7788 15604
rect 7852 15540 7853 15604
rect 7787 15539 7853 15540
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 7790 3773 7850 15539
rect 8440 15264 8760 16288
rect 9259 16284 9325 16285
rect 9259 16220 9260 16284
rect 9324 16220 9325 16284
rect 9259 16219 9325 16220
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 9262 12205 9322 16219
rect 9259 12204 9325 12205
rect 9259 12140 9260 12204
rect 9324 12140 9325 12204
rect 9259 12139 9325 12140
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 9446 9621 9506 16491
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10179 15332 10245 15333
rect 10179 15268 10180 15332
rect 10244 15268 10245 15332
rect 10179 15267 10245 15268
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 9995 4860 10061 4861
rect 9995 4796 9996 4860
rect 10060 4796 10061 4860
rect 9995 4795 10061 4796
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 7787 3772 7853 3773
rect 7787 3708 7788 3772
rect 7852 3708 7853 3772
rect 7787 3707 7853 3708
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2128 6886 2688
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 9998 2277 10058 4795
rect 10182 2957 10242 15267
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10179 2956 10245 2957
rect 10179 2892 10180 2956
rect 10244 2892 10245 2956
rect 10179 2891 10245 2892
rect 10314 2752 10634 3776
rect 10734 3093 10794 17171
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12019 15876 12085 15877
rect 12019 15812 12020 15876
rect 12084 15812 12085 15876
rect 12019 15811 12085 15812
rect 11099 15060 11165 15061
rect 11099 14996 11100 15060
rect 11164 14996 11165 15060
rect 11099 14995 11165 14996
rect 11102 10573 11162 14995
rect 11099 10572 11165 10573
rect 11099 10508 11100 10572
rect 11164 10508 11165 10572
rect 11099 10507 11165 10508
rect 12022 10029 12082 15811
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12019 10028 12085 10029
rect 12019 9964 12020 10028
rect 12084 9964 12085 10028
rect 12019 9963 12085 9964
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14779 16556 14845 16557
rect 14779 16492 14780 16556
rect 14844 16492 14845 16556
rect 14779 16491 14845 16492
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 12571 9620 12637 9621
rect 12571 9556 12572 9620
rect 12636 9556 12637 9620
rect 12571 9555 12637 9556
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12574 8397 12634 9555
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 12571 8396 12637 8397
rect 12571 8332 12572 8396
rect 12636 8332 12637 8396
rect 12571 8331 12637 8332
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12574 3773 12634 8331
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14782 4861 14842 16491
rect 14963 15876 15029 15877
rect 14963 15812 14964 15876
rect 15028 15812 15029 15876
rect 14963 15811 15029 15812
rect 14779 4860 14845 4861
rect 14779 4796 14780 4860
rect 14844 4796 14845 4860
rect 14779 4795 14845 4796
rect 14966 4045 15026 15811
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 12571 3772 12637 3773
rect 12571 3708 12572 3772
rect 12636 3708 12637 3772
rect 12571 3707 12637 3708
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 10731 3092 10797 3093
rect 10731 3028 10732 3092
rect 10796 3028 10797 3092
rect 10731 3027 10797 3028
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 9995 2276 10061 2277
rect 9995 2212 9996 2276
rect 10060 2212 10061 2276
rect 9995 2211 10061 2212
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2128 10634 2688
rect 12188 2208 12508 3232
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform -1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 7360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 5520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 3220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform -1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform -1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 12512 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_A
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform -1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 10120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14168 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 13984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_153 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_84
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_128
timestamp 1649977179
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_101
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_152
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1649977179
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_150
timestamp 1649977179
transform 1 0 14904 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_67
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_14
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_61
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_118
timestamp 1649977179
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_10
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_147
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_144
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_129
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1649977179
transform 1 0 14260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_34
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_10
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_22
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_122
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_76
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_103
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_136
timestamp 1649977179
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_152
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_10
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1649977179
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_144
timestamp 1649977179
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_156
timestamp 1649977179
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_14
timestamp 1649977179
transform 1 0 2392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_56
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_101
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_102
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_158
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_46
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_150
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_10
timestamp 1649977179
transform 1 0 2024 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_98
timestamp 1649977179
transform 1 0 10120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_132
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_11
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_19
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_102
timestamp 1649977179
transform 1 0 10488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_106
timestamp 1649977179
transform 1 0 10856 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_158
timestamp 1649977179
transform 1 0 15640 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_21
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_44
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_98
timestamp 1649977179
transform 1 0 10120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_128
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_25
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1649977179
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_31
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_143
timestamp 1649977179
transform 1 0 14260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_35
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_95
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_107
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform -1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform -1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform -1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform -1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1649977179
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 4416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform -1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform -1 0 3036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 2852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform -1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform -1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform -1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform -1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform -1 0 9660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform -1 0 5520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform -1 0 5888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform -1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform -1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform -1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform -1 0 9292 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform -1 0 13248 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform -1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 14352 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5336 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5704 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8740 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6992 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5796 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13432 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12696 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8924 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7268 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11500 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6164 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5520 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3864 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13248 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6164 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12696 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7912 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7912 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8556 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10212 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9844 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11316 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10856 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14720 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8924 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13800 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13892 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3588 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13984 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13064 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform 1 0 15088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 590 592
<< labels >>
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 16400 2048 17200 2168 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 5 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 6 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 7 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 8 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 9 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 10 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 11 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 12 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 13 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 14 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 15 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 16 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 17 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 18 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 19 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 20 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 21 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 22 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 23 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 24 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 25 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 26 nsew signal tristate
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 27 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 28 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 29 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 30 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 31 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 32 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 33 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 34 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 35 nsew signal tristate
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 36 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 37 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 38 nsew signal tristate
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 39 nsew signal tristate
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 40 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 41 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 42 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 43 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 44 nsew signal tristate
flabel metal2 s 8758 19200 8814 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 45 nsew signal input
flabel metal2 s 12438 19200 12494 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 46 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 47 nsew signal input
flabel metal2 s 13174 19200 13230 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 48 nsew signal input
flabel metal2 s 13542 19200 13598 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 49 nsew signal input
flabel metal2 s 13910 19200 13966 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 50 nsew signal input
flabel metal2 s 14278 19200 14334 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 51 nsew signal input
flabel metal2 s 14646 19200 14702 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 52 nsew signal input
flabel metal2 s 15014 19200 15070 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 53 nsew signal input
flabel metal2 s 15382 19200 15438 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 54 nsew signal input
flabel metal2 s 15750 19200 15806 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 55 nsew signal input
flabel metal2 s 9126 19200 9182 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 56 nsew signal input
flabel metal2 s 9494 19200 9550 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 57 nsew signal input
flabel metal2 s 9862 19200 9918 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 58 nsew signal input
flabel metal2 s 10230 19200 10286 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 59 nsew signal input
flabel metal2 s 10598 19200 10654 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 60 nsew signal input
flabel metal2 s 10966 19200 11022 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 61 nsew signal input
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 62 nsew signal input
flabel metal2 s 11702 19200 11758 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 63 nsew signal input
flabel metal2 s 12070 19200 12126 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 64 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 65 nsew signal tristate
flabel metal2 s 5078 19200 5134 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 66 nsew signal tristate
flabel metal2 s 5446 19200 5502 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 67 nsew signal tristate
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 68 nsew signal tristate
flabel metal2 s 6182 19200 6238 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 69 nsew signal tristate
flabel metal2 s 6550 19200 6606 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 70 nsew signal tristate
flabel metal2 s 6918 19200 6974 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 71 nsew signal tristate
flabel metal2 s 7286 19200 7342 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 72 nsew signal tristate
flabel metal2 s 7654 19200 7710 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 73 nsew signal tristate
flabel metal2 s 8022 19200 8078 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 74 nsew signal tristate
flabel metal2 s 8390 19200 8446 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 75 nsew signal tristate
flabel metal2 s 1766 19200 1822 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 76 nsew signal tristate
flabel metal2 s 2134 19200 2190 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 77 nsew signal tristate
flabel metal2 s 2502 19200 2558 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 78 nsew signal tristate
flabel metal2 s 2870 19200 2926 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 79 nsew signal tristate
flabel metal2 s 3238 19200 3294 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 80 nsew signal tristate
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 81 nsew signal tristate
flabel metal2 s 3974 19200 4030 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 82 nsew signal tristate
flabel metal2 s 4342 19200 4398 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 83 nsew signal tristate
flabel metal2 s 4710 19200 4766 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 84 nsew signal tristate
flabel metal3 s 16400 9936 17200 10056 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
flabel metal3 s 16400 13880 17200 14000 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
flabel metal3 s 16400 17824 17200 17944 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_grid_pin_16_
port 88 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 left_grid_pin_17_
port 89 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 left_grid_pin_18_
port 90 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 left_grid_pin_19_
port 91 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 left_grid_pin_20_
port 92 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 left_grid_pin_21_
port 93 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 left_grid_pin_22_
port 94 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 left_grid_pin_23_
port 95 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 left_grid_pin_24_
port 96 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 left_grid_pin_25_
port 97 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 left_grid_pin_26_
port 98 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 left_grid_pin_27_
port 99 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 left_grid_pin_28_
port 100 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 left_grid_pin_29_
port 101 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 left_grid_pin_30_
port 102 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 left_grid_pin_31_
port 103 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_0_
port 104 nsew signal input
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_1_lower
port 105 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_1_upper
port 106 nsew signal tristate
flabel metal2 s 16118 19200 16174 20000 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 107 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 108 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 prog_clk_0_W_in
port 109 nsew signal input
flabel metal3 s 16400 5992 17200 6112 0 FreeSans 480 0 0 0 right_grid_pin_0_
port 110 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
