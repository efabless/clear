//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Nov 24 18:04:19 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- Verilog module for fpga_top -----
module fpga_top(prog_clk,
                Test_en,
                IO_ISOL_N,
                clk,
                gfpga_pad_EMBEDDED_IO_HD_SOC_IN,
                gfpga_pad_EMBEDDED_IO_HD_SOC_OUT,
                gfpga_pad_EMBEDDED_IO_HD_SOC_DIR,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GLOBAL PORTS -----
input [0:0] IO_ISOL_N;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIN PORTS -----
input [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
//----- GPOUT PORTS -----
output [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
//----- GPOUT PORTS -----
output [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__0_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:19] cbx_1__0__0_chanx_left_out;
wire [0:19] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:19] cbx_1__0__1_chanx_left_out;
wire [0:19] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__2_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:19] cbx_1__0__2_chanx_left_out;
wire [0:19] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__3_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:19] cbx_1__0__3_chanx_left_out;
wire [0:19] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__4_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:19] cbx_1__0__4_chanx_left_out;
wire [0:19] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__5_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:19] cbx_1__0__5_chanx_left_out;
wire [0:19] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__0__6_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__6_ccff_tail;
wire [0:19] cbx_1__0__6_chanx_left_out;
wire [0:19] cbx_1__0__6_chanx_right_out;
wire [0:0] cbx_1__0__7_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_10_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_12_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_14_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_16_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_2_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_4_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_6_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_8_;
wire [0:0] cbx_1__0__7_ccff_tail;
wire [0:19] cbx_1__0__7_chanx_left_out;
wire [0:19] cbx_1__0__7_chanx_right_out;
wire [0:0] cbx_1__1__0_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__0_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:19] cbx_1__1__0_chanx_left_out;
wire [0:19] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__10_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__10_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__10_ccff_tail;
wire [0:19] cbx_1__1__10_chanx_left_out;
wire [0:19] cbx_1__1__10_chanx_right_out;
wire [0:0] cbx_1__1__11_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__11_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__11_ccff_tail;
wire [0:19] cbx_1__1__11_chanx_left_out;
wire [0:19] cbx_1__1__11_chanx_right_out;
wire [0:0] cbx_1__1__12_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__12_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__12_ccff_tail;
wire [0:19] cbx_1__1__12_chanx_left_out;
wire [0:19] cbx_1__1__12_chanx_right_out;
wire [0:0] cbx_1__1__13_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__13_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__13_ccff_tail;
wire [0:19] cbx_1__1__13_chanx_left_out;
wire [0:19] cbx_1__1__13_chanx_right_out;
wire [0:0] cbx_1__1__14_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__14_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__14_ccff_tail;
wire [0:19] cbx_1__1__14_chanx_left_out;
wire [0:19] cbx_1__1__14_chanx_right_out;
wire [0:0] cbx_1__1__15_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__15_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__15_ccff_tail;
wire [0:19] cbx_1__1__15_chanx_left_out;
wire [0:19] cbx_1__1__15_chanx_right_out;
wire [0:0] cbx_1__1__16_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__16_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__16_ccff_tail;
wire [0:19] cbx_1__1__16_chanx_left_out;
wire [0:19] cbx_1__1__16_chanx_right_out;
wire [0:0] cbx_1__1__17_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__17_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__17_ccff_tail;
wire [0:19] cbx_1__1__17_chanx_left_out;
wire [0:19] cbx_1__1__17_chanx_right_out;
wire [0:0] cbx_1__1__18_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__18_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__18_ccff_tail;
wire [0:19] cbx_1__1__18_chanx_left_out;
wire [0:19] cbx_1__1__18_chanx_right_out;
wire [0:0] cbx_1__1__19_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__19_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__19_ccff_tail;
wire [0:19] cbx_1__1__19_chanx_left_out;
wire [0:19] cbx_1__1__19_chanx_right_out;
wire [0:0] cbx_1__1__1_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__1_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:19] cbx_1__1__1_chanx_left_out;
wire [0:19] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__1__20_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__20_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__20_ccff_tail;
wire [0:19] cbx_1__1__20_chanx_left_out;
wire [0:19] cbx_1__1__20_chanx_right_out;
wire [0:0] cbx_1__1__21_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__21_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__21_ccff_tail;
wire [0:19] cbx_1__1__21_chanx_left_out;
wire [0:19] cbx_1__1__21_chanx_right_out;
wire [0:0] cbx_1__1__22_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__22_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__22_ccff_tail;
wire [0:19] cbx_1__1__22_chanx_left_out;
wire [0:19] cbx_1__1__22_chanx_right_out;
wire [0:0] cbx_1__1__23_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__23_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__23_ccff_tail;
wire [0:19] cbx_1__1__23_chanx_left_out;
wire [0:19] cbx_1__1__23_chanx_right_out;
wire [0:0] cbx_1__1__24_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__24_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__24_ccff_tail;
wire [0:19] cbx_1__1__24_chanx_left_out;
wire [0:19] cbx_1__1__24_chanx_right_out;
wire [0:0] cbx_1__1__25_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__25_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__25_ccff_tail;
wire [0:19] cbx_1__1__25_chanx_left_out;
wire [0:19] cbx_1__1__25_chanx_right_out;
wire [0:0] cbx_1__1__26_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__26_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__26_ccff_tail;
wire [0:19] cbx_1__1__26_chanx_left_out;
wire [0:19] cbx_1__1__26_chanx_right_out;
wire [0:0] cbx_1__1__27_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__27_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__27_ccff_tail;
wire [0:19] cbx_1__1__27_chanx_left_out;
wire [0:19] cbx_1__1__27_chanx_right_out;
wire [0:0] cbx_1__1__28_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__28_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__28_ccff_tail;
wire [0:19] cbx_1__1__28_chanx_left_out;
wire [0:19] cbx_1__1__28_chanx_right_out;
wire [0:0] cbx_1__1__29_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__29_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__29_ccff_tail;
wire [0:19] cbx_1__1__29_chanx_left_out;
wire [0:19] cbx_1__1__29_chanx_right_out;
wire [0:0] cbx_1__1__2_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__2_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__2_ccff_tail;
wire [0:19] cbx_1__1__2_chanx_left_out;
wire [0:19] cbx_1__1__2_chanx_right_out;
wire [0:0] cbx_1__1__30_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__30_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__30_ccff_tail;
wire [0:19] cbx_1__1__30_chanx_left_out;
wire [0:19] cbx_1__1__30_chanx_right_out;
wire [0:0] cbx_1__1__31_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__31_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__31_ccff_tail;
wire [0:19] cbx_1__1__31_chanx_left_out;
wire [0:19] cbx_1__1__31_chanx_right_out;
wire [0:0] cbx_1__1__32_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__32_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__32_ccff_tail;
wire [0:19] cbx_1__1__32_chanx_left_out;
wire [0:19] cbx_1__1__32_chanx_right_out;
wire [0:0] cbx_1__1__33_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__33_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__33_ccff_tail;
wire [0:19] cbx_1__1__33_chanx_left_out;
wire [0:19] cbx_1__1__33_chanx_right_out;
wire [0:0] cbx_1__1__34_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__34_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__34_ccff_tail;
wire [0:19] cbx_1__1__34_chanx_left_out;
wire [0:19] cbx_1__1__34_chanx_right_out;
wire [0:0] cbx_1__1__35_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__35_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__35_ccff_tail;
wire [0:19] cbx_1__1__35_chanx_left_out;
wire [0:19] cbx_1__1__35_chanx_right_out;
wire [0:0] cbx_1__1__36_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__36_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__36_ccff_tail;
wire [0:19] cbx_1__1__36_chanx_left_out;
wire [0:19] cbx_1__1__36_chanx_right_out;
wire [0:0] cbx_1__1__37_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__37_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__37_ccff_tail;
wire [0:19] cbx_1__1__37_chanx_left_out;
wire [0:19] cbx_1__1__37_chanx_right_out;
wire [0:0] cbx_1__1__38_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__38_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__38_ccff_tail;
wire [0:19] cbx_1__1__38_chanx_left_out;
wire [0:19] cbx_1__1__38_chanx_right_out;
wire [0:0] cbx_1__1__39_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__39_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__39_ccff_tail;
wire [0:19] cbx_1__1__39_chanx_left_out;
wire [0:19] cbx_1__1__39_chanx_right_out;
wire [0:0] cbx_1__1__3_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__3_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__3_ccff_tail;
wire [0:19] cbx_1__1__3_chanx_left_out;
wire [0:19] cbx_1__1__3_chanx_right_out;
wire [0:0] cbx_1__1__40_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__40_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__40_ccff_tail;
wire [0:19] cbx_1__1__40_chanx_left_out;
wire [0:19] cbx_1__1__40_chanx_right_out;
wire [0:0] cbx_1__1__41_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__41_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__41_ccff_tail;
wire [0:19] cbx_1__1__41_chanx_left_out;
wire [0:19] cbx_1__1__41_chanx_right_out;
wire [0:0] cbx_1__1__42_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__42_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__42_ccff_tail;
wire [0:19] cbx_1__1__42_chanx_left_out;
wire [0:19] cbx_1__1__42_chanx_right_out;
wire [0:0] cbx_1__1__43_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__43_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__43_ccff_tail;
wire [0:19] cbx_1__1__43_chanx_left_out;
wire [0:19] cbx_1__1__43_chanx_right_out;
wire [0:0] cbx_1__1__44_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__44_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__44_ccff_tail;
wire [0:19] cbx_1__1__44_chanx_left_out;
wire [0:19] cbx_1__1__44_chanx_right_out;
wire [0:0] cbx_1__1__45_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__45_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__45_ccff_tail;
wire [0:19] cbx_1__1__45_chanx_left_out;
wire [0:19] cbx_1__1__45_chanx_right_out;
wire [0:0] cbx_1__1__46_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__46_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__46_ccff_tail;
wire [0:19] cbx_1__1__46_chanx_left_out;
wire [0:19] cbx_1__1__46_chanx_right_out;
wire [0:0] cbx_1__1__47_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__47_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__47_ccff_tail;
wire [0:19] cbx_1__1__47_chanx_left_out;
wire [0:19] cbx_1__1__47_chanx_right_out;
wire [0:0] cbx_1__1__48_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__48_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__48_ccff_tail;
wire [0:19] cbx_1__1__48_chanx_left_out;
wire [0:19] cbx_1__1__48_chanx_right_out;
wire [0:0] cbx_1__1__49_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__49_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__49_ccff_tail;
wire [0:19] cbx_1__1__49_chanx_left_out;
wire [0:19] cbx_1__1__49_chanx_right_out;
wire [0:0] cbx_1__1__4_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__4_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__4_ccff_tail;
wire [0:19] cbx_1__1__4_chanx_left_out;
wire [0:19] cbx_1__1__4_chanx_right_out;
wire [0:0] cbx_1__1__50_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__50_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__50_ccff_tail;
wire [0:19] cbx_1__1__50_chanx_left_out;
wire [0:19] cbx_1__1__50_chanx_right_out;
wire [0:0] cbx_1__1__51_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__51_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__51_ccff_tail;
wire [0:19] cbx_1__1__51_chanx_left_out;
wire [0:19] cbx_1__1__51_chanx_right_out;
wire [0:0] cbx_1__1__52_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__52_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__52_ccff_tail;
wire [0:19] cbx_1__1__52_chanx_left_out;
wire [0:19] cbx_1__1__52_chanx_right_out;
wire [0:0] cbx_1__1__53_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__53_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__53_ccff_tail;
wire [0:19] cbx_1__1__53_chanx_left_out;
wire [0:19] cbx_1__1__53_chanx_right_out;
wire [0:0] cbx_1__1__54_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__54_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__54_ccff_tail;
wire [0:19] cbx_1__1__54_chanx_left_out;
wire [0:19] cbx_1__1__54_chanx_right_out;
wire [0:0] cbx_1__1__55_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__55_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__55_ccff_tail;
wire [0:19] cbx_1__1__55_chanx_left_out;
wire [0:19] cbx_1__1__55_chanx_right_out;
wire [0:0] cbx_1__1__5_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__5_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__5_ccff_tail;
wire [0:19] cbx_1__1__5_chanx_left_out;
wire [0:19] cbx_1__1__5_chanx_right_out;
wire [0:0] cbx_1__1__6_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__6_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__6_ccff_tail;
wire [0:19] cbx_1__1__6_chanx_left_out;
wire [0:19] cbx_1__1__6_chanx_right_out;
wire [0:0] cbx_1__1__7_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__7_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__7_ccff_tail;
wire [0:19] cbx_1__1__7_chanx_left_out;
wire [0:19] cbx_1__1__7_chanx_right_out;
wire [0:0] cbx_1__1__8_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__8_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__8_ccff_tail;
wire [0:19] cbx_1__1__8_chanx_left_out;
wire [0:19] cbx_1__1__8_chanx_right_out;
wire [0:0] cbx_1__1__9_bottom_grid_pin_0_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_10_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_11_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_12_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_13_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_14_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_15_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_1_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_2_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_3_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_4_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_5_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_6_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_7_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_8_;
wire [0:0] cbx_1__1__9_bottom_grid_pin_9_;
wire [0:0] cbx_1__1__9_ccff_tail;
wire [0:19] cbx_1__1__9_chanx_left_out;
wire [0:19] cbx_1__1__9_chanx_right_out;
wire [0:0] cbx_1__8__0_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__0_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__0_ccff_tail;
wire [0:19] cbx_1__8__0_chanx_left_out;
wire [0:19] cbx_1__8__0_chanx_right_out;
wire [0:0] cbx_1__8__0_top_grid_pin_0_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__1_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__1_ccff_tail;
wire [0:19] cbx_1__8__1_chanx_left_out;
wire [0:19] cbx_1__8__1_chanx_right_out;
wire [0:0] cbx_1__8__1_top_grid_pin_0_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__2_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__2_ccff_tail;
wire [0:19] cbx_1__8__2_chanx_left_out;
wire [0:19] cbx_1__8__2_chanx_right_out;
wire [0:0] cbx_1__8__2_top_grid_pin_0_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__3_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__3_ccff_tail;
wire [0:19] cbx_1__8__3_chanx_left_out;
wire [0:19] cbx_1__8__3_chanx_right_out;
wire [0:0] cbx_1__8__3_top_grid_pin_0_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__4_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__4_ccff_tail;
wire [0:19] cbx_1__8__4_chanx_left_out;
wire [0:19] cbx_1__8__4_chanx_right_out;
wire [0:0] cbx_1__8__4_top_grid_pin_0_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__5_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__5_ccff_tail;
wire [0:19] cbx_1__8__5_chanx_left_out;
wire [0:19] cbx_1__8__5_chanx_right_out;
wire [0:0] cbx_1__8__5_top_grid_pin_0_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__6_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__6_ccff_tail;
wire [0:19] cbx_1__8__6_chanx_left_out;
wire [0:19] cbx_1__8__6_chanx_right_out;
wire [0:0] cbx_1__8__6_top_grid_pin_0_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_0_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_10_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_11_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_12_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_13_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_14_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_15_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_1_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_2_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_3_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_4_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_5_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_6_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_7_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_8_;
wire [0:0] cbx_1__8__7_bottom_grid_pin_9_;
wire [0:0] cbx_1__8__7_ccff_tail;
wire [0:19] cbx_1__8__7_chanx_left_out;
wire [0:19] cbx_1__8__7_chanx_right_out;
wire [0:0] cbx_1__8__7_top_grid_pin_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:19] cby_0__1__0_chany_bottom_out;
wire [0:19] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_pin_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:19] cby_0__1__1_chany_bottom_out;
wire [0:19] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_pin_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:19] cby_0__1__2_chany_bottom_out;
wire [0:19] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_pin_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:19] cby_0__1__3_chany_bottom_out;
wire [0:19] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_pin_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:19] cby_0__1__4_chany_bottom_out;
wire [0:19] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_pin_0_;
wire [0:0] cby_0__1__5_ccff_tail;
wire [0:19] cby_0__1__5_chany_bottom_out;
wire [0:19] cby_0__1__5_chany_top_out;
wire [0:0] cby_0__1__5_left_grid_pin_0_;
wire [0:0] cby_0__1__6_ccff_tail;
wire [0:19] cby_0__1__6_chany_bottom_out;
wire [0:19] cby_0__1__6_chany_top_out;
wire [0:0] cby_0__1__6_left_grid_pin_0_;
wire [0:0] cby_0__1__7_ccff_tail;
wire [0:19] cby_0__1__7_chany_bottom_out;
wire [0:19] cby_0__1__7_chany_top_out;
wire [0:0] cby_0__1__7_left_grid_pin_0_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:19] cby_1__1__0_chany_bottom_out;
wire [0:19] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_pin_16_;
wire [0:0] cby_1__1__0_left_grid_pin_17_;
wire [0:0] cby_1__1__0_left_grid_pin_18_;
wire [0:0] cby_1__1__0_left_grid_pin_19_;
wire [0:0] cby_1__1__0_left_grid_pin_20_;
wire [0:0] cby_1__1__0_left_grid_pin_21_;
wire [0:0] cby_1__1__0_left_grid_pin_22_;
wire [0:0] cby_1__1__0_left_grid_pin_23_;
wire [0:0] cby_1__1__0_left_grid_pin_24_;
wire [0:0] cby_1__1__0_left_grid_pin_25_;
wire [0:0] cby_1__1__0_left_grid_pin_26_;
wire [0:0] cby_1__1__0_left_grid_pin_27_;
wire [0:0] cby_1__1__0_left_grid_pin_28_;
wire [0:0] cby_1__1__0_left_grid_pin_29_;
wire [0:0] cby_1__1__0_left_grid_pin_30_;
wire [0:0] cby_1__1__0_left_grid_pin_31_;
wire [0:0] cby_1__1__10_ccff_tail;
wire [0:19] cby_1__1__10_chany_bottom_out;
wire [0:19] cby_1__1__10_chany_top_out;
wire [0:0] cby_1__1__10_left_grid_pin_16_;
wire [0:0] cby_1__1__10_left_grid_pin_17_;
wire [0:0] cby_1__1__10_left_grid_pin_18_;
wire [0:0] cby_1__1__10_left_grid_pin_19_;
wire [0:0] cby_1__1__10_left_grid_pin_20_;
wire [0:0] cby_1__1__10_left_grid_pin_21_;
wire [0:0] cby_1__1__10_left_grid_pin_22_;
wire [0:0] cby_1__1__10_left_grid_pin_23_;
wire [0:0] cby_1__1__10_left_grid_pin_24_;
wire [0:0] cby_1__1__10_left_grid_pin_25_;
wire [0:0] cby_1__1__10_left_grid_pin_26_;
wire [0:0] cby_1__1__10_left_grid_pin_27_;
wire [0:0] cby_1__1__10_left_grid_pin_28_;
wire [0:0] cby_1__1__10_left_grid_pin_29_;
wire [0:0] cby_1__1__10_left_grid_pin_30_;
wire [0:0] cby_1__1__10_left_grid_pin_31_;
wire [0:0] cby_1__1__11_ccff_tail;
wire [0:19] cby_1__1__11_chany_bottom_out;
wire [0:19] cby_1__1__11_chany_top_out;
wire [0:0] cby_1__1__11_left_grid_pin_16_;
wire [0:0] cby_1__1__11_left_grid_pin_17_;
wire [0:0] cby_1__1__11_left_grid_pin_18_;
wire [0:0] cby_1__1__11_left_grid_pin_19_;
wire [0:0] cby_1__1__11_left_grid_pin_20_;
wire [0:0] cby_1__1__11_left_grid_pin_21_;
wire [0:0] cby_1__1__11_left_grid_pin_22_;
wire [0:0] cby_1__1__11_left_grid_pin_23_;
wire [0:0] cby_1__1__11_left_grid_pin_24_;
wire [0:0] cby_1__1__11_left_grid_pin_25_;
wire [0:0] cby_1__1__11_left_grid_pin_26_;
wire [0:0] cby_1__1__11_left_grid_pin_27_;
wire [0:0] cby_1__1__11_left_grid_pin_28_;
wire [0:0] cby_1__1__11_left_grid_pin_29_;
wire [0:0] cby_1__1__11_left_grid_pin_30_;
wire [0:0] cby_1__1__11_left_grid_pin_31_;
wire [0:0] cby_1__1__12_ccff_tail;
wire [0:19] cby_1__1__12_chany_bottom_out;
wire [0:19] cby_1__1__12_chany_top_out;
wire [0:0] cby_1__1__12_left_grid_pin_16_;
wire [0:0] cby_1__1__12_left_grid_pin_17_;
wire [0:0] cby_1__1__12_left_grid_pin_18_;
wire [0:0] cby_1__1__12_left_grid_pin_19_;
wire [0:0] cby_1__1__12_left_grid_pin_20_;
wire [0:0] cby_1__1__12_left_grid_pin_21_;
wire [0:0] cby_1__1__12_left_grid_pin_22_;
wire [0:0] cby_1__1__12_left_grid_pin_23_;
wire [0:0] cby_1__1__12_left_grid_pin_24_;
wire [0:0] cby_1__1__12_left_grid_pin_25_;
wire [0:0] cby_1__1__12_left_grid_pin_26_;
wire [0:0] cby_1__1__12_left_grid_pin_27_;
wire [0:0] cby_1__1__12_left_grid_pin_28_;
wire [0:0] cby_1__1__12_left_grid_pin_29_;
wire [0:0] cby_1__1__12_left_grid_pin_30_;
wire [0:0] cby_1__1__12_left_grid_pin_31_;
wire [0:0] cby_1__1__13_ccff_tail;
wire [0:19] cby_1__1__13_chany_bottom_out;
wire [0:19] cby_1__1__13_chany_top_out;
wire [0:0] cby_1__1__13_left_grid_pin_16_;
wire [0:0] cby_1__1__13_left_grid_pin_17_;
wire [0:0] cby_1__1__13_left_grid_pin_18_;
wire [0:0] cby_1__1__13_left_grid_pin_19_;
wire [0:0] cby_1__1__13_left_grid_pin_20_;
wire [0:0] cby_1__1__13_left_grid_pin_21_;
wire [0:0] cby_1__1__13_left_grid_pin_22_;
wire [0:0] cby_1__1__13_left_grid_pin_23_;
wire [0:0] cby_1__1__13_left_grid_pin_24_;
wire [0:0] cby_1__1__13_left_grid_pin_25_;
wire [0:0] cby_1__1__13_left_grid_pin_26_;
wire [0:0] cby_1__1__13_left_grid_pin_27_;
wire [0:0] cby_1__1__13_left_grid_pin_28_;
wire [0:0] cby_1__1__13_left_grid_pin_29_;
wire [0:0] cby_1__1__13_left_grid_pin_30_;
wire [0:0] cby_1__1__13_left_grid_pin_31_;
wire [0:0] cby_1__1__14_ccff_tail;
wire [0:19] cby_1__1__14_chany_bottom_out;
wire [0:19] cby_1__1__14_chany_top_out;
wire [0:0] cby_1__1__14_left_grid_pin_16_;
wire [0:0] cby_1__1__14_left_grid_pin_17_;
wire [0:0] cby_1__1__14_left_grid_pin_18_;
wire [0:0] cby_1__1__14_left_grid_pin_19_;
wire [0:0] cby_1__1__14_left_grid_pin_20_;
wire [0:0] cby_1__1__14_left_grid_pin_21_;
wire [0:0] cby_1__1__14_left_grid_pin_22_;
wire [0:0] cby_1__1__14_left_grid_pin_23_;
wire [0:0] cby_1__1__14_left_grid_pin_24_;
wire [0:0] cby_1__1__14_left_grid_pin_25_;
wire [0:0] cby_1__1__14_left_grid_pin_26_;
wire [0:0] cby_1__1__14_left_grid_pin_27_;
wire [0:0] cby_1__1__14_left_grid_pin_28_;
wire [0:0] cby_1__1__14_left_grid_pin_29_;
wire [0:0] cby_1__1__14_left_grid_pin_30_;
wire [0:0] cby_1__1__14_left_grid_pin_31_;
wire [0:0] cby_1__1__15_ccff_tail;
wire [0:19] cby_1__1__15_chany_bottom_out;
wire [0:19] cby_1__1__15_chany_top_out;
wire [0:0] cby_1__1__15_left_grid_pin_16_;
wire [0:0] cby_1__1__15_left_grid_pin_17_;
wire [0:0] cby_1__1__15_left_grid_pin_18_;
wire [0:0] cby_1__1__15_left_grid_pin_19_;
wire [0:0] cby_1__1__15_left_grid_pin_20_;
wire [0:0] cby_1__1__15_left_grid_pin_21_;
wire [0:0] cby_1__1__15_left_grid_pin_22_;
wire [0:0] cby_1__1__15_left_grid_pin_23_;
wire [0:0] cby_1__1__15_left_grid_pin_24_;
wire [0:0] cby_1__1__15_left_grid_pin_25_;
wire [0:0] cby_1__1__15_left_grid_pin_26_;
wire [0:0] cby_1__1__15_left_grid_pin_27_;
wire [0:0] cby_1__1__15_left_grid_pin_28_;
wire [0:0] cby_1__1__15_left_grid_pin_29_;
wire [0:0] cby_1__1__15_left_grid_pin_30_;
wire [0:0] cby_1__1__15_left_grid_pin_31_;
wire [0:0] cby_1__1__16_ccff_tail;
wire [0:19] cby_1__1__16_chany_bottom_out;
wire [0:19] cby_1__1__16_chany_top_out;
wire [0:0] cby_1__1__16_left_grid_pin_16_;
wire [0:0] cby_1__1__16_left_grid_pin_17_;
wire [0:0] cby_1__1__16_left_grid_pin_18_;
wire [0:0] cby_1__1__16_left_grid_pin_19_;
wire [0:0] cby_1__1__16_left_grid_pin_20_;
wire [0:0] cby_1__1__16_left_grid_pin_21_;
wire [0:0] cby_1__1__16_left_grid_pin_22_;
wire [0:0] cby_1__1__16_left_grid_pin_23_;
wire [0:0] cby_1__1__16_left_grid_pin_24_;
wire [0:0] cby_1__1__16_left_grid_pin_25_;
wire [0:0] cby_1__1__16_left_grid_pin_26_;
wire [0:0] cby_1__1__16_left_grid_pin_27_;
wire [0:0] cby_1__1__16_left_grid_pin_28_;
wire [0:0] cby_1__1__16_left_grid_pin_29_;
wire [0:0] cby_1__1__16_left_grid_pin_30_;
wire [0:0] cby_1__1__16_left_grid_pin_31_;
wire [0:0] cby_1__1__17_ccff_tail;
wire [0:19] cby_1__1__17_chany_bottom_out;
wire [0:19] cby_1__1__17_chany_top_out;
wire [0:0] cby_1__1__17_left_grid_pin_16_;
wire [0:0] cby_1__1__17_left_grid_pin_17_;
wire [0:0] cby_1__1__17_left_grid_pin_18_;
wire [0:0] cby_1__1__17_left_grid_pin_19_;
wire [0:0] cby_1__1__17_left_grid_pin_20_;
wire [0:0] cby_1__1__17_left_grid_pin_21_;
wire [0:0] cby_1__1__17_left_grid_pin_22_;
wire [0:0] cby_1__1__17_left_grid_pin_23_;
wire [0:0] cby_1__1__17_left_grid_pin_24_;
wire [0:0] cby_1__1__17_left_grid_pin_25_;
wire [0:0] cby_1__1__17_left_grid_pin_26_;
wire [0:0] cby_1__1__17_left_grid_pin_27_;
wire [0:0] cby_1__1__17_left_grid_pin_28_;
wire [0:0] cby_1__1__17_left_grid_pin_29_;
wire [0:0] cby_1__1__17_left_grid_pin_30_;
wire [0:0] cby_1__1__17_left_grid_pin_31_;
wire [0:0] cby_1__1__18_ccff_tail;
wire [0:19] cby_1__1__18_chany_bottom_out;
wire [0:19] cby_1__1__18_chany_top_out;
wire [0:0] cby_1__1__18_left_grid_pin_16_;
wire [0:0] cby_1__1__18_left_grid_pin_17_;
wire [0:0] cby_1__1__18_left_grid_pin_18_;
wire [0:0] cby_1__1__18_left_grid_pin_19_;
wire [0:0] cby_1__1__18_left_grid_pin_20_;
wire [0:0] cby_1__1__18_left_grid_pin_21_;
wire [0:0] cby_1__1__18_left_grid_pin_22_;
wire [0:0] cby_1__1__18_left_grid_pin_23_;
wire [0:0] cby_1__1__18_left_grid_pin_24_;
wire [0:0] cby_1__1__18_left_grid_pin_25_;
wire [0:0] cby_1__1__18_left_grid_pin_26_;
wire [0:0] cby_1__1__18_left_grid_pin_27_;
wire [0:0] cby_1__1__18_left_grid_pin_28_;
wire [0:0] cby_1__1__18_left_grid_pin_29_;
wire [0:0] cby_1__1__18_left_grid_pin_30_;
wire [0:0] cby_1__1__18_left_grid_pin_31_;
wire [0:0] cby_1__1__19_ccff_tail;
wire [0:19] cby_1__1__19_chany_bottom_out;
wire [0:19] cby_1__1__19_chany_top_out;
wire [0:0] cby_1__1__19_left_grid_pin_16_;
wire [0:0] cby_1__1__19_left_grid_pin_17_;
wire [0:0] cby_1__1__19_left_grid_pin_18_;
wire [0:0] cby_1__1__19_left_grid_pin_19_;
wire [0:0] cby_1__1__19_left_grid_pin_20_;
wire [0:0] cby_1__1__19_left_grid_pin_21_;
wire [0:0] cby_1__1__19_left_grid_pin_22_;
wire [0:0] cby_1__1__19_left_grid_pin_23_;
wire [0:0] cby_1__1__19_left_grid_pin_24_;
wire [0:0] cby_1__1__19_left_grid_pin_25_;
wire [0:0] cby_1__1__19_left_grid_pin_26_;
wire [0:0] cby_1__1__19_left_grid_pin_27_;
wire [0:0] cby_1__1__19_left_grid_pin_28_;
wire [0:0] cby_1__1__19_left_grid_pin_29_;
wire [0:0] cby_1__1__19_left_grid_pin_30_;
wire [0:0] cby_1__1__19_left_grid_pin_31_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:19] cby_1__1__1_chany_bottom_out;
wire [0:19] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_pin_16_;
wire [0:0] cby_1__1__1_left_grid_pin_17_;
wire [0:0] cby_1__1__1_left_grid_pin_18_;
wire [0:0] cby_1__1__1_left_grid_pin_19_;
wire [0:0] cby_1__1__1_left_grid_pin_20_;
wire [0:0] cby_1__1__1_left_grid_pin_21_;
wire [0:0] cby_1__1__1_left_grid_pin_22_;
wire [0:0] cby_1__1__1_left_grid_pin_23_;
wire [0:0] cby_1__1__1_left_grid_pin_24_;
wire [0:0] cby_1__1__1_left_grid_pin_25_;
wire [0:0] cby_1__1__1_left_grid_pin_26_;
wire [0:0] cby_1__1__1_left_grid_pin_27_;
wire [0:0] cby_1__1__1_left_grid_pin_28_;
wire [0:0] cby_1__1__1_left_grid_pin_29_;
wire [0:0] cby_1__1__1_left_grid_pin_30_;
wire [0:0] cby_1__1__1_left_grid_pin_31_;
wire [0:0] cby_1__1__20_ccff_tail;
wire [0:19] cby_1__1__20_chany_bottom_out;
wire [0:19] cby_1__1__20_chany_top_out;
wire [0:0] cby_1__1__20_left_grid_pin_16_;
wire [0:0] cby_1__1__20_left_grid_pin_17_;
wire [0:0] cby_1__1__20_left_grid_pin_18_;
wire [0:0] cby_1__1__20_left_grid_pin_19_;
wire [0:0] cby_1__1__20_left_grid_pin_20_;
wire [0:0] cby_1__1__20_left_grid_pin_21_;
wire [0:0] cby_1__1__20_left_grid_pin_22_;
wire [0:0] cby_1__1__20_left_grid_pin_23_;
wire [0:0] cby_1__1__20_left_grid_pin_24_;
wire [0:0] cby_1__1__20_left_grid_pin_25_;
wire [0:0] cby_1__1__20_left_grid_pin_26_;
wire [0:0] cby_1__1__20_left_grid_pin_27_;
wire [0:0] cby_1__1__20_left_grid_pin_28_;
wire [0:0] cby_1__1__20_left_grid_pin_29_;
wire [0:0] cby_1__1__20_left_grid_pin_30_;
wire [0:0] cby_1__1__20_left_grid_pin_31_;
wire [0:0] cby_1__1__21_ccff_tail;
wire [0:19] cby_1__1__21_chany_bottom_out;
wire [0:19] cby_1__1__21_chany_top_out;
wire [0:0] cby_1__1__21_left_grid_pin_16_;
wire [0:0] cby_1__1__21_left_grid_pin_17_;
wire [0:0] cby_1__1__21_left_grid_pin_18_;
wire [0:0] cby_1__1__21_left_grid_pin_19_;
wire [0:0] cby_1__1__21_left_grid_pin_20_;
wire [0:0] cby_1__1__21_left_grid_pin_21_;
wire [0:0] cby_1__1__21_left_grid_pin_22_;
wire [0:0] cby_1__1__21_left_grid_pin_23_;
wire [0:0] cby_1__1__21_left_grid_pin_24_;
wire [0:0] cby_1__1__21_left_grid_pin_25_;
wire [0:0] cby_1__1__21_left_grid_pin_26_;
wire [0:0] cby_1__1__21_left_grid_pin_27_;
wire [0:0] cby_1__1__21_left_grid_pin_28_;
wire [0:0] cby_1__1__21_left_grid_pin_29_;
wire [0:0] cby_1__1__21_left_grid_pin_30_;
wire [0:0] cby_1__1__21_left_grid_pin_31_;
wire [0:0] cby_1__1__22_ccff_tail;
wire [0:19] cby_1__1__22_chany_bottom_out;
wire [0:19] cby_1__1__22_chany_top_out;
wire [0:0] cby_1__1__22_left_grid_pin_16_;
wire [0:0] cby_1__1__22_left_grid_pin_17_;
wire [0:0] cby_1__1__22_left_grid_pin_18_;
wire [0:0] cby_1__1__22_left_grid_pin_19_;
wire [0:0] cby_1__1__22_left_grid_pin_20_;
wire [0:0] cby_1__1__22_left_grid_pin_21_;
wire [0:0] cby_1__1__22_left_grid_pin_22_;
wire [0:0] cby_1__1__22_left_grid_pin_23_;
wire [0:0] cby_1__1__22_left_grid_pin_24_;
wire [0:0] cby_1__1__22_left_grid_pin_25_;
wire [0:0] cby_1__1__22_left_grid_pin_26_;
wire [0:0] cby_1__1__22_left_grid_pin_27_;
wire [0:0] cby_1__1__22_left_grid_pin_28_;
wire [0:0] cby_1__1__22_left_grid_pin_29_;
wire [0:0] cby_1__1__22_left_grid_pin_30_;
wire [0:0] cby_1__1__22_left_grid_pin_31_;
wire [0:0] cby_1__1__23_ccff_tail;
wire [0:19] cby_1__1__23_chany_bottom_out;
wire [0:19] cby_1__1__23_chany_top_out;
wire [0:0] cby_1__1__23_left_grid_pin_16_;
wire [0:0] cby_1__1__23_left_grid_pin_17_;
wire [0:0] cby_1__1__23_left_grid_pin_18_;
wire [0:0] cby_1__1__23_left_grid_pin_19_;
wire [0:0] cby_1__1__23_left_grid_pin_20_;
wire [0:0] cby_1__1__23_left_grid_pin_21_;
wire [0:0] cby_1__1__23_left_grid_pin_22_;
wire [0:0] cby_1__1__23_left_grid_pin_23_;
wire [0:0] cby_1__1__23_left_grid_pin_24_;
wire [0:0] cby_1__1__23_left_grid_pin_25_;
wire [0:0] cby_1__1__23_left_grid_pin_26_;
wire [0:0] cby_1__1__23_left_grid_pin_27_;
wire [0:0] cby_1__1__23_left_grid_pin_28_;
wire [0:0] cby_1__1__23_left_grid_pin_29_;
wire [0:0] cby_1__1__23_left_grid_pin_30_;
wire [0:0] cby_1__1__23_left_grid_pin_31_;
wire [0:0] cby_1__1__24_ccff_tail;
wire [0:19] cby_1__1__24_chany_bottom_out;
wire [0:19] cby_1__1__24_chany_top_out;
wire [0:0] cby_1__1__24_left_grid_pin_16_;
wire [0:0] cby_1__1__24_left_grid_pin_17_;
wire [0:0] cby_1__1__24_left_grid_pin_18_;
wire [0:0] cby_1__1__24_left_grid_pin_19_;
wire [0:0] cby_1__1__24_left_grid_pin_20_;
wire [0:0] cby_1__1__24_left_grid_pin_21_;
wire [0:0] cby_1__1__24_left_grid_pin_22_;
wire [0:0] cby_1__1__24_left_grid_pin_23_;
wire [0:0] cby_1__1__24_left_grid_pin_24_;
wire [0:0] cby_1__1__24_left_grid_pin_25_;
wire [0:0] cby_1__1__24_left_grid_pin_26_;
wire [0:0] cby_1__1__24_left_grid_pin_27_;
wire [0:0] cby_1__1__24_left_grid_pin_28_;
wire [0:0] cby_1__1__24_left_grid_pin_29_;
wire [0:0] cby_1__1__24_left_grid_pin_30_;
wire [0:0] cby_1__1__24_left_grid_pin_31_;
wire [0:0] cby_1__1__25_ccff_tail;
wire [0:19] cby_1__1__25_chany_bottom_out;
wire [0:19] cby_1__1__25_chany_top_out;
wire [0:0] cby_1__1__25_left_grid_pin_16_;
wire [0:0] cby_1__1__25_left_grid_pin_17_;
wire [0:0] cby_1__1__25_left_grid_pin_18_;
wire [0:0] cby_1__1__25_left_grid_pin_19_;
wire [0:0] cby_1__1__25_left_grid_pin_20_;
wire [0:0] cby_1__1__25_left_grid_pin_21_;
wire [0:0] cby_1__1__25_left_grid_pin_22_;
wire [0:0] cby_1__1__25_left_grid_pin_23_;
wire [0:0] cby_1__1__25_left_grid_pin_24_;
wire [0:0] cby_1__1__25_left_grid_pin_25_;
wire [0:0] cby_1__1__25_left_grid_pin_26_;
wire [0:0] cby_1__1__25_left_grid_pin_27_;
wire [0:0] cby_1__1__25_left_grid_pin_28_;
wire [0:0] cby_1__1__25_left_grid_pin_29_;
wire [0:0] cby_1__1__25_left_grid_pin_30_;
wire [0:0] cby_1__1__25_left_grid_pin_31_;
wire [0:0] cby_1__1__26_ccff_tail;
wire [0:19] cby_1__1__26_chany_bottom_out;
wire [0:19] cby_1__1__26_chany_top_out;
wire [0:0] cby_1__1__26_left_grid_pin_16_;
wire [0:0] cby_1__1__26_left_grid_pin_17_;
wire [0:0] cby_1__1__26_left_grid_pin_18_;
wire [0:0] cby_1__1__26_left_grid_pin_19_;
wire [0:0] cby_1__1__26_left_grid_pin_20_;
wire [0:0] cby_1__1__26_left_grid_pin_21_;
wire [0:0] cby_1__1__26_left_grid_pin_22_;
wire [0:0] cby_1__1__26_left_grid_pin_23_;
wire [0:0] cby_1__1__26_left_grid_pin_24_;
wire [0:0] cby_1__1__26_left_grid_pin_25_;
wire [0:0] cby_1__1__26_left_grid_pin_26_;
wire [0:0] cby_1__1__26_left_grid_pin_27_;
wire [0:0] cby_1__1__26_left_grid_pin_28_;
wire [0:0] cby_1__1__26_left_grid_pin_29_;
wire [0:0] cby_1__1__26_left_grid_pin_30_;
wire [0:0] cby_1__1__26_left_grid_pin_31_;
wire [0:0] cby_1__1__27_ccff_tail;
wire [0:19] cby_1__1__27_chany_bottom_out;
wire [0:19] cby_1__1__27_chany_top_out;
wire [0:0] cby_1__1__27_left_grid_pin_16_;
wire [0:0] cby_1__1__27_left_grid_pin_17_;
wire [0:0] cby_1__1__27_left_grid_pin_18_;
wire [0:0] cby_1__1__27_left_grid_pin_19_;
wire [0:0] cby_1__1__27_left_grid_pin_20_;
wire [0:0] cby_1__1__27_left_grid_pin_21_;
wire [0:0] cby_1__1__27_left_grid_pin_22_;
wire [0:0] cby_1__1__27_left_grid_pin_23_;
wire [0:0] cby_1__1__27_left_grid_pin_24_;
wire [0:0] cby_1__1__27_left_grid_pin_25_;
wire [0:0] cby_1__1__27_left_grid_pin_26_;
wire [0:0] cby_1__1__27_left_grid_pin_27_;
wire [0:0] cby_1__1__27_left_grid_pin_28_;
wire [0:0] cby_1__1__27_left_grid_pin_29_;
wire [0:0] cby_1__1__27_left_grid_pin_30_;
wire [0:0] cby_1__1__27_left_grid_pin_31_;
wire [0:0] cby_1__1__28_ccff_tail;
wire [0:19] cby_1__1__28_chany_bottom_out;
wire [0:19] cby_1__1__28_chany_top_out;
wire [0:0] cby_1__1__28_left_grid_pin_16_;
wire [0:0] cby_1__1__28_left_grid_pin_17_;
wire [0:0] cby_1__1__28_left_grid_pin_18_;
wire [0:0] cby_1__1__28_left_grid_pin_19_;
wire [0:0] cby_1__1__28_left_grid_pin_20_;
wire [0:0] cby_1__1__28_left_grid_pin_21_;
wire [0:0] cby_1__1__28_left_grid_pin_22_;
wire [0:0] cby_1__1__28_left_grid_pin_23_;
wire [0:0] cby_1__1__28_left_grid_pin_24_;
wire [0:0] cby_1__1__28_left_grid_pin_25_;
wire [0:0] cby_1__1__28_left_grid_pin_26_;
wire [0:0] cby_1__1__28_left_grid_pin_27_;
wire [0:0] cby_1__1__28_left_grid_pin_28_;
wire [0:0] cby_1__1__28_left_grid_pin_29_;
wire [0:0] cby_1__1__28_left_grid_pin_30_;
wire [0:0] cby_1__1__28_left_grid_pin_31_;
wire [0:0] cby_1__1__29_ccff_tail;
wire [0:19] cby_1__1__29_chany_bottom_out;
wire [0:19] cby_1__1__29_chany_top_out;
wire [0:0] cby_1__1__29_left_grid_pin_16_;
wire [0:0] cby_1__1__29_left_grid_pin_17_;
wire [0:0] cby_1__1__29_left_grid_pin_18_;
wire [0:0] cby_1__1__29_left_grid_pin_19_;
wire [0:0] cby_1__1__29_left_grid_pin_20_;
wire [0:0] cby_1__1__29_left_grid_pin_21_;
wire [0:0] cby_1__1__29_left_grid_pin_22_;
wire [0:0] cby_1__1__29_left_grid_pin_23_;
wire [0:0] cby_1__1__29_left_grid_pin_24_;
wire [0:0] cby_1__1__29_left_grid_pin_25_;
wire [0:0] cby_1__1__29_left_grid_pin_26_;
wire [0:0] cby_1__1__29_left_grid_pin_27_;
wire [0:0] cby_1__1__29_left_grid_pin_28_;
wire [0:0] cby_1__1__29_left_grid_pin_29_;
wire [0:0] cby_1__1__29_left_grid_pin_30_;
wire [0:0] cby_1__1__29_left_grid_pin_31_;
wire [0:0] cby_1__1__2_ccff_tail;
wire [0:19] cby_1__1__2_chany_bottom_out;
wire [0:19] cby_1__1__2_chany_top_out;
wire [0:0] cby_1__1__2_left_grid_pin_16_;
wire [0:0] cby_1__1__2_left_grid_pin_17_;
wire [0:0] cby_1__1__2_left_grid_pin_18_;
wire [0:0] cby_1__1__2_left_grid_pin_19_;
wire [0:0] cby_1__1__2_left_grid_pin_20_;
wire [0:0] cby_1__1__2_left_grid_pin_21_;
wire [0:0] cby_1__1__2_left_grid_pin_22_;
wire [0:0] cby_1__1__2_left_grid_pin_23_;
wire [0:0] cby_1__1__2_left_grid_pin_24_;
wire [0:0] cby_1__1__2_left_grid_pin_25_;
wire [0:0] cby_1__1__2_left_grid_pin_26_;
wire [0:0] cby_1__1__2_left_grid_pin_27_;
wire [0:0] cby_1__1__2_left_grid_pin_28_;
wire [0:0] cby_1__1__2_left_grid_pin_29_;
wire [0:0] cby_1__1__2_left_grid_pin_30_;
wire [0:0] cby_1__1__2_left_grid_pin_31_;
wire [0:0] cby_1__1__30_ccff_tail;
wire [0:19] cby_1__1__30_chany_bottom_out;
wire [0:19] cby_1__1__30_chany_top_out;
wire [0:0] cby_1__1__30_left_grid_pin_16_;
wire [0:0] cby_1__1__30_left_grid_pin_17_;
wire [0:0] cby_1__1__30_left_grid_pin_18_;
wire [0:0] cby_1__1__30_left_grid_pin_19_;
wire [0:0] cby_1__1__30_left_grid_pin_20_;
wire [0:0] cby_1__1__30_left_grid_pin_21_;
wire [0:0] cby_1__1__30_left_grid_pin_22_;
wire [0:0] cby_1__1__30_left_grid_pin_23_;
wire [0:0] cby_1__1__30_left_grid_pin_24_;
wire [0:0] cby_1__1__30_left_grid_pin_25_;
wire [0:0] cby_1__1__30_left_grid_pin_26_;
wire [0:0] cby_1__1__30_left_grid_pin_27_;
wire [0:0] cby_1__1__30_left_grid_pin_28_;
wire [0:0] cby_1__1__30_left_grid_pin_29_;
wire [0:0] cby_1__1__30_left_grid_pin_30_;
wire [0:0] cby_1__1__30_left_grid_pin_31_;
wire [0:0] cby_1__1__31_ccff_tail;
wire [0:19] cby_1__1__31_chany_bottom_out;
wire [0:19] cby_1__1__31_chany_top_out;
wire [0:0] cby_1__1__31_left_grid_pin_16_;
wire [0:0] cby_1__1__31_left_grid_pin_17_;
wire [0:0] cby_1__1__31_left_grid_pin_18_;
wire [0:0] cby_1__1__31_left_grid_pin_19_;
wire [0:0] cby_1__1__31_left_grid_pin_20_;
wire [0:0] cby_1__1__31_left_grid_pin_21_;
wire [0:0] cby_1__1__31_left_grid_pin_22_;
wire [0:0] cby_1__1__31_left_grid_pin_23_;
wire [0:0] cby_1__1__31_left_grid_pin_24_;
wire [0:0] cby_1__1__31_left_grid_pin_25_;
wire [0:0] cby_1__1__31_left_grid_pin_26_;
wire [0:0] cby_1__1__31_left_grid_pin_27_;
wire [0:0] cby_1__1__31_left_grid_pin_28_;
wire [0:0] cby_1__1__31_left_grid_pin_29_;
wire [0:0] cby_1__1__31_left_grid_pin_30_;
wire [0:0] cby_1__1__31_left_grid_pin_31_;
wire [0:0] cby_1__1__32_ccff_tail;
wire [0:19] cby_1__1__32_chany_bottom_out;
wire [0:19] cby_1__1__32_chany_top_out;
wire [0:0] cby_1__1__32_left_grid_pin_16_;
wire [0:0] cby_1__1__32_left_grid_pin_17_;
wire [0:0] cby_1__1__32_left_grid_pin_18_;
wire [0:0] cby_1__1__32_left_grid_pin_19_;
wire [0:0] cby_1__1__32_left_grid_pin_20_;
wire [0:0] cby_1__1__32_left_grid_pin_21_;
wire [0:0] cby_1__1__32_left_grid_pin_22_;
wire [0:0] cby_1__1__32_left_grid_pin_23_;
wire [0:0] cby_1__1__32_left_grid_pin_24_;
wire [0:0] cby_1__1__32_left_grid_pin_25_;
wire [0:0] cby_1__1__32_left_grid_pin_26_;
wire [0:0] cby_1__1__32_left_grid_pin_27_;
wire [0:0] cby_1__1__32_left_grid_pin_28_;
wire [0:0] cby_1__1__32_left_grid_pin_29_;
wire [0:0] cby_1__1__32_left_grid_pin_30_;
wire [0:0] cby_1__1__32_left_grid_pin_31_;
wire [0:0] cby_1__1__33_ccff_tail;
wire [0:19] cby_1__1__33_chany_bottom_out;
wire [0:19] cby_1__1__33_chany_top_out;
wire [0:0] cby_1__1__33_left_grid_pin_16_;
wire [0:0] cby_1__1__33_left_grid_pin_17_;
wire [0:0] cby_1__1__33_left_grid_pin_18_;
wire [0:0] cby_1__1__33_left_grid_pin_19_;
wire [0:0] cby_1__1__33_left_grid_pin_20_;
wire [0:0] cby_1__1__33_left_grid_pin_21_;
wire [0:0] cby_1__1__33_left_grid_pin_22_;
wire [0:0] cby_1__1__33_left_grid_pin_23_;
wire [0:0] cby_1__1__33_left_grid_pin_24_;
wire [0:0] cby_1__1__33_left_grid_pin_25_;
wire [0:0] cby_1__1__33_left_grid_pin_26_;
wire [0:0] cby_1__1__33_left_grid_pin_27_;
wire [0:0] cby_1__1__33_left_grid_pin_28_;
wire [0:0] cby_1__1__33_left_grid_pin_29_;
wire [0:0] cby_1__1__33_left_grid_pin_30_;
wire [0:0] cby_1__1__33_left_grid_pin_31_;
wire [0:0] cby_1__1__34_ccff_tail;
wire [0:19] cby_1__1__34_chany_bottom_out;
wire [0:19] cby_1__1__34_chany_top_out;
wire [0:0] cby_1__1__34_left_grid_pin_16_;
wire [0:0] cby_1__1__34_left_grid_pin_17_;
wire [0:0] cby_1__1__34_left_grid_pin_18_;
wire [0:0] cby_1__1__34_left_grid_pin_19_;
wire [0:0] cby_1__1__34_left_grid_pin_20_;
wire [0:0] cby_1__1__34_left_grid_pin_21_;
wire [0:0] cby_1__1__34_left_grid_pin_22_;
wire [0:0] cby_1__1__34_left_grid_pin_23_;
wire [0:0] cby_1__1__34_left_grid_pin_24_;
wire [0:0] cby_1__1__34_left_grid_pin_25_;
wire [0:0] cby_1__1__34_left_grid_pin_26_;
wire [0:0] cby_1__1__34_left_grid_pin_27_;
wire [0:0] cby_1__1__34_left_grid_pin_28_;
wire [0:0] cby_1__1__34_left_grid_pin_29_;
wire [0:0] cby_1__1__34_left_grid_pin_30_;
wire [0:0] cby_1__1__34_left_grid_pin_31_;
wire [0:0] cby_1__1__35_ccff_tail;
wire [0:19] cby_1__1__35_chany_bottom_out;
wire [0:19] cby_1__1__35_chany_top_out;
wire [0:0] cby_1__1__35_left_grid_pin_16_;
wire [0:0] cby_1__1__35_left_grid_pin_17_;
wire [0:0] cby_1__1__35_left_grid_pin_18_;
wire [0:0] cby_1__1__35_left_grid_pin_19_;
wire [0:0] cby_1__1__35_left_grid_pin_20_;
wire [0:0] cby_1__1__35_left_grid_pin_21_;
wire [0:0] cby_1__1__35_left_grid_pin_22_;
wire [0:0] cby_1__1__35_left_grid_pin_23_;
wire [0:0] cby_1__1__35_left_grid_pin_24_;
wire [0:0] cby_1__1__35_left_grid_pin_25_;
wire [0:0] cby_1__1__35_left_grid_pin_26_;
wire [0:0] cby_1__1__35_left_grid_pin_27_;
wire [0:0] cby_1__1__35_left_grid_pin_28_;
wire [0:0] cby_1__1__35_left_grid_pin_29_;
wire [0:0] cby_1__1__35_left_grid_pin_30_;
wire [0:0] cby_1__1__35_left_grid_pin_31_;
wire [0:0] cby_1__1__36_ccff_tail;
wire [0:19] cby_1__1__36_chany_bottom_out;
wire [0:19] cby_1__1__36_chany_top_out;
wire [0:0] cby_1__1__36_left_grid_pin_16_;
wire [0:0] cby_1__1__36_left_grid_pin_17_;
wire [0:0] cby_1__1__36_left_grid_pin_18_;
wire [0:0] cby_1__1__36_left_grid_pin_19_;
wire [0:0] cby_1__1__36_left_grid_pin_20_;
wire [0:0] cby_1__1__36_left_grid_pin_21_;
wire [0:0] cby_1__1__36_left_grid_pin_22_;
wire [0:0] cby_1__1__36_left_grid_pin_23_;
wire [0:0] cby_1__1__36_left_grid_pin_24_;
wire [0:0] cby_1__1__36_left_grid_pin_25_;
wire [0:0] cby_1__1__36_left_grid_pin_26_;
wire [0:0] cby_1__1__36_left_grid_pin_27_;
wire [0:0] cby_1__1__36_left_grid_pin_28_;
wire [0:0] cby_1__1__36_left_grid_pin_29_;
wire [0:0] cby_1__1__36_left_grid_pin_30_;
wire [0:0] cby_1__1__36_left_grid_pin_31_;
wire [0:0] cby_1__1__37_ccff_tail;
wire [0:19] cby_1__1__37_chany_bottom_out;
wire [0:19] cby_1__1__37_chany_top_out;
wire [0:0] cby_1__1__37_left_grid_pin_16_;
wire [0:0] cby_1__1__37_left_grid_pin_17_;
wire [0:0] cby_1__1__37_left_grid_pin_18_;
wire [0:0] cby_1__1__37_left_grid_pin_19_;
wire [0:0] cby_1__1__37_left_grid_pin_20_;
wire [0:0] cby_1__1__37_left_grid_pin_21_;
wire [0:0] cby_1__1__37_left_grid_pin_22_;
wire [0:0] cby_1__1__37_left_grid_pin_23_;
wire [0:0] cby_1__1__37_left_grid_pin_24_;
wire [0:0] cby_1__1__37_left_grid_pin_25_;
wire [0:0] cby_1__1__37_left_grid_pin_26_;
wire [0:0] cby_1__1__37_left_grid_pin_27_;
wire [0:0] cby_1__1__37_left_grid_pin_28_;
wire [0:0] cby_1__1__37_left_grid_pin_29_;
wire [0:0] cby_1__1__37_left_grid_pin_30_;
wire [0:0] cby_1__1__37_left_grid_pin_31_;
wire [0:0] cby_1__1__38_ccff_tail;
wire [0:19] cby_1__1__38_chany_bottom_out;
wire [0:19] cby_1__1__38_chany_top_out;
wire [0:0] cby_1__1__38_left_grid_pin_16_;
wire [0:0] cby_1__1__38_left_grid_pin_17_;
wire [0:0] cby_1__1__38_left_grid_pin_18_;
wire [0:0] cby_1__1__38_left_grid_pin_19_;
wire [0:0] cby_1__1__38_left_grid_pin_20_;
wire [0:0] cby_1__1__38_left_grid_pin_21_;
wire [0:0] cby_1__1__38_left_grid_pin_22_;
wire [0:0] cby_1__1__38_left_grid_pin_23_;
wire [0:0] cby_1__1__38_left_grid_pin_24_;
wire [0:0] cby_1__1__38_left_grid_pin_25_;
wire [0:0] cby_1__1__38_left_grid_pin_26_;
wire [0:0] cby_1__1__38_left_grid_pin_27_;
wire [0:0] cby_1__1__38_left_grid_pin_28_;
wire [0:0] cby_1__1__38_left_grid_pin_29_;
wire [0:0] cby_1__1__38_left_grid_pin_30_;
wire [0:0] cby_1__1__38_left_grid_pin_31_;
wire [0:0] cby_1__1__39_ccff_tail;
wire [0:19] cby_1__1__39_chany_bottom_out;
wire [0:19] cby_1__1__39_chany_top_out;
wire [0:0] cby_1__1__39_left_grid_pin_16_;
wire [0:0] cby_1__1__39_left_grid_pin_17_;
wire [0:0] cby_1__1__39_left_grid_pin_18_;
wire [0:0] cby_1__1__39_left_grid_pin_19_;
wire [0:0] cby_1__1__39_left_grid_pin_20_;
wire [0:0] cby_1__1__39_left_grid_pin_21_;
wire [0:0] cby_1__1__39_left_grid_pin_22_;
wire [0:0] cby_1__1__39_left_grid_pin_23_;
wire [0:0] cby_1__1__39_left_grid_pin_24_;
wire [0:0] cby_1__1__39_left_grid_pin_25_;
wire [0:0] cby_1__1__39_left_grid_pin_26_;
wire [0:0] cby_1__1__39_left_grid_pin_27_;
wire [0:0] cby_1__1__39_left_grid_pin_28_;
wire [0:0] cby_1__1__39_left_grid_pin_29_;
wire [0:0] cby_1__1__39_left_grid_pin_30_;
wire [0:0] cby_1__1__39_left_grid_pin_31_;
wire [0:0] cby_1__1__3_ccff_tail;
wire [0:19] cby_1__1__3_chany_bottom_out;
wire [0:19] cby_1__1__3_chany_top_out;
wire [0:0] cby_1__1__3_left_grid_pin_16_;
wire [0:0] cby_1__1__3_left_grid_pin_17_;
wire [0:0] cby_1__1__3_left_grid_pin_18_;
wire [0:0] cby_1__1__3_left_grid_pin_19_;
wire [0:0] cby_1__1__3_left_grid_pin_20_;
wire [0:0] cby_1__1__3_left_grid_pin_21_;
wire [0:0] cby_1__1__3_left_grid_pin_22_;
wire [0:0] cby_1__1__3_left_grid_pin_23_;
wire [0:0] cby_1__1__3_left_grid_pin_24_;
wire [0:0] cby_1__1__3_left_grid_pin_25_;
wire [0:0] cby_1__1__3_left_grid_pin_26_;
wire [0:0] cby_1__1__3_left_grid_pin_27_;
wire [0:0] cby_1__1__3_left_grid_pin_28_;
wire [0:0] cby_1__1__3_left_grid_pin_29_;
wire [0:0] cby_1__1__3_left_grid_pin_30_;
wire [0:0] cby_1__1__3_left_grid_pin_31_;
wire [0:0] cby_1__1__40_ccff_tail;
wire [0:19] cby_1__1__40_chany_bottom_out;
wire [0:19] cby_1__1__40_chany_top_out;
wire [0:0] cby_1__1__40_left_grid_pin_16_;
wire [0:0] cby_1__1__40_left_grid_pin_17_;
wire [0:0] cby_1__1__40_left_grid_pin_18_;
wire [0:0] cby_1__1__40_left_grid_pin_19_;
wire [0:0] cby_1__1__40_left_grid_pin_20_;
wire [0:0] cby_1__1__40_left_grid_pin_21_;
wire [0:0] cby_1__1__40_left_grid_pin_22_;
wire [0:0] cby_1__1__40_left_grid_pin_23_;
wire [0:0] cby_1__1__40_left_grid_pin_24_;
wire [0:0] cby_1__1__40_left_grid_pin_25_;
wire [0:0] cby_1__1__40_left_grid_pin_26_;
wire [0:0] cby_1__1__40_left_grid_pin_27_;
wire [0:0] cby_1__1__40_left_grid_pin_28_;
wire [0:0] cby_1__1__40_left_grid_pin_29_;
wire [0:0] cby_1__1__40_left_grid_pin_30_;
wire [0:0] cby_1__1__40_left_grid_pin_31_;
wire [0:0] cby_1__1__41_ccff_tail;
wire [0:19] cby_1__1__41_chany_bottom_out;
wire [0:19] cby_1__1__41_chany_top_out;
wire [0:0] cby_1__1__41_left_grid_pin_16_;
wire [0:0] cby_1__1__41_left_grid_pin_17_;
wire [0:0] cby_1__1__41_left_grid_pin_18_;
wire [0:0] cby_1__1__41_left_grid_pin_19_;
wire [0:0] cby_1__1__41_left_grid_pin_20_;
wire [0:0] cby_1__1__41_left_grid_pin_21_;
wire [0:0] cby_1__1__41_left_grid_pin_22_;
wire [0:0] cby_1__1__41_left_grid_pin_23_;
wire [0:0] cby_1__1__41_left_grid_pin_24_;
wire [0:0] cby_1__1__41_left_grid_pin_25_;
wire [0:0] cby_1__1__41_left_grid_pin_26_;
wire [0:0] cby_1__1__41_left_grid_pin_27_;
wire [0:0] cby_1__1__41_left_grid_pin_28_;
wire [0:0] cby_1__1__41_left_grid_pin_29_;
wire [0:0] cby_1__1__41_left_grid_pin_30_;
wire [0:0] cby_1__1__41_left_grid_pin_31_;
wire [0:0] cby_1__1__42_ccff_tail;
wire [0:19] cby_1__1__42_chany_bottom_out;
wire [0:19] cby_1__1__42_chany_top_out;
wire [0:0] cby_1__1__42_left_grid_pin_16_;
wire [0:0] cby_1__1__42_left_grid_pin_17_;
wire [0:0] cby_1__1__42_left_grid_pin_18_;
wire [0:0] cby_1__1__42_left_grid_pin_19_;
wire [0:0] cby_1__1__42_left_grid_pin_20_;
wire [0:0] cby_1__1__42_left_grid_pin_21_;
wire [0:0] cby_1__1__42_left_grid_pin_22_;
wire [0:0] cby_1__1__42_left_grid_pin_23_;
wire [0:0] cby_1__1__42_left_grid_pin_24_;
wire [0:0] cby_1__1__42_left_grid_pin_25_;
wire [0:0] cby_1__1__42_left_grid_pin_26_;
wire [0:0] cby_1__1__42_left_grid_pin_27_;
wire [0:0] cby_1__1__42_left_grid_pin_28_;
wire [0:0] cby_1__1__42_left_grid_pin_29_;
wire [0:0] cby_1__1__42_left_grid_pin_30_;
wire [0:0] cby_1__1__42_left_grid_pin_31_;
wire [0:0] cby_1__1__43_ccff_tail;
wire [0:19] cby_1__1__43_chany_bottom_out;
wire [0:19] cby_1__1__43_chany_top_out;
wire [0:0] cby_1__1__43_left_grid_pin_16_;
wire [0:0] cby_1__1__43_left_grid_pin_17_;
wire [0:0] cby_1__1__43_left_grid_pin_18_;
wire [0:0] cby_1__1__43_left_grid_pin_19_;
wire [0:0] cby_1__1__43_left_grid_pin_20_;
wire [0:0] cby_1__1__43_left_grid_pin_21_;
wire [0:0] cby_1__1__43_left_grid_pin_22_;
wire [0:0] cby_1__1__43_left_grid_pin_23_;
wire [0:0] cby_1__1__43_left_grid_pin_24_;
wire [0:0] cby_1__1__43_left_grid_pin_25_;
wire [0:0] cby_1__1__43_left_grid_pin_26_;
wire [0:0] cby_1__1__43_left_grid_pin_27_;
wire [0:0] cby_1__1__43_left_grid_pin_28_;
wire [0:0] cby_1__1__43_left_grid_pin_29_;
wire [0:0] cby_1__1__43_left_grid_pin_30_;
wire [0:0] cby_1__1__43_left_grid_pin_31_;
wire [0:0] cby_1__1__44_ccff_tail;
wire [0:19] cby_1__1__44_chany_bottom_out;
wire [0:19] cby_1__1__44_chany_top_out;
wire [0:0] cby_1__1__44_left_grid_pin_16_;
wire [0:0] cby_1__1__44_left_grid_pin_17_;
wire [0:0] cby_1__1__44_left_grid_pin_18_;
wire [0:0] cby_1__1__44_left_grid_pin_19_;
wire [0:0] cby_1__1__44_left_grid_pin_20_;
wire [0:0] cby_1__1__44_left_grid_pin_21_;
wire [0:0] cby_1__1__44_left_grid_pin_22_;
wire [0:0] cby_1__1__44_left_grid_pin_23_;
wire [0:0] cby_1__1__44_left_grid_pin_24_;
wire [0:0] cby_1__1__44_left_grid_pin_25_;
wire [0:0] cby_1__1__44_left_grid_pin_26_;
wire [0:0] cby_1__1__44_left_grid_pin_27_;
wire [0:0] cby_1__1__44_left_grid_pin_28_;
wire [0:0] cby_1__1__44_left_grid_pin_29_;
wire [0:0] cby_1__1__44_left_grid_pin_30_;
wire [0:0] cby_1__1__44_left_grid_pin_31_;
wire [0:0] cby_1__1__45_ccff_tail;
wire [0:19] cby_1__1__45_chany_bottom_out;
wire [0:19] cby_1__1__45_chany_top_out;
wire [0:0] cby_1__1__45_left_grid_pin_16_;
wire [0:0] cby_1__1__45_left_grid_pin_17_;
wire [0:0] cby_1__1__45_left_grid_pin_18_;
wire [0:0] cby_1__1__45_left_grid_pin_19_;
wire [0:0] cby_1__1__45_left_grid_pin_20_;
wire [0:0] cby_1__1__45_left_grid_pin_21_;
wire [0:0] cby_1__1__45_left_grid_pin_22_;
wire [0:0] cby_1__1__45_left_grid_pin_23_;
wire [0:0] cby_1__1__45_left_grid_pin_24_;
wire [0:0] cby_1__1__45_left_grid_pin_25_;
wire [0:0] cby_1__1__45_left_grid_pin_26_;
wire [0:0] cby_1__1__45_left_grid_pin_27_;
wire [0:0] cby_1__1__45_left_grid_pin_28_;
wire [0:0] cby_1__1__45_left_grid_pin_29_;
wire [0:0] cby_1__1__45_left_grid_pin_30_;
wire [0:0] cby_1__1__45_left_grid_pin_31_;
wire [0:0] cby_1__1__46_ccff_tail;
wire [0:19] cby_1__1__46_chany_bottom_out;
wire [0:19] cby_1__1__46_chany_top_out;
wire [0:0] cby_1__1__46_left_grid_pin_16_;
wire [0:0] cby_1__1__46_left_grid_pin_17_;
wire [0:0] cby_1__1__46_left_grid_pin_18_;
wire [0:0] cby_1__1__46_left_grid_pin_19_;
wire [0:0] cby_1__1__46_left_grid_pin_20_;
wire [0:0] cby_1__1__46_left_grid_pin_21_;
wire [0:0] cby_1__1__46_left_grid_pin_22_;
wire [0:0] cby_1__1__46_left_grid_pin_23_;
wire [0:0] cby_1__1__46_left_grid_pin_24_;
wire [0:0] cby_1__1__46_left_grid_pin_25_;
wire [0:0] cby_1__1__46_left_grid_pin_26_;
wire [0:0] cby_1__1__46_left_grid_pin_27_;
wire [0:0] cby_1__1__46_left_grid_pin_28_;
wire [0:0] cby_1__1__46_left_grid_pin_29_;
wire [0:0] cby_1__1__46_left_grid_pin_30_;
wire [0:0] cby_1__1__46_left_grid_pin_31_;
wire [0:0] cby_1__1__47_ccff_tail;
wire [0:19] cby_1__1__47_chany_bottom_out;
wire [0:19] cby_1__1__47_chany_top_out;
wire [0:0] cby_1__1__47_left_grid_pin_16_;
wire [0:0] cby_1__1__47_left_grid_pin_17_;
wire [0:0] cby_1__1__47_left_grid_pin_18_;
wire [0:0] cby_1__1__47_left_grid_pin_19_;
wire [0:0] cby_1__1__47_left_grid_pin_20_;
wire [0:0] cby_1__1__47_left_grid_pin_21_;
wire [0:0] cby_1__1__47_left_grid_pin_22_;
wire [0:0] cby_1__1__47_left_grid_pin_23_;
wire [0:0] cby_1__1__47_left_grid_pin_24_;
wire [0:0] cby_1__1__47_left_grid_pin_25_;
wire [0:0] cby_1__1__47_left_grid_pin_26_;
wire [0:0] cby_1__1__47_left_grid_pin_27_;
wire [0:0] cby_1__1__47_left_grid_pin_28_;
wire [0:0] cby_1__1__47_left_grid_pin_29_;
wire [0:0] cby_1__1__47_left_grid_pin_30_;
wire [0:0] cby_1__1__47_left_grid_pin_31_;
wire [0:0] cby_1__1__48_ccff_tail;
wire [0:19] cby_1__1__48_chany_bottom_out;
wire [0:19] cby_1__1__48_chany_top_out;
wire [0:0] cby_1__1__48_left_grid_pin_16_;
wire [0:0] cby_1__1__48_left_grid_pin_17_;
wire [0:0] cby_1__1__48_left_grid_pin_18_;
wire [0:0] cby_1__1__48_left_grid_pin_19_;
wire [0:0] cby_1__1__48_left_grid_pin_20_;
wire [0:0] cby_1__1__48_left_grid_pin_21_;
wire [0:0] cby_1__1__48_left_grid_pin_22_;
wire [0:0] cby_1__1__48_left_grid_pin_23_;
wire [0:0] cby_1__1__48_left_grid_pin_24_;
wire [0:0] cby_1__1__48_left_grid_pin_25_;
wire [0:0] cby_1__1__48_left_grid_pin_26_;
wire [0:0] cby_1__1__48_left_grid_pin_27_;
wire [0:0] cby_1__1__48_left_grid_pin_28_;
wire [0:0] cby_1__1__48_left_grid_pin_29_;
wire [0:0] cby_1__1__48_left_grid_pin_30_;
wire [0:0] cby_1__1__48_left_grid_pin_31_;
wire [0:0] cby_1__1__49_ccff_tail;
wire [0:19] cby_1__1__49_chany_bottom_out;
wire [0:19] cby_1__1__49_chany_top_out;
wire [0:0] cby_1__1__49_left_grid_pin_16_;
wire [0:0] cby_1__1__49_left_grid_pin_17_;
wire [0:0] cby_1__1__49_left_grid_pin_18_;
wire [0:0] cby_1__1__49_left_grid_pin_19_;
wire [0:0] cby_1__1__49_left_grid_pin_20_;
wire [0:0] cby_1__1__49_left_grid_pin_21_;
wire [0:0] cby_1__1__49_left_grid_pin_22_;
wire [0:0] cby_1__1__49_left_grid_pin_23_;
wire [0:0] cby_1__1__49_left_grid_pin_24_;
wire [0:0] cby_1__1__49_left_grid_pin_25_;
wire [0:0] cby_1__1__49_left_grid_pin_26_;
wire [0:0] cby_1__1__49_left_grid_pin_27_;
wire [0:0] cby_1__1__49_left_grid_pin_28_;
wire [0:0] cby_1__1__49_left_grid_pin_29_;
wire [0:0] cby_1__1__49_left_grid_pin_30_;
wire [0:0] cby_1__1__49_left_grid_pin_31_;
wire [0:0] cby_1__1__4_ccff_tail;
wire [0:19] cby_1__1__4_chany_bottom_out;
wire [0:19] cby_1__1__4_chany_top_out;
wire [0:0] cby_1__1__4_left_grid_pin_16_;
wire [0:0] cby_1__1__4_left_grid_pin_17_;
wire [0:0] cby_1__1__4_left_grid_pin_18_;
wire [0:0] cby_1__1__4_left_grid_pin_19_;
wire [0:0] cby_1__1__4_left_grid_pin_20_;
wire [0:0] cby_1__1__4_left_grid_pin_21_;
wire [0:0] cby_1__1__4_left_grid_pin_22_;
wire [0:0] cby_1__1__4_left_grid_pin_23_;
wire [0:0] cby_1__1__4_left_grid_pin_24_;
wire [0:0] cby_1__1__4_left_grid_pin_25_;
wire [0:0] cby_1__1__4_left_grid_pin_26_;
wire [0:0] cby_1__1__4_left_grid_pin_27_;
wire [0:0] cby_1__1__4_left_grid_pin_28_;
wire [0:0] cby_1__1__4_left_grid_pin_29_;
wire [0:0] cby_1__1__4_left_grid_pin_30_;
wire [0:0] cby_1__1__4_left_grid_pin_31_;
wire [0:0] cby_1__1__50_ccff_tail;
wire [0:19] cby_1__1__50_chany_bottom_out;
wire [0:19] cby_1__1__50_chany_top_out;
wire [0:0] cby_1__1__50_left_grid_pin_16_;
wire [0:0] cby_1__1__50_left_grid_pin_17_;
wire [0:0] cby_1__1__50_left_grid_pin_18_;
wire [0:0] cby_1__1__50_left_grid_pin_19_;
wire [0:0] cby_1__1__50_left_grid_pin_20_;
wire [0:0] cby_1__1__50_left_grid_pin_21_;
wire [0:0] cby_1__1__50_left_grid_pin_22_;
wire [0:0] cby_1__1__50_left_grid_pin_23_;
wire [0:0] cby_1__1__50_left_grid_pin_24_;
wire [0:0] cby_1__1__50_left_grid_pin_25_;
wire [0:0] cby_1__1__50_left_grid_pin_26_;
wire [0:0] cby_1__1__50_left_grid_pin_27_;
wire [0:0] cby_1__1__50_left_grid_pin_28_;
wire [0:0] cby_1__1__50_left_grid_pin_29_;
wire [0:0] cby_1__1__50_left_grid_pin_30_;
wire [0:0] cby_1__1__50_left_grid_pin_31_;
wire [0:0] cby_1__1__51_ccff_tail;
wire [0:19] cby_1__1__51_chany_bottom_out;
wire [0:19] cby_1__1__51_chany_top_out;
wire [0:0] cby_1__1__51_left_grid_pin_16_;
wire [0:0] cby_1__1__51_left_grid_pin_17_;
wire [0:0] cby_1__1__51_left_grid_pin_18_;
wire [0:0] cby_1__1__51_left_grid_pin_19_;
wire [0:0] cby_1__1__51_left_grid_pin_20_;
wire [0:0] cby_1__1__51_left_grid_pin_21_;
wire [0:0] cby_1__1__51_left_grid_pin_22_;
wire [0:0] cby_1__1__51_left_grid_pin_23_;
wire [0:0] cby_1__1__51_left_grid_pin_24_;
wire [0:0] cby_1__1__51_left_grid_pin_25_;
wire [0:0] cby_1__1__51_left_grid_pin_26_;
wire [0:0] cby_1__1__51_left_grid_pin_27_;
wire [0:0] cby_1__1__51_left_grid_pin_28_;
wire [0:0] cby_1__1__51_left_grid_pin_29_;
wire [0:0] cby_1__1__51_left_grid_pin_30_;
wire [0:0] cby_1__1__51_left_grid_pin_31_;
wire [0:0] cby_1__1__52_ccff_tail;
wire [0:19] cby_1__1__52_chany_bottom_out;
wire [0:19] cby_1__1__52_chany_top_out;
wire [0:0] cby_1__1__52_left_grid_pin_16_;
wire [0:0] cby_1__1__52_left_grid_pin_17_;
wire [0:0] cby_1__1__52_left_grid_pin_18_;
wire [0:0] cby_1__1__52_left_grid_pin_19_;
wire [0:0] cby_1__1__52_left_grid_pin_20_;
wire [0:0] cby_1__1__52_left_grid_pin_21_;
wire [0:0] cby_1__1__52_left_grid_pin_22_;
wire [0:0] cby_1__1__52_left_grid_pin_23_;
wire [0:0] cby_1__1__52_left_grid_pin_24_;
wire [0:0] cby_1__1__52_left_grid_pin_25_;
wire [0:0] cby_1__1__52_left_grid_pin_26_;
wire [0:0] cby_1__1__52_left_grid_pin_27_;
wire [0:0] cby_1__1__52_left_grid_pin_28_;
wire [0:0] cby_1__1__52_left_grid_pin_29_;
wire [0:0] cby_1__1__52_left_grid_pin_30_;
wire [0:0] cby_1__1__52_left_grid_pin_31_;
wire [0:0] cby_1__1__53_ccff_tail;
wire [0:19] cby_1__1__53_chany_bottom_out;
wire [0:19] cby_1__1__53_chany_top_out;
wire [0:0] cby_1__1__53_left_grid_pin_16_;
wire [0:0] cby_1__1__53_left_grid_pin_17_;
wire [0:0] cby_1__1__53_left_grid_pin_18_;
wire [0:0] cby_1__1__53_left_grid_pin_19_;
wire [0:0] cby_1__1__53_left_grid_pin_20_;
wire [0:0] cby_1__1__53_left_grid_pin_21_;
wire [0:0] cby_1__1__53_left_grid_pin_22_;
wire [0:0] cby_1__1__53_left_grid_pin_23_;
wire [0:0] cby_1__1__53_left_grid_pin_24_;
wire [0:0] cby_1__1__53_left_grid_pin_25_;
wire [0:0] cby_1__1__53_left_grid_pin_26_;
wire [0:0] cby_1__1__53_left_grid_pin_27_;
wire [0:0] cby_1__1__53_left_grid_pin_28_;
wire [0:0] cby_1__1__53_left_grid_pin_29_;
wire [0:0] cby_1__1__53_left_grid_pin_30_;
wire [0:0] cby_1__1__53_left_grid_pin_31_;
wire [0:0] cby_1__1__54_ccff_tail;
wire [0:19] cby_1__1__54_chany_bottom_out;
wire [0:19] cby_1__1__54_chany_top_out;
wire [0:0] cby_1__1__54_left_grid_pin_16_;
wire [0:0] cby_1__1__54_left_grid_pin_17_;
wire [0:0] cby_1__1__54_left_grid_pin_18_;
wire [0:0] cby_1__1__54_left_grid_pin_19_;
wire [0:0] cby_1__1__54_left_grid_pin_20_;
wire [0:0] cby_1__1__54_left_grid_pin_21_;
wire [0:0] cby_1__1__54_left_grid_pin_22_;
wire [0:0] cby_1__1__54_left_grid_pin_23_;
wire [0:0] cby_1__1__54_left_grid_pin_24_;
wire [0:0] cby_1__1__54_left_grid_pin_25_;
wire [0:0] cby_1__1__54_left_grid_pin_26_;
wire [0:0] cby_1__1__54_left_grid_pin_27_;
wire [0:0] cby_1__1__54_left_grid_pin_28_;
wire [0:0] cby_1__1__54_left_grid_pin_29_;
wire [0:0] cby_1__1__54_left_grid_pin_30_;
wire [0:0] cby_1__1__54_left_grid_pin_31_;
wire [0:0] cby_1__1__55_ccff_tail;
wire [0:19] cby_1__1__55_chany_bottom_out;
wire [0:19] cby_1__1__55_chany_top_out;
wire [0:0] cby_1__1__55_left_grid_pin_16_;
wire [0:0] cby_1__1__55_left_grid_pin_17_;
wire [0:0] cby_1__1__55_left_grid_pin_18_;
wire [0:0] cby_1__1__55_left_grid_pin_19_;
wire [0:0] cby_1__1__55_left_grid_pin_20_;
wire [0:0] cby_1__1__55_left_grid_pin_21_;
wire [0:0] cby_1__1__55_left_grid_pin_22_;
wire [0:0] cby_1__1__55_left_grid_pin_23_;
wire [0:0] cby_1__1__55_left_grid_pin_24_;
wire [0:0] cby_1__1__55_left_grid_pin_25_;
wire [0:0] cby_1__1__55_left_grid_pin_26_;
wire [0:0] cby_1__1__55_left_grid_pin_27_;
wire [0:0] cby_1__1__55_left_grid_pin_28_;
wire [0:0] cby_1__1__55_left_grid_pin_29_;
wire [0:0] cby_1__1__55_left_grid_pin_30_;
wire [0:0] cby_1__1__55_left_grid_pin_31_;
wire [0:0] cby_1__1__5_ccff_tail;
wire [0:19] cby_1__1__5_chany_bottom_out;
wire [0:19] cby_1__1__5_chany_top_out;
wire [0:0] cby_1__1__5_left_grid_pin_16_;
wire [0:0] cby_1__1__5_left_grid_pin_17_;
wire [0:0] cby_1__1__5_left_grid_pin_18_;
wire [0:0] cby_1__1__5_left_grid_pin_19_;
wire [0:0] cby_1__1__5_left_grid_pin_20_;
wire [0:0] cby_1__1__5_left_grid_pin_21_;
wire [0:0] cby_1__1__5_left_grid_pin_22_;
wire [0:0] cby_1__1__5_left_grid_pin_23_;
wire [0:0] cby_1__1__5_left_grid_pin_24_;
wire [0:0] cby_1__1__5_left_grid_pin_25_;
wire [0:0] cby_1__1__5_left_grid_pin_26_;
wire [0:0] cby_1__1__5_left_grid_pin_27_;
wire [0:0] cby_1__1__5_left_grid_pin_28_;
wire [0:0] cby_1__1__5_left_grid_pin_29_;
wire [0:0] cby_1__1__5_left_grid_pin_30_;
wire [0:0] cby_1__1__5_left_grid_pin_31_;
wire [0:0] cby_1__1__6_ccff_tail;
wire [0:19] cby_1__1__6_chany_bottom_out;
wire [0:19] cby_1__1__6_chany_top_out;
wire [0:0] cby_1__1__6_left_grid_pin_16_;
wire [0:0] cby_1__1__6_left_grid_pin_17_;
wire [0:0] cby_1__1__6_left_grid_pin_18_;
wire [0:0] cby_1__1__6_left_grid_pin_19_;
wire [0:0] cby_1__1__6_left_grid_pin_20_;
wire [0:0] cby_1__1__6_left_grid_pin_21_;
wire [0:0] cby_1__1__6_left_grid_pin_22_;
wire [0:0] cby_1__1__6_left_grid_pin_23_;
wire [0:0] cby_1__1__6_left_grid_pin_24_;
wire [0:0] cby_1__1__6_left_grid_pin_25_;
wire [0:0] cby_1__1__6_left_grid_pin_26_;
wire [0:0] cby_1__1__6_left_grid_pin_27_;
wire [0:0] cby_1__1__6_left_grid_pin_28_;
wire [0:0] cby_1__1__6_left_grid_pin_29_;
wire [0:0] cby_1__1__6_left_grid_pin_30_;
wire [0:0] cby_1__1__6_left_grid_pin_31_;
wire [0:0] cby_1__1__7_ccff_tail;
wire [0:19] cby_1__1__7_chany_bottom_out;
wire [0:19] cby_1__1__7_chany_top_out;
wire [0:0] cby_1__1__7_left_grid_pin_16_;
wire [0:0] cby_1__1__7_left_grid_pin_17_;
wire [0:0] cby_1__1__7_left_grid_pin_18_;
wire [0:0] cby_1__1__7_left_grid_pin_19_;
wire [0:0] cby_1__1__7_left_grid_pin_20_;
wire [0:0] cby_1__1__7_left_grid_pin_21_;
wire [0:0] cby_1__1__7_left_grid_pin_22_;
wire [0:0] cby_1__1__7_left_grid_pin_23_;
wire [0:0] cby_1__1__7_left_grid_pin_24_;
wire [0:0] cby_1__1__7_left_grid_pin_25_;
wire [0:0] cby_1__1__7_left_grid_pin_26_;
wire [0:0] cby_1__1__7_left_grid_pin_27_;
wire [0:0] cby_1__1__7_left_grid_pin_28_;
wire [0:0] cby_1__1__7_left_grid_pin_29_;
wire [0:0] cby_1__1__7_left_grid_pin_30_;
wire [0:0] cby_1__1__7_left_grid_pin_31_;
wire [0:0] cby_1__1__8_ccff_tail;
wire [0:19] cby_1__1__8_chany_bottom_out;
wire [0:19] cby_1__1__8_chany_top_out;
wire [0:0] cby_1__1__8_left_grid_pin_16_;
wire [0:0] cby_1__1__8_left_grid_pin_17_;
wire [0:0] cby_1__1__8_left_grid_pin_18_;
wire [0:0] cby_1__1__8_left_grid_pin_19_;
wire [0:0] cby_1__1__8_left_grid_pin_20_;
wire [0:0] cby_1__1__8_left_grid_pin_21_;
wire [0:0] cby_1__1__8_left_grid_pin_22_;
wire [0:0] cby_1__1__8_left_grid_pin_23_;
wire [0:0] cby_1__1__8_left_grid_pin_24_;
wire [0:0] cby_1__1__8_left_grid_pin_25_;
wire [0:0] cby_1__1__8_left_grid_pin_26_;
wire [0:0] cby_1__1__8_left_grid_pin_27_;
wire [0:0] cby_1__1__8_left_grid_pin_28_;
wire [0:0] cby_1__1__8_left_grid_pin_29_;
wire [0:0] cby_1__1__8_left_grid_pin_30_;
wire [0:0] cby_1__1__8_left_grid_pin_31_;
wire [0:0] cby_1__1__9_ccff_tail;
wire [0:19] cby_1__1__9_chany_bottom_out;
wire [0:19] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__1__9_left_grid_pin_16_;
wire [0:0] cby_1__1__9_left_grid_pin_17_;
wire [0:0] cby_1__1__9_left_grid_pin_18_;
wire [0:0] cby_1__1__9_left_grid_pin_19_;
wire [0:0] cby_1__1__9_left_grid_pin_20_;
wire [0:0] cby_1__1__9_left_grid_pin_21_;
wire [0:0] cby_1__1__9_left_grid_pin_22_;
wire [0:0] cby_1__1__9_left_grid_pin_23_;
wire [0:0] cby_1__1__9_left_grid_pin_24_;
wire [0:0] cby_1__1__9_left_grid_pin_25_;
wire [0:0] cby_1__1__9_left_grid_pin_26_;
wire [0:0] cby_1__1__9_left_grid_pin_27_;
wire [0:0] cby_1__1__9_left_grid_pin_28_;
wire [0:0] cby_1__1__9_left_grid_pin_29_;
wire [0:0] cby_1__1__9_left_grid_pin_30_;
wire [0:0] cby_1__1__9_left_grid_pin_31_;
wire [0:0] cby_8__1__0_ccff_tail;
wire [0:19] cby_8__1__0_chany_bottom_out;
wire [0:19] cby_8__1__0_chany_top_out;
wire [0:0] cby_8__1__0_left_grid_pin_16_;
wire [0:0] cby_8__1__0_left_grid_pin_17_;
wire [0:0] cby_8__1__0_left_grid_pin_18_;
wire [0:0] cby_8__1__0_left_grid_pin_19_;
wire [0:0] cby_8__1__0_left_grid_pin_20_;
wire [0:0] cby_8__1__0_left_grid_pin_21_;
wire [0:0] cby_8__1__0_left_grid_pin_22_;
wire [0:0] cby_8__1__0_left_grid_pin_23_;
wire [0:0] cby_8__1__0_left_grid_pin_24_;
wire [0:0] cby_8__1__0_left_grid_pin_25_;
wire [0:0] cby_8__1__0_left_grid_pin_26_;
wire [0:0] cby_8__1__0_left_grid_pin_27_;
wire [0:0] cby_8__1__0_left_grid_pin_28_;
wire [0:0] cby_8__1__0_left_grid_pin_29_;
wire [0:0] cby_8__1__0_left_grid_pin_30_;
wire [0:0] cby_8__1__0_left_grid_pin_31_;
wire [0:0] cby_8__1__0_right_grid_pin_0_;
wire [0:0] cby_8__1__1_ccff_tail;
wire [0:19] cby_8__1__1_chany_bottom_out;
wire [0:19] cby_8__1__1_chany_top_out;
wire [0:0] cby_8__1__1_left_grid_pin_16_;
wire [0:0] cby_8__1__1_left_grid_pin_17_;
wire [0:0] cby_8__1__1_left_grid_pin_18_;
wire [0:0] cby_8__1__1_left_grid_pin_19_;
wire [0:0] cby_8__1__1_left_grid_pin_20_;
wire [0:0] cby_8__1__1_left_grid_pin_21_;
wire [0:0] cby_8__1__1_left_grid_pin_22_;
wire [0:0] cby_8__1__1_left_grid_pin_23_;
wire [0:0] cby_8__1__1_left_grid_pin_24_;
wire [0:0] cby_8__1__1_left_grid_pin_25_;
wire [0:0] cby_8__1__1_left_grid_pin_26_;
wire [0:0] cby_8__1__1_left_grid_pin_27_;
wire [0:0] cby_8__1__1_left_grid_pin_28_;
wire [0:0] cby_8__1__1_left_grid_pin_29_;
wire [0:0] cby_8__1__1_left_grid_pin_30_;
wire [0:0] cby_8__1__1_left_grid_pin_31_;
wire [0:0] cby_8__1__1_right_grid_pin_0_;
wire [0:0] cby_8__1__2_ccff_tail;
wire [0:19] cby_8__1__2_chany_bottom_out;
wire [0:19] cby_8__1__2_chany_top_out;
wire [0:0] cby_8__1__2_left_grid_pin_16_;
wire [0:0] cby_8__1__2_left_grid_pin_17_;
wire [0:0] cby_8__1__2_left_grid_pin_18_;
wire [0:0] cby_8__1__2_left_grid_pin_19_;
wire [0:0] cby_8__1__2_left_grid_pin_20_;
wire [0:0] cby_8__1__2_left_grid_pin_21_;
wire [0:0] cby_8__1__2_left_grid_pin_22_;
wire [0:0] cby_8__1__2_left_grid_pin_23_;
wire [0:0] cby_8__1__2_left_grid_pin_24_;
wire [0:0] cby_8__1__2_left_grid_pin_25_;
wire [0:0] cby_8__1__2_left_grid_pin_26_;
wire [0:0] cby_8__1__2_left_grid_pin_27_;
wire [0:0] cby_8__1__2_left_grid_pin_28_;
wire [0:0] cby_8__1__2_left_grid_pin_29_;
wire [0:0] cby_8__1__2_left_grid_pin_30_;
wire [0:0] cby_8__1__2_left_grid_pin_31_;
wire [0:0] cby_8__1__2_right_grid_pin_0_;
wire [0:0] cby_8__1__3_ccff_tail;
wire [0:19] cby_8__1__3_chany_bottom_out;
wire [0:19] cby_8__1__3_chany_top_out;
wire [0:0] cby_8__1__3_left_grid_pin_16_;
wire [0:0] cby_8__1__3_left_grid_pin_17_;
wire [0:0] cby_8__1__3_left_grid_pin_18_;
wire [0:0] cby_8__1__3_left_grid_pin_19_;
wire [0:0] cby_8__1__3_left_grid_pin_20_;
wire [0:0] cby_8__1__3_left_grid_pin_21_;
wire [0:0] cby_8__1__3_left_grid_pin_22_;
wire [0:0] cby_8__1__3_left_grid_pin_23_;
wire [0:0] cby_8__1__3_left_grid_pin_24_;
wire [0:0] cby_8__1__3_left_grid_pin_25_;
wire [0:0] cby_8__1__3_left_grid_pin_26_;
wire [0:0] cby_8__1__3_left_grid_pin_27_;
wire [0:0] cby_8__1__3_left_grid_pin_28_;
wire [0:0] cby_8__1__3_left_grid_pin_29_;
wire [0:0] cby_8__1__3_left_grid_pin_30_;
wire [0:0] cby_8__1__3_left_grid_pin_31_;
wire [0:0] cby_8__1__3_right_grid_pin_0_;
wire [0:0] cby_8__1__4_ccff_tail;
wire [0:19] cby_8__1__4_chany_bottom_out;
wire [0:19] cby_8__1__4_chany_top_out;
wire [0:0] cby_8__1__4_left_grid_pin_16_;
wire [0:0] cby_8__1__4_left_grid_pin_17_;
wire [0:0] cby_8__1__4_left_grid_pin_18_;
wire [0:0] cby_8__1__4_left_grid_pin_19_;
wire [0:0] cby_8__1__4_left_grid_pin_20_;
wire [0:0] cby_8__1__4_left_grid_pin_21_;
wire [0:0] cby_8__1__4_left_grid_pin_22_;
wire [0:0] cby_8__1__4_left_grid_pin_23_;
wire [0:0] cby_8__1__4_left_grid_pin_24_;
wire [0:0] cby_8__1__4_left_grid_pin_25_;
wire [0:0] cby_8__1__4_left_grid_pin_26_;
wire [0:0] cby_8__1__4_left_grid_pin_27_;
wire [0:0] cby_8__1__4_left_grid_pin_28_;
wire [0:0] cby_8__1__4_left_grid_pin_29_;
wire [0:0] cby_8__1__4_left_grid_pin_30_;
wire [0:0] cby_8__1__4_left_grid_pin_31_;
wire [0:0] cby_8__1__4_right_grid_pin_0_;
wire [0:0] cby_8__1__5_ccff_tail;
wire [0:19] cby_8__1__5_chany_bottom_out;
wire [0:19] cby_8__1__5_chany_top_out;
wire [0:0] cby_8__1__5_left_grid_pin_16_;
wire [0:0] cby_8__1__5_left_grid_pin_17_;
wire [0:0] cby_8__1__5_left_grid_pin_18_;
wire [0:0] cby_8__1__5_left_grid_pin_19_;
wire [0:0] cby_8__1__5_left_grid_pin_20_;
wire [0:0] cby_8__1__5_left_grid_pin_21_;
wire [0:0] cby_8__1__5_left_grid_pin_22_;
wire [0:0] cby_8__1__5_left_grid_pin_23_;
wire [0:0] cby_8__1__5_left_grid_pin_24_;
wire [0:0] cby_8__1__5_left_grid_pin_25_;
wire [0:0] cby_8__1__5_left_grid_pin_26_;
wire [0:0] cby_8__1__5_left_grid_pin_27_;
wire [0:0] cby_8__1__5_left_grid_pin_28_;
wire [0:0] cby_8__1__5_left_grid_pin_29_;
wire [0:0] cby_8__1__5_left_grid_pin_30_;
wire [0:0] cby_8__1__5_left_grid_pin_31_;
wire [0:0] cby_8__1__5_right_grid_pin_0_;
wire [0:0] cby_8__1__6_ccff_tail;
wire [0:19] cby_8__1__6_chany_bottom_out;
wire [0:19] cby_8__1__6_chany_top_out;
wire [0:0] cby_8__1__6_left_grid_pin_16_;
wire [0:0] cby_8__1__6_left_grid_pin_17_;
wire [0:0] cby_8__1__6_left_grid_pin_18_;
wire [0:0] cby_8__1__6_left_grid_pin_19_;
wire [0:0] cby_8__1__6_left_grid_pin_20_;
wire [0:0] cby_8__1__6_left_grid_pin_21_;
wire [0:0] cby_8__1__6_left_grid_pin_22_;
wire [0:0] cby_8__1__6_left_grid_pin_23_;
wire [0:0] cby_8__1__6_left_grid_pin_24_;
wire [0:0] cby_8__1__6_left_grid_pin_25_;
wire [0:0] cby_8__1__6_left_grid_pin_26_;
wire [0:0] cby_8__1__6_left_grid_pin_27_;
wire [0:0] cby_8__1__6_left_grid_pin_28_;
wire [0:0] cby_8__1__6_left_grid_pin_29_;
wire [0:0] cby_8__1__6_left_grid_pin_30_;
wire [0:0] cby_8__1__6_left_grid_pin_31_;
wire [0:0] cby_8__1__6_right_grid_pin_0_;
wire [0:0] cby_8__1__7_ccff_tail;
wire [0:19] cby_8__1__7_chany_bottom_out;
wire [0:19] cby_8__1__7_chany_top_out;
wire [0:0] cby_8__1__7_left_grid_pin_16_;
wire [0:0] cby_8__1__7_left_grid_pin_17_;
wire [0:0] cby_8__1__7_left_grid_pin_18_;
wire [0:0] cby_8__1__7_left_grid_pin_19_;
wire [0:0] cby_8__1__7_left_grid_pin_20_;
wire [0:0] cby_8__1__7_left_grid_pin_21_;
wire [0:0] cby_8__1__7_left_grid_pin_22_;
wire [0:0] cby_8__1__7_left_grid_pin_23_;
wire [0:0] cby_8__1__7_left_grid_pin_24_;
wire [0:0] cby_8__1__7_left_grid_pin_25_;
wire [0:0] cby_8__1__7_left_grid_pin_26_;
wire [0:0] cby_8__1__7_left_grid_pin_27_;
wire [0:0] cby_8__1__7_left_grid_pin_28_;
wire [0:0] cby_8__1__7_left_grid_pin_29_;
wire [0:0] cby_8__1__7_left_grid_pin_30_;
wire [0:0] cby_8__1__7_left_grid_pin_31_;
wire [0:0] cby_8__1__7_right_grid_pin_0_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_100_out;
wire [0:0] direct_interc_101_out;
wire [0:0] direct_interc_102_out;
wire [0:0] direct_interc_103_out;
wire [0:0] direct_interc_104_out;
wire [0:0] direct_interc_105_out;
wire [0:0] direct_interc_106_out;
wire [0:0] direct_interc_107_out;
wire [0:0] direct_interc_108_out;
wire [0:0] direct_interc_109_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_110_out;
wire [0:0] direct_interc_111_out;
wire [0:0] direct_interc_112_out;
wire [0:0] direct_interc_113_out;
wire [0:0] direct_interc_114_out;
wire [0:0] direct_interc_115_out;
wire [0:0] direct_interc_116_out;
wire [0:0] direct_interc_117_out;
wire [0:0] direct_interc_118_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_44_out;
wire [0:0] direct_interc_45_out;
wire [0:0] direct_interc_46_out;
wire [0:0] direct_interc_47_out;
wire [0:0] direct_interc_48_out;
wire [0:0] direct_interc_49_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_50_out;
wire [0:0] direct_interc_51_out;
wire [0:0] direct_interc_52_out;
wire [0:0] direct_interc_53_out;
wire [0:0] direct_interc_54_out;
wire [0:0] direct_interc_55_out;
wire [0:0] direct_interc_56_out;
wire [0:0] direct_interc_57_out;
wire [0:0] direct_interc_58_out;
wire [0:0] direct_interc_59_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_60_out;
wire [0:0] direct_interc_61_out;
wire [0:0] direct_interc_62_out;
wire [0:0] direct_interc_63_out;
wire [0:0] direct_interc_64_out;
wire [0:0] direct_interc_65_out;
wire [0:0] direct_interc_66_out;
wire [0:0] direct_interc_67_out;
wire [0:0] direct_interc_68_out;
wire [0:0] direct_interc_69_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_70_out;
wire [0:0] direct_interc_71_out;
wire [0:0] direct_interc_72_out;
wire [0:0] direct_interc_73_out;
wire [0:0] direct_interc_74_out;
wire [0:0] direct_interc_75_out;
wire [0:0] direct_interc_76_out;
wire [0:0] direct_interc_77_out;
wire [0:0] direct_interc_78_out;
wire [0:0] direct_interc_79_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_80_out;
wire [0:0] direct_interc_81_out;
wire [0:0] direct_interc_82_out;
wire [0:0] direct_interc_83_out;
wire [0:0] direct_interc_84_out;
wire [0:0] direct_interc_85_out;
wire [0:0] direct_interc_86_out;
wire [0:0] direct_interc_87_out;
wire [0:0] direct_interc_88_out;
wire [0:0] direct_interc_89_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_90_out;
wire [0:0] direct_interc_91_out;
wire [0:0] direct_interc_92_out;
wire [0:0] direct_interc_93_out;
wire [0:0] direct_interc_94_out;
wire [0:0] direct_interc_95_out;
wire [0:0] direct_interc_96_out;
wire [0:0] direct_interc_97_out;
wire [0:0] direct_interc_98_out;
wire [0:0] direct_interc_99_out;
wire [0:0] direct_interc_9_out;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_1__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_1__8__undriven_top_width_0_height_0__pin_33_;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_22_ccff_tail;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_23_ccff_tail;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_24_ccff_tail;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_25_ccff_tail;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_26_ccff_tail;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_27_ccff_tail;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_28_ccff_tail;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_29_ccff_tail;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_2__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_30_ccff_tail;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_31_ccff_tail;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_32_ccff_tail;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_33_ccff_tail;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_34_ccff_tail;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_35_ccff_tail;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_36_ccff_tail;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_37_ccff_tail;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_38_ccff_tail;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_39_ccff_tail;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_3__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_40_ccff_tail;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_41_ccff_tail;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_42_ccff_tail;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_43_ccff_tail;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_44_ccff_tail;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_45_ccff_tail;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_46_ccff_tail;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_47_ccff_tail;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_48_ccff_tail;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_49_ccff_tail;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_4__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_50_ccff_tail;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_51_ccff_tail;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_52_ccff_tail;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_53_ccff_tail;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_54_ccff_tail;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_55_ccff_tail;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_56_ccff_tail;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_57_ccff_tail;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_58_ccff_tail;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_59_ccff_tail;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_5__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_60_ccff_tail;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_61_ccff_tail;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_62_ccff_tail;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_63_ccff_tail;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_6__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_7__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_8__8__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_upper;
wire [0:0] grid_io_bottom_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_6_ccff_tail;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_bottom_bottom_7_ccff_tail;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_upper;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_lower;
wire [0:0] grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_upper;
wire [0:0] grid_io_left_left_0_ccff_tail;
wire [0:0] grid_io_left_left_0_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_0_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_1_ccff_tail;
wire [0:0] grid_io_left_left_1_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_1_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_2_ccff_tail;
wire [0:0] grid_io_left_left_2_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_2_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_3_ccff_tail;
wire [0:0] grid_io_left_left_3_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_3_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_4_ccff_tail;
wire [0:0] grid_io_left_left_4_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_4_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_5_ccff_tail;
wire [0:0] grid_io_left_left_5_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_5_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_6_ccff_tail;
wire [0:0] grid_io_left_left_6_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_6_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_left_7_ccff_tail;
wire [0:0] grid_io_left_left_7_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_left_7_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_0_ccff_tail;
wire [0:0] grid_io_right_right_0_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_0_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_1_ccff_tail;
wire [0:0] grid_io_right_right_1_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_1_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_2_ccff_tail;
wire [0:0] grid_io_right_right_2_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_2_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_3_ccff_tail;
wire [0:0] grid_io_right_right_3_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_3_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_4_ccff_tail;
wire [0:0] grid_io_right_right_4_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_4_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_5_ccff_tail;
wire [0:0] grid_io_right_right_5_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_5_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_6_ccff_tail;
wire [0:0] grid_io_right_right_6_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_6_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_right_7_ccff_tail;
wire [0:0] grid_io_right_right_7_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_right_7_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_0_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_0_ccff_tail;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_1_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_1_ccff_tail;
wire [0:0] grid_io_top_top_2_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_2_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_2_ccff_tail;
wire [0:0] grid_io_top_top_3_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_3_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_3_ccff_tail;
wire [0:0] grid_io_top_top_4_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_4_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_4_ccff_tail;
wire [0:0] grid_io_top_top_5_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_5_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_5_ccff_tail;
wire [0:0] grid_io_top_top_6_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_6_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_6_ccff_tail;
wire [0:0] grid_io_top_top_7_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_top_7_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_top_7_ccff_tail;
wire [0:19] sb_0__0__0_chanx_right_out;
wire [0:19] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:19] sb_0__1__0_chanx_right_out;
wire [0:19] sb_0__1__0_chany_bottom_out;
wire [0:19] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:19] sb_0__1__1_chanx_right_out;
wire [0:19] sb_0__1__1_chany_bottom_out;
wire [0:19] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__1__2_ccff_tail;
wire [0:19] sb_0__1__2_chanx_right_out;
wire [0:19] sb_0__1__2_chany_bottom_out;
wire [0:19] sb_0__1__2_chany_top_out;
wire [0:0] sb_0__1__3_ccff_tail;
wire [0:19] sb_0__1__3_chanx_right_out;
wire [0:19] sb_0__1__3_chany_bottom_out;
wire [0:19] sb_0__1__3_chany_top_out;
wire [0:0] sb_0__1__4_ccff_tail;
wire [0:19] sb_0__1__4_chanx_right_out;
wire [0:19] sb_0__1__4_chany_bottom_out;
wire [0:19] sb_0__1__4_chany_top_out;
wire [0:0] sb_0__1__5_ccff_tail;
wire [0:19] sb_0__1__5_chanx_right_out;
wire [0:19] sb_0__1__5_chany_bottom_out;
wire [0:19] sb_0__1__5_chany_top_out;
wire [0:0] sb_0__1__6_ccff_tail;
wire [0:19] sb_0__1__6_chanx_right_out;
wire [0:19] sb_0__1__6_chany_bottom_out;
wire [0:19] sb_0__1__6_chany_top_out;
wire [0:0] sb_0__8__0_ccff_tail;
wire [0:19] sb_0__8__0_chanx_right_out;
wire [0:19] sb_0__8__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:19] sb_1__0__0_chanx_left_out;
wire [0:19] sb_1__0__0_chanx_right_out;
wire [0:19] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:19] sb_1__0__1_chanx_left_out;
wire [0:19] sb_1__0__1_chanx_right_out;
wire [0:19] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:19] sb_1__0__2_chanx_left_out;
wire [0:19] sb_1__0__2_chanx_right_out;
wire [0:19] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:19] sb_1__0__3_chanx_left_out;
wire [0:19] sb_1__0__3_chanx_right_out;
wire [0:19] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:19] sb_1__0__4_chanx_left_out;
wire [0:19] sb_1__0__4_chanx_right_out;
wire [0:19] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__0__5_ccff_tail;
wire [0:19] sb_1__0__5_chanx_left_out;
wire [0:19] sb_1__0__5_chanx_right_out;
wire [0:19] sb_1__0__5_chany_top_out;
wire [0:0] sb_1__0__6_ccff_tail;
wire [0:19] sb_1__0__6_chanx_left_out;
wire [0:19] sb_1__0__6_chanx_right_out;
wire [0:19] sb_1__0__6_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:19] sb_1__1__0_chanx_left_out;
wire [0:19] sb_1__1__0_chanx_right_out;
wire [0:19] sb_1__1__0_chany_bottom_out;
wire [0:19] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__10_ccff_tail;
wire [0:19] sb_1__1__10_chanx_left_out;
wire [0:19] sb_1__1__10_chanx_right_out;
wire [0:19] sb_1__1__10_chany_bottom_out;
wire [0:19] sb_1__1__10_chany_top_out;
wire [0:0] sb_1__1__11_ccff_tail;
wire [0:19] sb_1__1__11_chanx_left_out;
wire [0:19] sb_1__1__11_chanx_right_out;
wire [0:19] sb_1__1__11_chany_bottom_out;
wire [0:19] sb_1__1__11_chany_top_out;
wire [0:0] sb_1__1__12_ccff_tail;
wire [0:19] sb_1__1__12_chanx_left_out;
wire [0:19] sb_1__1__12_chanx_right_out;
wire [0:19] sb_1__1__12_chany_bottom_out;
wire [0:19] sb_1__1__12_chany_top_out;
wire [0:0] sb_1__1__13_ccff_tail;
wire [0:19] sb_1__1__13_chanx_left_out;
wire [0:19] sb_1__1__13_chanx_right_out;
wire [0:19] sb_1__1__13_chany_bottom_out;
wire [0:19] sb_1__1__13_chany_top_out;
wire [0:0] sb_1__1__14_ccff_tail;
wire [0:19] sb_1__1__14_chanx_left_out;
wire [0:19] sb_1__1__14_chanx_right_out;
wire [0:19] sb_1__1__14_chany_bottom_out;
wire [0:19] sb_1__1__14_chany_top_out;
wire [0:0] sb_1__1__15_ccff_tail;
wire [0:19] sb_1__1__15_chanx_left_out;
wire [0:19] sb_1__1__15_chanx_right_out;
wire [0:19] sb_1__1__15_chany_bottom_out;
wire [0:19] sb_1__1__15_chany_top_out;
wire [0:0] sb_1__1__16_ccff_tail;
wire [0:19] sb_1__1__16_chanx_left_out;
wire [0:19] sb_1__1__16_chanx_right_out;
wire [0:19] sb_1__1__16_chany_bottom_out;
wire [0:19] sb_1__1__16_chany_top_out;
wire [0:0] sb_1__1__17_ccff_tail;
wire [0:19] sb_1__1__17_chanx_left_out;
wire [0:19] sb_1__1__17_chanx_right_out;
wire [0:19] sb_1__1__17_chany_bottom_out;
wire [0:19] sb_1__1__17_chany_top_out;
wire [0:0] sb_1__1__18_ccff_tail;
wire [0:19] sb_1__1__18_chanx_left_out;
wire [0:19] sb_1__1__18_chanx_right_out;
wire [0:19] sb_1__1__18_chany_bottom_out;
wire [0:19] sb_1__1__18_chany_top_out;
wire [0:0] sb_1__1__19_ccff_tail;
wire [0:19] sb_1__1__19_chanx_left_out;
wire [0:19] sb_1__1__19_chanx_right_out;
wire [0:19] sb_1__1__19_chany_bottom_out;
wire [0:19] sb_1__1__19_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:19] sb_1__1__1_chanx_left_out;
wire [0:19] sb_1__1__1_chanx_right_out;
wire [0:19] sb_1__1__1_chany_bottom_out;
wire [0:19] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__20_ccff_tail;
wire [0:19] sb_1__1__20_chanx_left_out;
wire [0:19] sb_1__1__20_chanx_right_out;
wire [0:19] sb_1__1__20_chany_bottom_out;
wire [0:19] sb_1__1__20_chany_top_out;
wire [0:0] sb_1__1__21_ccff_tail;
wire [0:19] sb_1__1__21_chanx_left_out;
wire [0:19] sb_1__1__21_chanx_right_out;
wire [0:19] sb_1__1__21_chany_bottom_out;
wire [0:19] sb_1__1__21_chany_top_out;
wire [0:0] sb_1__1__22_ccff_tail;
wire [0:19] sb_1__1__22_chanx_left_out;
wire [0:19] sb_1__1__22_chanx_right_out;
wire [0:19] sb_1__1__22_chany_bottom_out;
wire [0:19] sb_1__1__22_chany_top_out;
wire [0:0] sb_1__1__23_ccff_tail;
wire [0:19] sb_1__1__23_chanx_left_out;
wire [0:19] sb_1__1__23_chanx_right_out;
wire [0:19] sb_1__1__23_chany_bottom_out;
wire [0:19] sb_1__1__23_chany_top_out;
wire [0:0] sb_1__1__24_ccff_tail;
wire [0:19] sb_1__1__24_chanx_left_out;
wire [0:19] sb_1__1__24_chanx_right_out;
wire [0:19] sb_1__1__24_chany_bottom_out;
wire [0:19] sb_1__1__24_chany_top_out;
wire [0:0] sb_1__1__25_ccff_tail;
wire [0:19] sb_1__1__25_chanx_left_out;
wire [0:19] sb_1__1__25_chanx_right_out;
wire [0:19] sb_1__1__25_chany_bottom_out;
wire [0:19] sb_1__1__25_chany_top_out;
wire [0:0] sb_1__1__26_ccff_tail;
wire [0:19] sb_1__1__26_chanx_left_out;
wire [0:19] sb_1__1__26_chanx_right_out;
wire [0:19] sb_1__1__26_chany_bottom_out;
wire [0:19] sb_1__1__26_chany_top_out;
wire [0:0] sb_1__1__27_ccff_tail;
wire [0:19] sb_1__1__27_chanx_left_out;
wire [0:19] sb_1__1__27_chanx_right_out;
wire [0:19] sb_1__1__27_chany_bottom_out;
wire [0:19] sb_1__1__27_chany_top_out;
wire [0:0] sb_1__1__28_ccff_tail;
wire [0:19] sb_1__1__28_chanx_left_out;
wire [0:19] sb_1__1__28_chanx_right_out;
wire [0:19] sb_1__1__28_chany_bottom_out;
wire [0:19] sb_1__1__28_chany_top_out;
wire [0:0] sb_1__1__29_ccff_tail;
wire [0:19] sb_1__1__29_chanx_left_out;
wire [0:19] sb_1__1__29_chanx_right_out;
wire [0:19] sb_1__1__29_chany_bottom_out;
wire [0:19] sb_1__1__29_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:19] sb_1__1__2_chanx_left_out;
wire [0:19] sb_1__1__2_chanx_right_out;
wire [0:19] sb_1__1__2_chany_bottom_out;
wire [0:19] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__30_ccff_tail;
wire [0:19] sb_1__1__30_chanx_left_out;
wire [0:19] sb_1__1__30_chanx_right_out;
wire [0:19] sb_1__1__30_chany_bottom_out;
wire [0:19] sb_1__1__30_chany_top_out;
wire [0:0] sb_1__1__31_ccff_tail;
wire [0:19] sb_1__1__31_chanx_left_out;
wire [0:19] sb_1__1__31_chanx_right_out;
wire [0:19] sb_1__1__31_chany_bottom_out;
wire [0:19] sb_1__1__31_chany_top_out;
wire [0:0] sb_1__1__32_ccff_tail;
wire [0:19] sb_1__1__32_chanx_left_out;
wire [0:19] sb_1__1__32_chanx_right_out;
wire [0:19] sb_1__1__32_chany_bottom_out;
wire [0:19] sb_1__1__32_chany_top_out;
wire [0:0] sb_1__1__33_ccff_tail;
wire [0:19] sb_1__1__33_chanx_left_out;
wire [0:19] sb_1__1__33_chanx_right_out;
wire [0:19] sb_1__1__33_chany_bottom_out;
wire [0:19] sb_1__1__33_chany_top_out;
wire [0:0] sb_1__1__34_ccff_tail;
wire [0:19] sb_1__1__34_chanx_left_out;
wire [0:19] sb_1__1__34_chanx_right_out;
wire [0:19] sb_1__1__34_chany_bottom_out;
wire [0:19] sb_1__1__34_chany_top_out;
wire [0:0] sb_1__1__35_ccff_tail;
wire [0:19] sb_1__1__35_chanx_left_out;
wire [0:19] sb_1__1__35_chanx_right_out;
wire [0:19] sb_1__1__35_chany_bottom_out;
wire [0:19] sb_1__1__35_chany_top_out;
wire [0:0] sb_1__1__36_ccff_tail;
wire [0:19] sb_1__1__36_chanx_left_out;
wire [0:19] sb_1__1__36_chanx_right_out;
wire [0:19] sb_1__1__36_chany_bottom_out;
wire [0:19] sb_1__1__36_chany_top_out;
wire [0:0] sb_1__1__37_ccff_tail;
wire [0:19] sb_1__1__37_chanx_left_out;
wire [0:19] sb_1__1__37_chanx_right_out;
wire [0:19] sb_1__1__37_chany_bottom_out;
wire [0:19] sb_1__1__37_chany_top_out;
wire [0:0] sb_1__1__38_ccff_tail;
wire [0:19] sb_1__1__38_chanx_left_out;
wire [0:19] sb_1__1__38_chanx_right_out;
wire [0:19] sb_1__1__38_chany_bottom_out;
wire [0:19] sb_1__1__38_chany_top_out;
wire [0:0] sb_1__1__39_ccff_tail;
wire [0:19] sb_1__1__39_chanx_left_out;
wire [0:19] sb_1__1__39_chanx_right_out;
wire [0:19] sb_1__1__39_chany_bottom_out;
wire [0:19] sb_1__1__39_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:19] sb_1__1__3_chanx_left_out;
wire [0:19] sb_1__1__3_chanx_right_out;
wire [0:19] sb_1__1__3_chany_bottom_out;
wire [0:19] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__40_ccff_tail;
wire [0:19] sb_1__1__40_chanx_left_out;
wire [0:19] sb_1__1__40_chanx_right_out;
wire [0:19] sb_1__1__40_chany_bottom_out;
wire [0:19] sb_1__1__40_chany_top_out;
wire [0:0] sb_1__1__41_ccff_tail;
wire [0:19] sb_1__1__41_chanx_left_out;
wire [0:19] sb_1__1__41_chanx_right_out;
wire [0:19] sb_1__1__41_chany_bottom_out;
wire [0:19] sb_1__1__41_chany_top_out;
wire [0:0] sb_1__1__42_ccff_tail;
wire [0:19] sb_1__1__42_chanx_left_out;
wire [0:19] sb_1__1__42_chanx_right_out;
wire [0:19] sb_1__1__42_chany_bottom_out;
wire [0:19] sb_1__1__42_chany_top_out;
wire [0:0] sb_1__1__43_ccff_tail;
wire [0:19] sb_1__1__43_chanx_left_out;
wire [0:19] sb_1__1__43_chanx_right_out;
wire [0:19] sb_1__1__43_chany_bottom_out;
wire [0:19] sb_1__1__43_chany_top_out;
wire [0:0] sb_1__1__44_ccff_tail;
wire [0:19] sb_1__1__44_chanx_left_out;
wire [0:19] sb_1__1__44_chanx_right_out;
wire [0:19] sb_1__1__44_chany_bottom_out;
wire [0:19] sb_1__1__44_chany_top_out;
wire [0:0] sb_1__1__45_ccff_tail;
wire [0:19] sb_1__1__45_chanx_left_out;
wire [0:19] sb_1__1__45_chanx_right_out;
wire [0:19] sb_1__1__45_chany_bottom_out;
wire [0:19] sb_1__1__45_chany_top_out;
wire [0:0] sb_1__1__46_ccff_tail;
wire [0:19] sb_1__1__46_chanx_left_out;
wire [0:19] sb_1__1__46_chanx_right_out;
wire [0:19] sb_1__1__46_chany_bottom_out;
wire [0:19] sb_1__1__46_chany_top_out;
wire [0:0] sb_1__1__47_ccff_tail;
wire [0:19] sb_1__1__47_chanx_left_out;
wire [0:19] sb_1__1__47_chanx_right_out;
wire [0:19] sb_1__1__47_chany_bottom_out;
wire [0:19] sb_1__1__47_chany_top_out;
wire [0:0] sb_1__1__48_ccff_tail;
wire [0:19] sb_1__1__48_chanx_left_out;
wire [0:19] sb_1__1__48_chanx_right_out;
wire [0:19] sb_1__1__48_chany_bottom_out;
wire [0:19] sb_1__1__48_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:19] sb_1__1__4_chanx_left_out;
wire [0:19] sb_1__1__4_chanx_right_out;
wire [0:19] sb_1__1__4_chany_bottom_out;
wire [0:19] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:19] sb_1__1__5_chanx_left_out;
wire [0:19] sb_1__1__5_chanx_right_out;
wire [0:19] sb_1__1__5_chany_bottom_out;
wire [0:19] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:19] sb_1__1__6_chanx_left_out;
wire [0:19] sb_1__1__6_chanx_right_out;
wire [0:19] sb_1__1__6_chany_bottom_out;
wire [0:19] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:19] sb_1__1__7_chanx_left_out;
wire [0:19] sb_1__1__7_chanx_right_out;
wire [0:19] sb_1__1__7_chany_bottom_out;
wire [0:19] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:19] sb_1__1__8_chanx_left_out;
wire [0:19] sb_1__1__8_chanx_right_out;
wire [0:19] sb_1__1__8_chany_bottom_out;
wire [0:19] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__1__9_ccff_tail;
wire [0:19] sb_1__1__9_chanx_left_out;
wire [0:19] sb_1__1__9_chanx_right_out;
wire [0:19] sb_1__1__9_chany_bottom_out;
wire [0:19] sb_1__1__9_chany_top_out;
wire [0:0] sb_1__8__0_ccff_tail;
wire [0:19] sb_1__8__0_chanx_left_out;
wire [0:19] sb_1__8__0_chanx_right_out;
wire [0:19] sb_1__8__0_chany_bottom_out;
wire [0:0] sb_1__8__1_ccff_tail;
wire [0:19] sb_1__8__1_chanx_left_out;
wire [0:19] sb_1__8__1_chanx_right_out;
wire [0:19] sb_1__8__1_chany_bottom_out;
wire [0:0] sb_1__8__2_ccff_tail;
wire [0:19] sb_1__8__2_chanx_left_out;
wire [0:19] sb_1__8__2_chanx_right_out;
wire [0:19] sb_1__8__2_chany_bottom_out;
wire [0:0] sb_1__8__3_ccff_tail;
wire [0:19] sb_1__8__3_chanx_left_out;
wire [0:19] sb_1__8__3_chanx_right_out;
wire [0:19] sb_1__8__3_chany_bottom_out;
wire [0:0] sb_1__8__4_ccff_tail;
wire [0:19] sb_1__8__4_chanx_left_out;
wire [0:19] sb_1__8__4_chanx_right_out;
wire [0:19] sb_1__8__4_chany_bottom_out;
wire [0:0] sb_1__8__5_ccff_tail;
wire [0:19] sb_1__8__5_chanx_left_out;
wire [0:19] sb_1__8__5_chanx_right_out;
wire [0:19] sb_1__8__5_chany_bottom_out;
wire [0:0] sb_1__8__6_ccff_tail;
wire [0:19] sb_1__8__6_chanx_left_out;
wire [0:19] sb_1__8__6_chanx_right_out;
wire [0:19] sb_1__8__6_chany_bottom_out;
wire [0:0] sb_8__0__0_ccff_tail;
wire [0:19] sb_8__0__0_chanx_left_out;
wire [0:19] sb_8__0__0_chany_top_out;
wire [0:0] sb_8__1__0_ccff_tail;
wire [0:19] sb_8__1__0_chanx_left_out;
wire [0:19] sb_8__1__0_chany_bottom_out;
wire [0:19] sb_8__1__0_chany_top_out;
wire [0:0] sb_8__1__1_ccff_tail;
wire [0:19] sb_8__1__1_chanx_left_out;
wire [0:19] sb_8__1__1_chany_bottom_out;
wire [0:19] sb_8__1__1_chany_top_out;
wire [0:0] sb_8__1__2_ccff_tail;
wire [0:19] sb_8__1__2_chanx_left_out;
wire [0:19] sb_8__1__2_chany_bottom_out;
wire [0:19] sb_8__1__2_chany_top_out;
wire [0:0] sb_8__1__3_ccff_tail;
wire [0:19] sb_8__1__3_chanx_left_out;
wire [0:19] sb_8__1__3_chany_bottom_out;
wire [0:19] sb_8__1__3_chany_top_out;
wire [0:0] sb_8__1__4_ccff_tail;
wire [0:19] sb_8__1__4_chanx_left_out;
wire [0:19] sb_8__1__4_chany_bottom_out;
wire [0:19] sb_8__1__4_chany_top_out;
wire [0:0] sb_8__1__5_ccff_tail;
wire [0:19] sb_8__1__5_chanx_left_out;
wire [0:19] sb_8__1__5_chany_bottom_out;
wire [0:19] sb_8__1__5_chany_top_out;
wire [0:0] sb_8__1__6_ccff_tail;
wire [0:19] sb_8__1__6_chanx_left_out;
wire [0:19] sb_8__1__6_chany_bottom_out;
wire [0:19] sb_8__1__6_chany_top_out;
wire [0:0] sb_8__8__0_ccff_tail;
wire [0:19] sb_8__8__0_chanx_left_out;
wire [0:19] sb_8__8__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_0_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_56_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_0_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_0_ccff_tail[0]));

	grid_clb grid_clb_1__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_1_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_57_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_1_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_1_ccff_tail[0]));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_2_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_58_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_2_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_2_ccff_tail[0]));

	grid_clb grid_clb_1__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_3_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_59_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_3_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_3_ccff_tail[0]));

	grid_clb grid_clb_1__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_4_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_60_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_4_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_4_ccff_tail[0]));

	grid_clb grid_clb_1__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_5_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_61_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_5_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_5_ccff_tail[0]));

	grid_clb grid_clb_1__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_6_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_62_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_6_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_6_ccff_tail[0]));

	grid_clb grid_clb_1__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__0_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__0_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__0_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__0_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__0_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__0_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__0_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__0_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__0_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__0_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__0_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__0_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__0_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__0_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__0_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__0_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_1__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(grid_clb_1__8__undriven_top_width_0_height_0__pin_33_[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(grid_io_left_left_7_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_7_ccff_tail[0]));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_7_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_63_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__0_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_8_ccff_tail[0]));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_8_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_64_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__1_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_9_ccff_tail[0]));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_9_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_65_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__2_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_10_ccff_tail[0]));

	grid_clb grid_clb_2__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_10_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_66_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__3_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_11_ccff_tail[0]));

	grid_clb grid_clb_2__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_11_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_67_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__4_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_12_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_12_ccff_tail[0]));

	grid_clb grid_clb_2__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_12_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_68_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__5_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_13_ccff_tail[0]));

	grid_clb grid_clb_2__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_13_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_69_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__6_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_14_ccff_tail[0]));

	grid_clb grid_clb_2__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__1_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__1_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__1_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__1_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__1_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__1_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__1_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__1_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__1_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__1_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__1_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__1_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__1_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__1_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__1_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__1_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_2__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_112_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__7_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_15_ccff_tail[0]));

	grid_clb grid_clb_3__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_14_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_70_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__8_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_16_ccff_tail[0]));

	grid_clb grid_clb_3__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_15_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_71_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__9_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_17_ccff_tail[0]));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_16_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_72_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__10_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_18_ccff_tail[0]));

	grid_clb grid_clb_3__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_17_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_73_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__11_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_19_ccff_tail[0]));

	grid_clb grid_clb_3__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_18_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_74_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__12_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_20_ccff_tail[0]));

	grid_clb grid_clb_3__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_19_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_75_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__13_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_21_ccff_tail[0]));

	grid_clb grid_clb_3__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_20_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_76_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__14_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_22_ccff_tail[0]));

	grid_clb grid_clb_3__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__2_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__2_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__2_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__2_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__2_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__2_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__2_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__2_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__2_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__2_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__2_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__2_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__2_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__2_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__2_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__2_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_3__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_113_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__15_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_23_ccff_tail[0]));

	grid_clb grid_clb_4__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_21_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_77_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__16_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_24_ccff_tail[0]));

	grid_clb grid_clb_4__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_22_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_78_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__17_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_25_ccff_tail[0]));

	grid_clb grid_clb_4__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_23_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_79_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__18_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_26_ccff_tail[0]));

	grid_clb grid_clb_4__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_24_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_80_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__19_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_27_ccff_tail[0]));

	grid_clb grid_clb_4__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_25_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_81_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__20_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_28_ccff_tail[0]));

	grid_clb grid_clb_4__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_26_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_82_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__21_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_29_ccff_tail[0]));

	grid_clb grid_clb_4__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_27_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_83_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__22_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_30_ccff_tail[0]));

	grid_clb grid_clb_4__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__3_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__3_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__3_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__3_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__3_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__3_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__3_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__3_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__3_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__3_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__3_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__3_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__3_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__3_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__3_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__3_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_4__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_114_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__23_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_31_ccff_tail[0]));

	grid_clb grid_clb_5__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_28_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_84_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__24_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_32_ccff_tail[0]));

	grid_clb grid_clb_5__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_29_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_85_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__25_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_33_ccff_tail[0]));

	grid_clb grid_clb_5__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_30_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_86_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__26_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_34_ccff_tail[0]));

	grid_clb grid_clb_5__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_31_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_87_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__27_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_35_ccff_tail[0]));

	grid_clb grid_clb_5__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_32_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_88_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__28_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_36_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_36_ccff_tail[0]));

	grid_clb grid_clb_5__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_33_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_89_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__29_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_37_ccff_tail[0]));

	grid_clb grid_clb_5__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_34_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_90_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__30_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_38_ccff_tail[0]));

	grid_clb grid_clb_5__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__4_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__4_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__4_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__4_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__4_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__4_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__4_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__4_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__4_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__4_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__4_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__4_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__4_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__4_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__4_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__4_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_5__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_115_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__31_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_39_ccff_tail[0]));

	grid_clb grid_clb_6__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_35_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_91_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__32_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_40_ccff_tail[0]));

	grid_clb grid_clb_6__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_36_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_92_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__33_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_41_ccff_tail[0]));

	grid_clb grid_clb_6__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_37_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_93_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__34_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_42_ccff_tail[0]));

	grid_clb grid_clb_6__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_38_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_94_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__35_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_43_ccff_tail[0]));

	grid_clb grid_clb_6__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_39_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_95_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__36_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_44_ccff_tail[0]));

	grid_clb grid_clb_6__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_40_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_96_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__37_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_45_ccff_tail[0]));

	grid_clb grid_clb_6__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_41_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_97_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__38_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_46_ccff_tail[0]));

	grid_clb grid_clb_6__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__5_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__5_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__5_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__5_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__5_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__5_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__5_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__5_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__5_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__5_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__5_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__5_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__5_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__5_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__5_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__5_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_6__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_116_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__39_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_47_ccff_tail[0]));

	grid_clb grid_clb_7__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_42_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_98_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__40_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_48_ccff_tail[0]));

	grid_clb grid_clb_7__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_43_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_99_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__41_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_49_ccff_tail[0]));

	grid_clb grid_clb_7__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_44_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_100_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__42_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_50_ccff_tail[0]));

	grid_clb grid_clb_7__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_45_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_101_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__43_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_51_ccff_tail[0]));

	grid_clb grid_clb_7__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_46_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_102_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__44_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_52_ccff_tail[0]));

	grid_clb grid_clb_7__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_47_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_103_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__45_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_53_ccff_tail[0]));

	grid_clb grid_clb_7__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_48_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_104_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__46_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_54_ccff_tail[0]));

	grid_clb grid_clb_7__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__6_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__6_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__6_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__6_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__6_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__6_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__6_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__6_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__6_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__6_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__6_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__6_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__6_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__6_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__6_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__6_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_7__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_117_out[0]),
		.right_width_0_height_0__pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__47_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_55_ccff_tail[0]));

	grid_clb grid_clb_8__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_49_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_105_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__0_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__0_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__0_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__0_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__0_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__0_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__0_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__0_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__0_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__0_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__0_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__0_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__0_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__0_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__0_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__0_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__48_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_56_ccff_tail[0]));

	grid_clb grid_clb_8__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_50_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_106_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__1_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__1_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__1_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__1_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__1_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__1_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__1_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__1_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__1_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__1_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__1_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__1_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__1_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__1_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__1_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__1_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__49_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_57_ccff_tail[0]));

	grid_clb grid_clb_8__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_51_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_107_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__2_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__2_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__2_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__2_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__2_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__2_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__2_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__2_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__2_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__2_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__2_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__2_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__2_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__2_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__2_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__2_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__50_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_58_ccff_tail[0]));

	grid_clb grid_clb_8__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_52_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_108_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__3_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__3_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__3_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__3_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__3_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__3_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__3_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__3_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__3_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__3_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__3_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__3_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__3_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__3_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__3_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__3_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__51_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_59_ccff_tail[0]));

	grid_clb grid_clb_8__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_53_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_109_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__4_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__4_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__4_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__4_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__4_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__4_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__4_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__4_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__4_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__4_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__4_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__4_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__4_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__4_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__4_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__4_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__52_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_60_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_60_ccff_tail[0]));

	grid_clb grid_clb_8__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_54_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_110_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__5_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__5_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__5_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__5_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__5_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__5_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__5_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__5_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__5_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__5_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__5_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__5_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__5_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__5_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__5_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__5_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__53_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_61_ccff_tail[0]));

	grid_clb grid_clb_8__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(direct_interc_55_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_111_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__6_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__6_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__6_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__6_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__6_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__6_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__6_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__6_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__6_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__6_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__6_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__6_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__6_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__6_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__6_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__6_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__54_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_62_ccff_tail[0]));

	grid_clb grid_clb_8__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.top_width_0_height_0__pin_0_(cbx_1__8__7_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_1_(cbx_1__8__7_bottom_grid_pin_1_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__8__7_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_3_(cbx_1__8__7_bottom_grid_pin_3_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__8__7_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_5_(cbx_1__8__7_bottom_grid_pin_5_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__8__7_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_7_(cbx_1__8__7_bottom_grid_pin_7_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__8__7_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_9_(cbx_1__8__7_bottom_grid_pin_9_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__8__7_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_11_(cbx_1__8__7_bottom_grid_pin_11_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__8__7_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_13_(cbx_1__8__7_bottom_grid_pin_13_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__8__7_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_15_(cbx_1__8__7_bottom_grid_pin_15_[0]),
		.top_width_0_height_0__pin_32_(grid_clb_8__8__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(direct_interc_118_out[0]),
		.right_width_0_height_0__pin_16_(cby_8__1__7_left_grid_pin_16_[0]),
		.right_width_0_height_0__pin_17_(cby_8__1__7_left_grid_pin_17_[0]),
		.right_width_0_height_0__pin_18_(cby_8__1__7_left_grid_pin_18_[0]),
		.right_width_0_height_0__pin_19_(cby_8__1__7_left_grid_pin_19_[0]),
		.right_width_0_height_0__pin_20_(cby_8__1__7_left_grid_pin_20_[0]),
		.right_width_0_height_0__pin_21_(cby_8__1__7_left_grid_pin_21_[0]),
		.right_width_0_height_0__pin_22_(cby_8__1__7_left_grid_pin_22_[0]),
		.right_width_0_height_0__pin_23_(cby_8__1__7_left_grid_pin_23_[0]),
		.right_width_0_height_0__pin_24_(cby_8__1__7_left_grid_pin_24_[0]),
		.right_width_0_height_0__pin_25_(cby_8__1__7_left_grid_pin_25_[0]),
		.right_width_0_height_0__pin_26_(cby_8__1__7_left_grid_pin_26_[0]),
		.right_width_0_height_0__pin_27_(cby_8__1__7_left_grid_pin_27_[0]),
		.right_width_0_height_0__pin_28_(cby_8__1__7_left_grid_pin_28_[0]),
		.right_width_0_height_0__pin_29_(cby_8__1__7_left_grid_pin_29_[0]),
		.right_width_0_height_0__pin_30_(cby_8__1__7_left_grid_pin_30_[0]),
		.right_width_0_height_0__pin_31_(cby_8__1__7_left_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(clk[0]),
		.ccff_head(cby_1__1__55_ccff_tail[0]),
		.top_width_0_height_0__pin_34_upper(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
		.top_width_0_height_0__pin_34_lower(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
		.top_width_0_height_0__pin_35_upper(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
		.top_width_0_height_0__pin_35_lower(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
		.top_width_0_height_0__pin_36_upper(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
		.top_width_0_height_0__pin_36_lower(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
		.top_width_0_height_0__pin_37_upper(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
		.top_width_0_height_0__pin_37_lower(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
		.top_width_0_height_0__pin_38_upper(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
		.top_width_0_height_0__pin_38_lower(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
		.top_width_0_height_0__pin_39_upper(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
		.top_width_0_height_0__pin_39_lower(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
		.top_width_0_height_0__pin_40_upper(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
		.top_width_0_height_0__pin_40_lower(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
		.top_width_0_height_0__pin_41_upper(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
		.top_width_0_height_0__pin_41_lower(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
		.right_width_0_height_0__pin_42_upper(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
		.right_width_0_height_0__pin_42_lower(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
		.right_width_0_height_0__pin_43_upper(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
		.right_width_0_height_0__pin_43_lower(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
		.right_width_0_height_0__pin_44_upper(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
		.right_width_0_height_0__pin_44_lower(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
		.right_width_0_height_0__pin_45_upper(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
		.right_width_0_height_0__pin_45_lower(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
		.right_width_0_height_0__pin_46_upper(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
		.right_width_0_height_0__pin_46_lower(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
		.right_width_0_height_0__pin_47_upper(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
		.right_width_0_height_0__pin_47_lower(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
		.right_width_0_height_0__pin_48_upper(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
		.right_width_0_height_0__pin_48_lower(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
		.right_width_0_height_0__pin_49_upper(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
		.right_width_0_height_0__pin_49_lower(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_63_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_1__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__0_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__0_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_0_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_2__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__1_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__1_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_1_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_3__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__2_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__2_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_2_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_2_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_2_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_4__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__3_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__3_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_3_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_3_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_3_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_5__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__4_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__4_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_4_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_4_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_4_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_6__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__5_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__5_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_5_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_5_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_5_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_7__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__6_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__6_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_6_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_6_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_6_ccff_tail[0]));

	grid_io_top_top grid_io_top_top_8__9_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
		.bottom_width_0_height_0__pin_0_(cbx_1__8__7_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__8__7_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_top_7_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_top_7_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_top_7_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__8_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
		.left_width_0_height_0__pin_0_(cby_8__1__7_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__7_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_0_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_0_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_0_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__7_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
		.left_width_0_height_0__pin_0_(cby_8__1__6_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__6_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_1_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_1_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_1_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__6_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]),
		.left_width_0_height_0__pin_0_(cby_8__1__5_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__5_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_2_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_2_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_2_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__5_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]),
		.left_width_0_height_0__pin_0_(cby_8__1__4_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__4_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_3_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_3_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_3_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__4_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]),
		.left_width_0_height_0__pin_0_(cby_8__1__3_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__3_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_4_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_4_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_4_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__3_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]),
		.left_width_0_height_0__pin_0_(cby_8__1__2_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__2_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_5_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_5_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_5_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__2_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]),
		.left_width_0_height_0__pin_0_(cby_8__1__1_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__1_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_6_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_6_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_6_ccff_tail[0]));

	grid_io_right_right grid_io_right_right_9__1_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]),
		.left_width_0_height_0__pin_0_(cby_8__1__0_right_grid_pin_0_[0]),
		.ccff_head(cby_8__1__0_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_right_7_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_right_7_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_right_7_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_8__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16:24]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16:24]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16:24]),
		.top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__7_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_0_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_7__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25:33]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25:33]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25:33]),
		.top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__6_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_1_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_6__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34:42]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34:42]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34:42]),
		.top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__5_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_2_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_5__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43:51]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43:51]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43:51]),
		.top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__4_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_3_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_4__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52:60]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52:60]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52:60]),
		.top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__3_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_4_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_3__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61:69]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61:69]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61:69]),
		.top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__2_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_5_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_2__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70:78]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70:78]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70:78]),
		.top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__1_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_6_ccff_tail[0]));

	grid_io_bottom_bottom grid_io_bottom_bottom_1__0_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79:87]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79:87]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79:87]),
		.top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.top_width_0_height_0__pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
		.top_width_0_height_0__pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
		.top_width_0_height_0__pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
		.top_width_0_height_0__pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
		.top_width_0_height_0__pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
		.top_width_0_height_0__pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
		.top_width_0_height_0__pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
		.top_width_0_height_0__pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
		.ccff_head(cbx_1__0__0_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_lower[0]),
		.top_width_0_height_0__pin_3_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_upper[0]),
		.top_width_0_height_0__pin_3_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_lower[0]),
		.top_width_0_height_0__pin_5_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_upper[0]),
		.top_width_0_height_0__pin_5_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_lower[0]),
		.top_width_0_height_0__pin_7_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_upper[0]),
		.top_width_0_height_0__pin_7_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_lower[0]),
		.top_width_0_height_0__pin_9_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_upper[0]),
		.top_width_0_height_0__pin_9_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_lower[0]),
		.top_width_0_height_0__pin_11_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_upper[0]),
		.top_width_0_height_0__pin_11_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_lower[0]),
		.top_width_0_height_0__pin_13_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_upper[0]),
		.top_width_0_height_0__pin_13_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_lower[0]),
		.top_width_0_height_0__pin_15_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_upper[0]),
		.top_width_0_height_0__pin_15_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_lower[0]),
		.top_width_0_height_0__pin_17_upper(grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_upper[0]),
		.top_width_0_height_0__pin_17_lower(grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_lower[0]),
		.ccff_tail(grid_io_bottom_bottom_7_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__1_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]),
		.right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__0_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_0_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_0_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_0_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__2_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]),
		.right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_1_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_1_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_1_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__3_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]),
		.right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__2_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_2_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_2_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_2_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__4_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]),
		.right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__3_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_3_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_3_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_3_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__5_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]),
		.right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__4_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_4_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_4_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_4_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__6_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]),
		.right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__5_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_5_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_5_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_5_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__7_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]),
		.right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__6_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_6_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_6_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_6_ccff_tail[0]));

	grid_io_left_left grid_io_left_left_0__8_ (
		.IO_ISOL_N(IO_ISOL_N[0]),
		.prog_clk(prog_clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]),
		.right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__7_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_left_7_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_left_7_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_left_7_ccff_tail[0]));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_0_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_upper[0]),
		.ccff_head(grid_io_bottom_bottom_7_ccff_tail[0]),
		.chany_top_out(sb_0__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
		.ccff_tail(ccff_tail[0]));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_1_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_0_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__0_ccff_tail[0]),
		.chany_top_out(sb_0__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__0_ccff_tail[0]));

	sb_0__1_ sb_0__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_2_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_1_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__1_ccff_tail[0]),
		.chany_top_out(sb_0__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__1_ccff_tail[0]));

	sb_0__1_ sb_0__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_3_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_2_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__2_ccff_tail[0]),
		.chany_top_out(sb_0__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__2_ccff_tail[0]));

	sb_0__1_ sb_0__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_4_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_3_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__3_ccff_tail[0]),
		.chany_top_out(sb_0__1__3_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__3_ccff_tail[0]));

	sb_0__1_ sb_0__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_5_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_4_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__4_ccff_tail[0]),
		.chany_top_out(sb_0__1__4_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__4_ccff_tail[0]));

	sb_0__1_ sb_0__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_6_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_5_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__5_ccff_tail[0]),
		.chany_top_out(sb_0__1__5_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__5_ccff_tail[0]));

	sb_0__1_ sb_0__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_left_7_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_6_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__6_ccff_tail[0]),
		.chany_top_out(sb_0__1__6_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__6_ccff_tail[0]));

	sb_0__8_ sb_0__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__0_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_left_7_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(grid_io_top_top_0_ccff_tail[0]),
		.chanx_right_out(sb_0__8__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__8__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__8__0_ccff_tail[0]));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_7_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_6_ccff_tail[0]),
		.chany_top_out(sb_1__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__0_ccff_tail[0]));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_6_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_5_ccff_tail[0]),
		.chany_top_out(sb_1__0__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__1_ccff_tail[0]));

	sb_1__0_ sb_3__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_5_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_4_ccff_tail[0]),
		.chany_top_out(sb_1__0__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__2_ccff_tail[0]));

	sb_1__0_ sb_4__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_4_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_3_ccff_tail[0]),
		.chany_top_out(sb_1__0__3_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__3_ccff_tail[0]));

	sb_1__0_ sb_5__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_3_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_2_ccff_tail[0]),
		.chany_top_out(sb_1__0__4_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__4_ccff_tail[0]));

	sb_1__0_ sb_6__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_2_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_1_ccff_tail[0]),
		.chany_top_out(sb_1__0__5_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__5_ccff_tail[0]));

	sb_1__0_ sb_7__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
		.right_bottom_grid_pin_1_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_3_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_upper[0]),
		.right_bottom_grid_pin_5_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_upper[0]),
		.right_bottom_grid_pin_7_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_upper[0]),
		.right_bottom_grid_pin_9_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_upper[0]),
		.right_bottom_grid_pin_11_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_upper[0]),
		.right_bottom_grid_pin_13_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_upper[0]),
		.right_bottom_grid_pin_15_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_upper[0]),
		.right_bottom_grid_pin_17_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_upper[0]),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_1_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_bottom_bottom_0_ccff_tail[0]),
		.chany_top_out(sb_1__0__6_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__6_ccff_tail[0]));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__7_ccff_tail[0]),
		.chany_top_out(sb_1__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__0_ccff_tail[0]));

	sb_1__1_ sb_1__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__8_ccff_tail[0]),
		.chany_top_out(sb_1__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__1_ccff_tail[0]));

	sb_1__1_ sb_1__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__9_ccff_tail[0]),
		.chany_top_out(sb_1__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__2_ccff_tail[0]));

	sb_1__1_ sb_1__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__10_ccff_tail[0]),
		.chany_top_out(sb_1__1__3_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__3_ccff_tail[0]));

	sb_1__1_ sb_1__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__11_ccff_tail[0]),
		.chany_top_out(sb_1__1__4_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__4_ccff_tail[0]));

	sb_1__1_ sb_1__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__12_ccff_tail[0]),
		.chany_top_out(sb_1__1__5_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__5_ccff_tail[0]));

	sb_1__1_ sb_1__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__13_ccff_tail[0]),
		.chany_top_out(sb_1__1__6_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__6_ccff_tail[0]));

	sb_1__1_ sb_2__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__14_ccff_tail[0]),
		.chany_top_out(sb_1__1__7_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__7_ccff_tail[0]));

	sb_1__1_ sb_2__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__15_ccff_tail[0]),
		.chany_top_out(sb_1__1__8_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__8_ccff_tail[0]));

	sb_1__1_ sb_2__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__16_ccff_tail[0]),
		.chany_top_out(sb_1__1__9_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__9_ccff_tail[0]));

	sb_1__1_ sb_2__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__17_ccff_tail[0]),
		.chany_top_out(sb_1__1__10_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__10_ccff_tail[0]));

	sb_1__1_ sb_2__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__18_ccff_tail[0]),
		.chany_top_out(sb_1__1__11_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__11_ccff_tail[0]));

	sb_1__1_ sb_2__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__19_ccff_tail[0]),
		.chany_top_out(sb_1__1__12_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__12_ccff_tail[0]));

	sb_1__1_ sb_2__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__20_ccff_tail[0]),
		.chany_top_out(sb_1__1__13_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__13_ccff_tail[0]));

	sb_1__1_ sb_3__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__21_ccff_tail[0]),
		.chany_top_out(sb_1__1__14_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__14_ccff_tail[0]));

	sb_1__1_ sb_3__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__22_ccff_tail[0]),
		.chany_top_out(sb_1__1__15_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__15_ccff_tail[0]));

	sb_1__1_ sb_3__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__23_ccff_tail[0]),
		.chany_top_out(sb_1__1__16_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__16_ccff_tail[0]));

	sb_1__1_ sb_3__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__24_ccff_tail[0]),
		.chany_top_out(sb_1__1__17_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__17_ccff_tail[0]));

	sb_1__1_ sb_3__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__25_ccff_tail[0]),
		.chany_top_out(sb_1__1__18_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__18_ccff_tail[0]));

	sb_1__1_ sb_3__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__26_ccff_tail[0]),
		.chany_top_out(sb_1__1__19_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__19_ccff_tail[0]));

	sb_1__1_ sb_3__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__27_ccff_tail[0]),
		.chany_top_out(sb_1__1__20_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__20_ccff_tail[0]));

	sb_1__1_ sb_4__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__28_ccff_tail[0]),
		.chany_top_out(sb_1__1__21_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__21_ccff_tail[0]));

	sb_1__1_ sb_4__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__29_ccff_tail[0]),
		.chany_top_out(sb_1__1__22_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__22_ccff_tail[0]));

	sb_1__1_ sb_4__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__30_ccff_tail[0]),
		.chany_top_out(sb_1__1__23_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__23_ccff_tail[0]));

	sb_1__1_ sb_4__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__31_ccff_tail[0]),
		.chany_top_out(sb_1__1__24_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__24_ccff_tail[0]));

	sb_1__1_ sb_4__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__32_ccff_tail[0]),
		.chany_top_out(sb_1__1__25_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__25_ccff_tail[0]));

	sb_1__1_ sb_4__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__33_ccff_tail[0]),
		.chany_top_out(sb_1__1__26_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__26_ccff_tail[0]));

	sb_1__1_ sb_4__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__34_ccff_tail[0]),
		.chany_top_out(sb_1__1__27_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__27_ccff_tail[0]));

	sb_1__1_ sb_5__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__35_ccff_tail[0]),
		.chany_top_out(sb_1__1__28_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__28_ccff_tail[0]));

	sb_1__1_ sb_5__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__36_ccff_tail[0]),
		.chany_top_out(sb_1__1__29_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__29_ccff_tail[0]));

	sb_1__1_ sb_5__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__37_ccff_tail[0]),
		.chany_top_out(sb_1__1__30_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__30_ccff_tail[0]));

	sb_1__1_ sb_5__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__38_ccff_tail[0]),
		.chany_top_out(sb_1__1__31_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__31_ccff_tail[0]));

	sb_1__1_ sb_5__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__39_ccff_tail[0]),
		.chany_top_out(sb_1__1__32_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__32_ccff_tail[0]));

	sb_1__1_ sb_5__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__40_ccff_tail[0]),
		.chany_top_out(sb_1__1__33_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__33_ccff_tail[0]));

	sb_1__1_ sb_5__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__41_ccff_tail[0]),
		.chany_top_out(sb_1__1__34_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__34_ccff_tail[0]));

	sb_1__1_ sb_6__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__42_ccff_tail[0]),
		.chany_top_out(sb_1__1__35_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__35_ccff_tail[0]));

	sb_1__1_ sb_6__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__43_ccff_tail[0]),
		.chany_top_out(sb_1__1__36_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__36_ccff_tail[0]));

	sb_1__1_ sb_6__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__44_ccff_tail[0]),
		.chany_top_out(sb_1__1__37_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__37_ccff_tail[0]));

	sb_1__1_ sb_6__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__45_ccff_tail[0]),
		.chany_top_out(sb_1__1__38_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__38_ccff_tail[0]));

	sb_1__1_ sb_6__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__46_ccff_tail[0]),
		.chany_top_out(sb_1__1__39_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__39_ccff_tail[0]));

	sb_1__1_ sb_6__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__47_ccff_tail[0]),
		.chany_top_out(sb_1__1__40_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__40_ccff_tail[0]));

	sb_1__1_ sb_6__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__48_ccff_tail[0]),
		.chany_top_out(sb_1__1__41_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__41_ccff_tail[0]));

	sb_1__1_ sb_7__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__49_ccff_tail[0]),
		.chany_top_out(sb_1__1__42_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__42_ccff_tail[0]));

	sb_1__1_ sb_7__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__50_ccff_tail[0]),
		.chany_top_out(sb_1__1__43_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__43_ccff_tail[0]));

	sb_1__1_ sb_7__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__51_ccff_tail[0]),
		.chany_top_out(sb_1__1__44_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__44_ccff_tail[0]));

	sb_1__1_ sb_7__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__52_ccff_tail[0]),
		.chany_top_out(sb_1__1__45_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__45_ccff_tail[0]));

	sb_1__1_ sb_7__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__53_ccff_tail[0]),
		.chany_top_out(sb_1__1__46_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__46_ccff_tail[0]));

	sb_1__1_ sb_7__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__54_ccff_tail[0]),
		.chany_top_out(sb_1__1__47_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__47_ccff_tail[0]));

	sb_1__1_ sb_7__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
		.chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
		.right_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(cbx_1__1__55_ccff_tail[0]),
		.chany_top_out(sb_1__1__48_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__48_ccff_tail[0]));

	sb_1__8_ sb_1__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__1_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__0_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_1_ccff_tail[0]),
		.chanx_right_out(sb_1__8__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__0_ccff_tail[0]));

	sb_1__8_ sb_2__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__2_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_2_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__1_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_2_ccff_tail[0]),
		.chanx_right_out(sb_1__8__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__1_ccff_tail[0]));

	sb_1__8_ sb_3__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__3_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_3_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__2_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_2_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_3_ccff_tail[0]),
		.chanx_right_out(sb_1__8__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__2_ccff_tail[0]));

	sb_1__8_ sb_4__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__4_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_4_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__3_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_3_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_4_ccff_tail[0]),
		.chanx_right_out(sb_1__8__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__3_ccff_tail[0]));

	sb_1__8_ sb_5__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__5_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_5_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__4_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_4_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_5_ccff_tail[0]),
		.chanx_right_out(sb_1__8__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__4_ccff_tail[0]));

	sb_1__8_ sb_6__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__6_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_6_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__5_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_5_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_6_ccff_tail[0]),
		.chanx_right_out(sb_1__8__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__5_ccff_tail[0]));

	sb_1__8_ sb_7__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__8__7_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_top_7_bottom_width_0_height_0__pin_1_upper[0]),
		.right_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
		.right_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
		.right_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
		.right_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
		.right_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
		.right_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
		.right_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
		.right_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
		.bottom_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__6_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_6_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_top_top_7_ccff_tail[0]),
		.chanx_right_out(sb_1__8__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__8__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__8__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__8__6_ccff_tail[0]));

	sb_8__0_ sb_8__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__0_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_7_left_width_0_height_0__pin_1_lower[0]),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
		.left_bottom_grid_pin_1_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_3_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_3_lower[0]),
		.left_bottom_grid_pin_5_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_5_lower[0]),
		.left_bottom_grid_pin_7_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_7_lower[0]),
		.left_bottom_grid_pin_9_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_9_lower[0]),
		.left_bottom_grid_pin_11_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_11_lower[0]),
		.left_bottom_grid_pin_13_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_13_lower[0]),
		.left_bottom_grid_pin_15_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_15_lower[0]),
		.left_bottom_grid_pin_17_(grid_io_bottom_bottom_0_top_width_0_height_0__pin_17_lower[0]),
		.ccff_head(grid_io_right_right_7_ccff_tail[0]),
		.chany_top_out(sb_8__0__0_chany_top_out[0:19]),
		.chanx_left_out(sb_8__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_8__0__0_ccff_tail[0]));

	sb_8__1_ sb_8__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__1_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_6_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__0_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_7_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_6_ccff_tail[0]),
		.chany_top_out(sb_8__1__0_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__0_ccff_tail[0]));

	sb_8__1_ sb_8__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__2_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_5_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__1_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_6_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_5_ccff_tail[0]),
		.chany_top_out(sb_8__1__1_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__1_ccff_tail[0]));

	sb_8__1_ sb_8__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__3_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_4_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__2_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_5_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_4_ccff_tail[0]),
		.chany_top_out(sb_8__1__2_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__2_ccff_tail[0]));

	sb_8__1_ sb_8__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__4_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_3_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__3_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_4_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_3_ccff_tail[0]),
		.chany_top_out(sb_8__1__3_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__3_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__3_ccff_tail[0]));

	sb_8__1_ sb_8__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__5_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_2_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__4_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_3_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_2_ccff_tail[0]),
		.chany_top_out(sb_8__1__4_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__4_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__4_ccff_tail[0]));

	sb_8__1_ sb_8__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__6_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_1_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__5_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_2_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_1_ccff_tail[0]),
		.chany_top_out(sb_8__1__5_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__5_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__5_ccff_tail[0]));

	sb_8__1_ sb_8__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_8__1__7_chany_bottom_out[0:19]),
		.top_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
		.top_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
		.top_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
		.top_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
		.top_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
		.top_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
		.top_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
		.top_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_right_0_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_8__1__6_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_1_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
		.left_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(grid_io_right_right_0_ccff_tail[0]),
		.chany_top_out(sb_8__1__6_chany_top_out[0:19]),
		.chany_bottom_out(sb_8__1__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__1__6_chanx_left_out[0:19]),
		.ccff_tail(sb_8__1__6_ccff_tail[0]));

	sb_8__8_ sb_8__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(cby_8__1__7_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_right_0_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
		.bottom_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
		.bottom_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
		.bottom_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
		.bottom_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
		.bottom_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
		.bottom_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
		.bottom_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
		.chanx_left_in(cbx_1__8__7_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_top_7_bottom_width_0_height_0__pin_1_lower[0]),
		.left_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
		.left_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
		.left_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
		.left_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
		.left_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
		.left_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
		.left_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
		.left_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
		.ccff_head(ccff_head[0]),
		.chany_bottom_out(sb_8__8__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_8__8__0_chanx_left_out[0:19]),
		.ccff_tail(sb_8__8__0_ccff_tail[0]));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__0_ccff_tail[0]));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__1_ccff_tail[0]));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__2_ccff_tail[0]));

	cbx_1__0_ cbx_4__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__3_ccff_tail[0]));

	cbx_1__0_ cbx_5__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__4_ccff_tail[0]));

	cbx_1__0_ cbx_6__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__5_ccff_tail[0]));

	cbx_1__0_ cbx_7__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__6_ccff_tail[0]));

	cbx_1__0_ cbx_8__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_8__0__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
		.ccff_tail(cbx_1__0__7_ccff_tail[0]));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__0_ccff_tail[0]));

	cbx_1__1_ cbx_1__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__1_ccff_tail[0]));

	cbx_1__1_ cbx_1__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__2_ccff_tail[0]));

	cbx_1__1_ cbx_1__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__3_ccff_tail[0]));

	cbx_1__1_ cbx_1__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__4_ccff_tail[0]));

	cbx_1__1_ cbx_1__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__5_ccff_tail[0]));

	cbx_1__1_ cbx_1__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__6_ccff_tail[0]));

	cbx_1__1_ cbx_2__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__7_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__7_ccff_tail[0]));

	cbx_1__1_ cbx_2__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__8_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__8_ccff_tail[0]));

	cbx_1__1_ cbx_2__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__9_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__9_ccff_tail[0]));

	cbx_1__1_ cbx_2__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__10_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__10_ccff_tail[0]));

	cbx_1__1_ cbx_2__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__11_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__11_ccff_tail[0]));

	cbx_1__1_ cbx_2__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__12_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__12_ccff_tail[0]));

	cbx_1__1_ cbx_2__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__13_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__13_ccff_tail[0]));

	cbx_1__1_ cbx_3__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__14_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__14_ccff_tail[0]));

	cbx_1__1_ cbx_3__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__15_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__15_ccff_tail[0]));

	cbx_1__1_ cbx_3__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__16_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__16_ccff_tail[0]));

	cbx_1__1_ cbx_3__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__17_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__17_ccff_tail[0]));

	cbx_1__1_ cbx_3__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__18_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__18_ccff_tail[0]));

	cbx_1__1_ cbx_3__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__19_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__19_ccff_tail[0]));

	cbx_1__1_ cbx_3__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__20_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__20_ccff_tail[0]));

	cbx_1__1_ cbx_4__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__21_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__21_ccff_tail[0]));

	cbx_1__1_ cbx_4__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__22_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__22_ccff_tail[0]));

	cbx_1__1_ cbx_4__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__23_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__23_ccff_tail[0]));

	cbx_1__1_ cbx_4__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__24_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__24_ccff_tail[0]));

	cbx_1__1_ cbx_4__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__25_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__25_ccff_tail[0]));

	cbx_1__1_ cbx_4__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__26_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__26_ccff_tail[0]));

	cbx_1__1_ cbx_4__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__27_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__27_ccff_tail[0]));

	cbx_1__1_ cbx_5__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__28_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__28_ccff_tail[0]));

	cbx_1__1_ cbx_5__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__29_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__29_ccff_tail[0]));

	cbx_1__1_ cbx_5__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__30_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__30_ccff_tail[0]));

	cbx_1__1_ cbx_5__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__31_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__31_ccff_tail[0]));

	cbx_1__1_ cbx_5__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__32_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__32_ccff_tail[0]));

	cbx_1__1_ cbx_5__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__33_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__33_ccff_tail[0]));

	cbx_1__1_ cbx_5__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__34_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__34_ccff_tail[0]));

	cbx_1__1_ cbx_6__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__35_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__35_ccff_tail[0]));

	cbx_1__1_ cbx_6__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__36_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__36_ccff_tail[0]));

	cbx_1__1_ cbx_6__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__37_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__37_ccff_tail[0]));

	cbx_1__1_ cbx_6__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__38_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__38_ccff_tail[0]));

	cbx_1__1_ cbx_6__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__39_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__39_ccff_tail[0]));

	cbx_1__1_ cbx_6__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__40_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__40_ccff_tail[0]));

	cbx_1__1_ cbx_6__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__41_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__41_ccff_tail[0]));

	cbx_1__1_ cbx_7__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__42_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__42_ccff_tail[0]));

	cbx_1__1_ cbx_7__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__43_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__43_ccff_tail[0]));

	cbx_1__1_ cbx_7__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__44_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__44_ccff_tail[0]));

	cbx_1__1_ cbx_7__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__45_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__45_ccff_tail[0]));

	cbx_1__1_ cbx_7__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__46_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__46_ccff_tail[0]));

	cbx_1__1_ cbx_7__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__47_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__47_ccff_tail[0]));

	cbx_1__1_ cbx_7__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__48_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__48_ccff_tail[0]));

	cbx_1__1_ cbx_8__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__49_ccff_tail[0]));

	cbx_1__1_ cbx_8__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__50_ccff_tail[0]));

	cbx_1__1_ cbx_8__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__51_ccff_tail[0]));

	cbx_1__1_ cbx_8__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__3_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__52_ccff_tail[0]));

	cbx_1__1_ cbx_8__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__4_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__53_ccff_tail[0]));

	cbx_1__1_ cbx_8__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__5_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__54_ccff_tail[0]));

	cbx_1__1_ cbx_8__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__1__6_chanx_left_out[0:19]),
		.ccff_head(sb_8__1__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
		.bottom_grid_pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__1__55_ccff_tail[0]));

	cbx_1__8_ cbx_1__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__8__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__0_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__0_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__0_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__0_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__0_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__0_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__0_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__0_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__0_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__0_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__0_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__0_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__0_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__0_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__0_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__0_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__0_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__0_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__0_ccff_tail[0]));

	cbx_1__8_ cbx_2__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__1_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__1_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__1_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__1_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__1_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__1_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__1_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__1_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__1_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__1_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__1_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__1_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__1_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__1_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__1_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__1_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__1_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__1_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__1_ccff_tail[0]));

	cbx_1__8_ cbx_3__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__2_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__2_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__2_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__2_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__2_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__2_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__2_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__2_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__2_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__2_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__2_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__2_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__2_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__2_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__2_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__2_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__2_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__2_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__2_ccff_tail[0]));

	cbx_1__8_ cbx_4__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__3_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__3_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__3_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__3_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__3_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__3_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__3_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__3_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__3_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__3_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__3_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__3_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__3_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__3_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__3_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__3_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__3_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__3_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__3_ccff_tail[0]));

	cbx_1__8_ cbx_5__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__4_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__4_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__4_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__4_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__4_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__4_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__4_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__4_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__4_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__4_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__4_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__4_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__4_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__4_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__4_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__4_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__4_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__4_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__4_ccff_tail[0]));

	cbx_1__8_ cbx_6__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__5_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__5_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__5_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__5_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__5_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__5_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__5_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__5_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__5_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__5_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__5_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__5_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__5_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__5_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__5_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__5_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__5_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__5_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__5_ccff_tail[0]));

	cbx_1__8_ cbx_7__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__8__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__8__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__6_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__6_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__6_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__6_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__6_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__6_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__6_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__6_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__6_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__6_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__6_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__6_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__6_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__6_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__6_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__6_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__6_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__6_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__6_ccff_tail[0]));

	cbx_1__8_ cbx_8__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__8__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_8__8__0_chanx_left_out[0:19]),
		.ccff_head(sb_8__8__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__8__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__8__7_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__8__7_top_grid_pin_0_[0]),
		.bottom_grid_pin_0_(cbx_1__8__7_bottom_grid_pin_0_[0]),
		.bottom_grid_pin_1_(cbx_1__8__7_bottom_grid_pin_1_[0]),
		.bottom_grid_pin_2_(cbx_1__8__7_bottom_grid_pin_2_[0]),
		.bottom_grid_pin_3_(cbx_1__8__7_bottom_grid_pin_3_[0]),
		.bottom_grid_pin_4_(cbx_1__8__7_bottom_grid_pin_4_[0]),
		.bottom_grid_pin_5_(cbx_1__8__7_bottom_grid_pin_5_[0]),
		.bottom_grid_pin_6_(cbx_1__8__7_bottom_grid_pin_6_[0]),
		.bottom_grid_pin_7_(cbx_1__8__7_bottom_grid_pin_7_[0]),
		.bottom_grid_pin_8_(cbx_1__8__7_bottom_grid_pin_8_[0]),
		.bottom_grid_pin_9_(cbx_1__8__7_bottom_grid_pin_9_[0]),
		.bottom_grid_pin_10_(cbx_1__8__7_bottom_grid_pin_10_[0]),
		.bottom_grid_pin_11_(cbx_1__8__7_bottom_grid_pin_11_[0]),
		.bottom_grid_pin_12_(cbx_1__8__7_bottom_grid_pin_12_[0]),
		.bottom_grid_pin_13_(cbx_1__8__7_bottom_grid_pin_13_[0]),
		.bottom_grid_pin_14_(cbx_1__8__7_bottom_grid_pin_14_[0]),
		.bottom_grid_pin_15_(cbx_1__8__7_bottom_grid_pin_15_[0]),
		.ccff_tail(cbx_1__8__7_ccff_tail[0]));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__0_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__0_ccff_tail[0]));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__1_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__1_ccff_tail[0]));

	cby_0__1_ cby_0__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__2_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__2_ccff_tail[0]));

	cby_0__1_ cby_0__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__3_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__3_ccff_tail[0]));

	cby_0__1_ cby_0__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__4_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__4_ccff_tail[0]));

	cby_0__1_ cby_0__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__5_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__5_ccff_tail[0]));

	cby_0__1_ cby_0__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__6_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__6_ccff_tail[0]));

	cby_0__1_ cby_0__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_0__8__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__8__0_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:19]),
		.left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__7_ccff_tail[0]));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_0_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__0_ccff_tail[0]));

	cby_1__1_ cby_1__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_1_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__1_ccff_tail[0]));

	cby_1__1_ cby_1__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_2_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__2_ccff_tail[0]));

	cby_1__1_ cby_1__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_3_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__3_ccff_tail[0]));

	cby_1__1_ cby_1__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_4_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__4_ccff_tail[0]));

	cby_1__1_ cby_1__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_5_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__5_ccff_tail[0]));

	cby_1__1_ cby_1__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_6_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__6_ccff_tail[0]));

	cby_1__1_ cby_1__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_7_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__7_ccff_tail[0]));

	cby_1__1_ cby_2__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_8_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__8_ccff_tail[0]));

	cby_1__1_ cby_2__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_9_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__9_ccff_tail[0]));

	cby_1__1_ cby_2__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_10_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__10_ccff_tail[0]));

	cby_1__1_ cby_2__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_11_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__11_ccff_tail[0]));

	cby_1__1_ cby_2__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_12_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__12_ccff_tail[0]));

	cby_1__1_ cby_2__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_13_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__13_ccff_tail[0]));

	cby_1__1_ cby_2__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_14_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__14_ccff_tail[0]));

	cby_1__1_ cby_2__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_15_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__15_ccff_tail[0]));

	cby_1__1_ cby_3__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_16_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__16_ccff_tail[0]));

	cby_1__1_ cby_3__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_17_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__17_ccff_tail[0]));

	cby_1__1_ cby_3__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_18_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__18_ccff_tail[0]));

	cby_1__1_ cby_3__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_19_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__19_ccff_tail[0]));

	cby_1__1_ cby_3__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_20_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__20_ccff_tail[0]));

	cby_1__1_ cby_3__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_21_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__21_ccff_tail[0]));

	cby_1__1_ cby_3__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_22_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__22_ccff_tail[0]));

	cby_1__1_ cby_3__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_23_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__23_ccff_tail[0]));

	cby_1__1_ cby_4__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_24_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__24_ccff_tail[0]));

	cby_1__1_ cby_4__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_25_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__25_ccff_tail[0]));

	cby_1__1_ cby_4__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_26_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__26_ccff_tail[0]));

	cby_1__1_ cby_4__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_27_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__27_ccff_tail[0]));

	cby_1__1_ cby_4__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_28_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__28_ccff_tail[0]));

	cby_1__1_ cby_4__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_29_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__29_ccff_tail[0]));

	cby_1__1_ cby_4__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_30_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__30_ccff_tail[0]));

	cby_1__1_ cby_4__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_31_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__31_ccff_tail[0]));

	cby_1__1_ cby_5__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_32_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__32_ccff_tail[0]));

	cby_1__1_ cby_5__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_33_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__33_ccff_tail[0]));

	cby_1__1_ cby_5__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_34_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__34_ccff_tail[0]));

	cby_1__1_ cby_5__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_35_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__35_ccff_tail[0]));

	cby_1__1_ cby_5__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_36_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__36_ccff_tail[0]));

	cby_1__1_ cby_5__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_37_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__37_ccff_tail[0]));

	cby_1__1_ cby_5__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_38_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__38_ccff_tail[0]));

	cby_1__1_ cby_5__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_39_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__39_ccff_tail[0]));

	cby_1__1_ cby_6__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_40_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__40_ccff_tail[0]));

	cby_1__1_ cby_6__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_41_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__41_ccff_tail[0]));

	cby_1__1_ cby_6__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_42_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__42_ccff_tail[0]));

	cby_1__1_ cby_6__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_43_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__43_ccff_tail[0]));

	cby_1__1_ cby_6__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_44_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__44_ccff_tail[0]));

	cby_1__1_ cby_6__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_45_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__45_ccff_tail[0]));

	cby_1__1_ cby_6__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_46_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__46_ccff_tail[0]));

	cby_1__1_ cby_6__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_47_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__47_ccff_tail[0]));

	cby_1__1_ cby_7__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_48_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__48_ccff_tail[0]));

	cby_1__1_ cby_7__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_49_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__49_ccff_tail[0]));

	cby_1__1_ cby_7__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_50_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__50_ccff_tail[0]));

	cby_1__1_ cby_7__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_51_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__51_ccff_tail[0]));

	cby_1__1_ cby_7__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_52_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__52_ccff_tail[0]));

	cby_1__1_ cby_7__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_53_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__53_ccff_tail[0]));

	cby_1__1_ cby_7__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_54_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__54_ccff_tail[0]));

	cby_1__1_ cby_7__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
		.chany_top_in(sb_1__8__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_55_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:19]),
		.left_grid_pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
		.ccff_tail(cby_1__1__55_ccff_tail[0]));

	cby_8__1_ cby_8__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_56_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__0_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__0_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__0_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__0_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__0_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__0_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__0_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__0_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__0_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__0_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__0_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__0_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__0_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__0_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__0_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__0_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__0_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__0_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__0_ccff_tail[0]));

	cby_8__1_ cby_8__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_57_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__1_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__1_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__1_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__1_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__1_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__1_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__1_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__1_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__1_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__1_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__1_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__1_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__1_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__1_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__1_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__1_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__1_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__1_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__1_ccff_tail[0]));

	cby_8__1_ cby_8__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_58_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__2_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__2_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__2_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__2_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__2_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__2_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__2_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__2_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__2_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__2_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__2_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__2_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__2_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__2_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__2_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__2_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__2_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__2_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__2_ccff_tail[0]));

	cby_8__1_ cby_8__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_59_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__3_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__3_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__3_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__3_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__3_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__3_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__3_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__3_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__3_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__3_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__3_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__3_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__3_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__3_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__3_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__3_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__3_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__3_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__3_ccff_tail[0]));

	cby_8__1_ cby_8__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_60_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__4_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__4_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__4_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__4_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__4_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__4_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__4_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__4_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__4_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__4_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__4_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__4_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__4_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__4_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__4_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__4_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__4_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__4_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__4_ccff_tail[0]));

	cby_8__1_ cby_8__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_61_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__5_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__5_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__5_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__5_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__5_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__5_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__5_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__5_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__5_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__5_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__5_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__5_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__5_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__5_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__5_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__5_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__5_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__5_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__5_ccff_tail[0]));

	cby_8__1_ cby_8__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_8__1__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_62_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__6_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__6_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__6_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__6_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__6_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__6_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__6_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__6_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__6_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__6_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__6_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__6_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__6_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__6_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__6_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__6_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__6_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__6_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__6_ccff_tail[0]));

	cby_8__1_ cby_8__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_8__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_8__8__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_63_ccff_tail[0]),
		.chany_bottom_out(cby_8__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_8__1__7_chany_top_out[0:19]),
		.right_grid_pin_0_(cby_8__1__7_right_grid_pin_0_[0]),
		.left_grid_pin_16_(cby_8__1__7_left_grid_pin_16_[0]),
		.left_grid_pin_17_(cby_8__1__7_left_grid_pin_17_[0]),
		.left_grid_pin_18_(cby_8__1__7_left_grid_pin_18_[0]),
		.left_grid_pin_19_(cby_8__1__7_left_grid_pin_19_[0]),
		.left_grid_pin_20_(cby_8__1__7_left_grid_pin_20_[0]),
		.left_grid_pin_21_(cby_8__1__7_left_grid_pin_21_[0]),
		.left_grid_pin_22_(cby_8__1__7_left_grid_pin_22_[0]),
		.left_grid_pin_23_(cby_8__1__7_left_grid_pin_23_[0]),
		.left_grid_pin_24_(cby_8__1__7_left_grid_pin_24_[0]),
		.left_grid_pin_25_(cby_8__1__7_left_grid_pin_25_[0]),
		.left_grid_pin_26_(cby_8__1__7_left_grid_pin_26_[0]),
		.left_grid_pin_27_(cby_8__1__7_left_grid_pin_27_[0]),
		.left_grid_pin_28_(cby_8__1__7_left_grid_pin_28_[0]),
		.left_grid_pin_29_(cby_8__1__7_left_grid_pin_29_[0]),
		.left_grid_pin_30_(cby_8__1__7_left_grid_pin_30_[0]),
		.left_grid_pin_31_(cby_8__1__7_left_grid_pin_31_[0]),
		.ccff_tail(cby_8__1__7_ccff_tail[0]));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_0_out[0]));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_1_out[0]));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_2_out[0]));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_3_out[0]));

	direct_interc direct_interc_4_ (
		.in(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_4_out[0]));

	direct_interc direct_interc_5_ (
		.in(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_5_out[0]));

	direct_interc direct_interc_6_ (
		.in(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_6_out[0]));

	direct_interc direct_interc_7_ (
		.in(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_7_out[0]));

	direct_interc direct_interc_8_ (
		.in(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_8_out[0]));

	direct_interc direct_interc_9_ (
		.in(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_9_out[0]));

	direct_interc direct_interc_10_ (
		.in(grid_clb_12_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_10_out[0]));

	direct_interc direct_interc_11_ (
		.in(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_11_out[0]));

	direct_interc direct_interc_12_ (
		.in(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_12_out[0]));

	direct_interc direct_interc_13_ (
		.in(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_13_out[0]));

	direct_interc direct_interc_14_ (
		.in(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_14_out[0]));

	direct_interc direct_interc_15_ (
		.in(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_15_out[0]));

	direct_interc direct_interc_16_ (
		.in(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_16_out[0]));

	direct_interc direct_interc_17_ (
		.in(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_17_out[0]));

	direct_interc direct_interc_18_ (
		.in(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_18_out[0]));

	direct_interc direct_interc_19_ (
		.in(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_19_out[0]));

	direct_interc direct_interc_20_ (
		.in(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_20_out[0]));

	direct_interc direct_interc_21_ (
		.in(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_21_out[0]));

	direct_interc direct_interc_22_ (
		.in(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_22_out[0]));

	direct_interc direct_interc_23_ (
		.in(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_23_out[0]));

	direct_interc direct_interc_24_ (
		.in(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_24_out[0]));

	direct_interc direct_interc_25_ (
		.in(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_25_out[0]));

	direct_interc direct_interc_26_ (
		.in(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_26_out[0]));

	direct_interc direct_interc_27_ (
		.in(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_27_out[0]));

	direct_interc direct_interc_28_ (
		.in(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_28_out[0]));

	direct_interc direct_interc_29_ (
		.in(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_29_out[0]));

	direct_interc direct_interc_30_ (
		.in(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_30_out[0]));

	direct_interc direct_interc_31_ (
		.in(grid_clb_36_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_31_out[0]));

	direct_interc direct_interc_32_ (
		.in(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_32_out[0]));

	direct_interc direct_interc_33_ (
		.in(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_33_out[0]));

	direct_interc direct_interc_34_ (
		.in(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_34_out[0]));

	direct_interc direct_interc_35_ (
		.in(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_35_out[0]));

	direct_interc direct_interc_36_ (
		.in(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_36_out[0]));

	direct_interc direct_interc_37_ (
		.in(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_37_out[0]));

	direct_interc direct_interc_38_ (
		.in(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_38_out[0]));

	direct_interc direct_interc_39_ (
		.in(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_39_out[0]));

	direct_interc direct_interc_40_ (
		.in(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_40_out[0]));

	direct_interc direct_interc_41_ (
		.in(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_41_out[0]));

	direct_interc direct_interc_42_ (
		.in(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_42_out[0]));

	direct_interc direct_interc_43_ (
		.in(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_43_out[0]));

	direct_interc direct_interc_44_ (
		.in(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_44_out[0]));

	direct_interc direct_interc_45_ (
		.in(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_45_out[0]));

	direct_interc direct_interc_46_ (
		.in(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_46_out[0]));

	direct_interc direct_interc_47_ (
		.in(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_47_out[0]));

	direct_interc direct_interc_48_ (
		.in(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_48_out[0]));

	direct_interc direct_interc_49_ (
		.in(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_49_out[0]));

	direct_interc direct_interc_50_ (
		.in(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_50_out[0]));

	direct_interc direct_interc_51_ (
		.in(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_51_out[0]));

	direct_interc direct_interc_52_ (
		.in(grid_clb_60_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_52_out[0]));

	direct_interc direct_interc_53_ (
		.in(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_53_out[0]));

	direct_interc direct_interc_54_ (
		.in(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_54_out[0]));

	direct_interc direct_interc_55_ (
		.in(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_55_out[0]));

	direct_interc direct_interc_56_ (
		.in(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_56_out[0]));

	direct_interc direct_interc_57_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_57_out[0]));

	direct_interc direct_interc_58_ (
		.in(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_58_out[0]));

	direct_interc direct_interc_59_ (
		.in(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_59_out[0]));

	direct_interc direct_interc_60_ (
		.in(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_60_out[0]));

	direct_interc direct_interc_61_ (
		.in(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_61_out[0]));

	direct_interc direct_interc_62_ (
		.in(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_62_out[0]));

	direct_interc direct_interc_63_ (
		.in(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_63_out[0]));

	direct_interc direct_interc_64_ (
		.in(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_64_out[0]));

	direct_interc direct_interc_65_ (
		.in(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_65_out[0]));

	direct_interc direct_interc_66_ (
		.in(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_66_out[0]));

	direct_interc direct_interc_67_ (
		.in(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_67_out[0]));

	direct_interc direct_interc_68_ (
		.in(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_68_out[0]));

	direct_interc direct_interc_69_ (
		.in(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_69_out[0]));

	direct_interc direct_interc_70_ (
		.in(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_70_out[0]));

	direct_interc direct_interc_71_ (
		.in(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_71_out[0]));

	direct_interc direct_interc_72_ (
		.in(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_72_out[0]));

	direct_interc direct_interc_73_ (
		.in(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_73_out[0]));

	direct_interc direct_interc_74_ (
		.in(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_74_out[0]));

	direct_interc direct_interc_75_ (
		.in(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_75_out[0]));

	direct_interc direct_interc_76_ (
		.in(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_76_out[0]));

	direct_interc direct_interc_77_ (
		.in(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_77_out[0]));

	direct_interc direct_interc_78_ (
		.in(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_78_out[0]));

	direct_interc direct_interc_79_ (
		.in(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_79_out[0]));

	direct_interc direct_interc_80_ (
		.in(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_80_out[0]));

	direct_interc direct_interc_81_ (
		.in(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_81_out[0]));

	direct_interc direct_interc_82_ (
		.in(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_82_out[0]));

	direct_interc direct_interc_83_ (
		.in(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_83_out[0]));

	direct_interc direct_interc_84_ (
		.in(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_84_out[0]));

	direct_interc direct_interc_85_ (
		.in(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_85_out[0]));

	direct_interc direct_interc_86_ (
		.in(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_86_out[0]));

	direct_interc direct_interc_87_ (
		.in(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_87_out[0]));

	direct_interc direct_interc_88_ (
		.in(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_88_out[0]));

	direct_interc direct_interc_89_ (
		.in(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_89_out[0]));

	direct_interc direct_interc_90_ (
		.in(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_90_out[0]));

	direct_interc direct_interc_91_ (
		.in(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_91_out[0]));

	direct_interc direct_interc_92_ (
		.in(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_92_out[0]));

	direct_interc direct_interc_93_ (
		.in(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_93_out[0]));

	direct_interc direct_interc_94_ (
		.in(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_94_out[0]));

	direct_interc direct_interc_95_ (
		.in(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_95_out[0]));

	direct_interc direct_interc_96_ (
		.in(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_96_out[0]));

	direct_interc direct_interc_97_ (
		.in(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_97_out[0]));

	direct_interc direct_interc_98_ (
		.in(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_98_out[0]));

	direct_interc direct_interc_99_ (
		.in(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_99_out[0]));

	direct_interc direct_interc_100_ (
		.in(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_100_out[0]));

	direct_interc direct_interc_101_ (
		.in(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_101_out[0]));

	direct_interc direct_interc_102_ (
		.in(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_102_out[0]));

	direct_interc direct_interc_103_ (
		.in(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_103_out[0]));

	direct_interc direct_interc_104_ (
		.in(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_104_out[0]));

	direct_interc direct_interc_105_ (
		.in(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_105_out[0]));

	direct_interc direct_interc_106_ (
		.in(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_106_out[0]));

	direct_interc direct_interc_107_ (
		.in(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_107_out[0]));

	direct_interc direct_interc_108_ (
		.in(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_108_out[0]));

	direct_interc direct_interc_109_ (
		.in(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_109_out[0]));

	direct_interc direct_interc_110_ (
		.in(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_110_out[0]));

	direct_interc direct_interc_111_ (
		.in(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_111_out[0]));

	direct_interc direct_interc_112_ (
		.in(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_112_out[0]));

	direct_interc direct_interc_113_ (
		.in(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_113_out[0]));

	direct_interc direct_interc_114_ (
		.in(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_114_out[0]));

	direct_interc direct_interc_115_ (
		.in(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_115_out[0]));

	direct_interc direct_interc_116_ (
		.in(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_116_out[0]));

	direct_interc direct_interc_117_ (
		.in(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_117_out[0]));

	direct_interc direct_interc_118_ (
		.in(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_118_out[0]));

endmodule
// ----- END Verilog module for fpga_top -----



