VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 123.000 BY 123.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 119.000 85.470 123.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 119.000 88.690 123.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 39.480 123.000 40.080 ;
    END
  END Test_en_E_in
  PIN Test_en_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 36.760 123.000 37.360 ;
    END
  END Test_en_E_out
  PIN Test_en_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END Test_en_W_in
  PIN Test_en_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END Test_en_W_out
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 32.710 10.640 34.310 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.700 10.640 62.300 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.690 10.640 90.290 111.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.715 10.640 20.315 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.705 10.640 48.305 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.695 10.640 76.295 111.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.685 10.640 104.285 111.760 ;
    END
  END VPWR
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 34.040 123.000 34.640 ;
    END
  END ccff_tail
  PIN clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 119.000 91.910 123.000 ;
    END
  END clk_0_N_in
  PIN clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END clk_0_S_in
  PIN prog_clk_0_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 44.920 123.000 45.520 ;
    END
  END prog_clk_0_E_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 42.200 123.000 42.800 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 119.000 95.130 123.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END prog_clk_0_W_out
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 47.640 123.000 48.240 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 50.360 123.000 50.960 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 53.080 123.000 53.680 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 55.800 123.000 56.400 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 58.520 123.000 59.120 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 61.240 123.000 61.840 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 63.960 123.000 64.560 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 66.680 123.000 67.280 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 69.400 123.000 70.000 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 72.120 123.000 72.720 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 74.840 123.000 75.440 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 77.560 123.000 78.160 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 80.280 123.000 80.880 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 83.000 123.000 83.600 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 85.720 123.000 86.320 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 88.440 123.000 89.040 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 12.280 123.000 12.880 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 91.160 123.000 91.760 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 15.000 123.000 15.600 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 93.880 123.000 94.480 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 17.720 123.000 18.320 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 96.600 123.000 97.200 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 20.440 123.000 21.040 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 99.320 123.000 99.920 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 23.160 123.000 23.760 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 102.040 123.000 102.640 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 25.880 123.000 26.480 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 104.760 123.000 105.360 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 28.600 123.000 29.200 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 107.480 123.000 108.080 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 31.320 123.000 31.920 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 110.200 123.000 110.800 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 119.000 27.510 123.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 119.000 59.710 123.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 119.000 62.930 123.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 119.000 66.150 123.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 119.000 69.370 123.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 119.000 72.590 123.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 119.000 75.810 123.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 119.000 30.730 123.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 119.000 33.950 123.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 119.000 79.030 123.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 119.000 82.250 123.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 119.000 98.350 123.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 119.000 1.750 123.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 119.000 101.570 123.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 119.000 4.970 123.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 119.000 104.790 123.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 119.000 8.190 123.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 119.000 108.010 123.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 119.000 11.410 123.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 119.000 111.230 123.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 119.000 14.630 123.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 119.000 114.450 123.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 119.000 17.850 123.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 119.000 37.170 123.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 119.000 117.670 123.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 119.000 21.070 123.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 119.000 120.890 123.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 119.000 24.290 123.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 119.000 40.390 123.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 119.000 43.610 123.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 119.000 46.830 123.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 119.000 50.050 123.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 119.000 53.270 123.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 119.000 56.490 123.000 ;
    END
  END top_width_0_height_0__pin_9_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 117.300 111.605 ;
      LAYER met1 ;
        RECT 1.450 10.640 120.910 114.200 ;
      LAYER met2 ;
        RECT 2.030 118.720 4.410 119.410 ;
        RECT 5.250 118.720 7.630 119.410 ;
        RECT 8.470 118.720 10.850 119.410 ;
        RECT 11.690 118.720 14.070 119.410 ;
        RECT 14.910 118.720 17.290 119.410 ;
        RECT 18.130 118.720 20.510 119.410 ;
        RECT 21.350 118.720 23.730 119.410 ;
        RECT 24.570 118.720 26.950 119.410 ;
        RECT 27.790 118.720 30.170 119.410 ;
        RECT 31.010 118.720 33.390 119.410 ;
        RECT 34.230 118.720 36.610 119.410 ;
        RECT 37.450 118.720 39.830 119.410 ;
        RECT 40.670 118.720 43.050 119.410 ;
        RECT 43.890 118.720 46.270 119.410 ;
        RECT 47.110 118.720 49.490 119.410 ;
        RECT 50.330 118.720 52.710 119.410 ;
        RECT 53.550 118.720 55.930 119.410 ;
        RECT 56.770 118.720 59.150 119.410 ;
        RECT 59.990 118.720 62.370 119.410 ;
        RECT 63.210 118.720 65.590 119.410 ;
        RECT 66.430 118.720 68.810 119.410 ;
        RECT 69.650 118.720 72.030 119.410 ;
        RECT 72.870 118.720 75.250 119.410 ;
        RECT 76.090 118.720 78.470 119.410 ;
        RECT 79.310 118.720 81.690 119.410 ;
        RECT 82.530 118.720 84.910 119.410 ;
        RECT 85.750 118.720 88.130 119.410 ;
        RECT 88.970 118.720 91.350 119.410 ;
        RECT 92.190 118.720 94.570 119.410 ;
        RECT 95.410 118.720 97.790 119.410 ;
        RECT 98.630 118.720 101.010 119.410 ;
        RECT 101.850 118.720 104.230 119.410 ;
        RECT 105.070 118.720 107.450 119.410 ;
        RECT 108.290 118.720 110.670 119.410 ;
        RECT 111.510 118.720 113.890 119.410 ;
        RECT 114.730 118.720 117.110 119.410 ;
        RECT 117.950 118.720 120.330 119.410 ;
        RECT 1.480 4.280 120.880 118.720 ;
        RECT 1.480 4.000 10.390 4.280 ;
        RECT 11.230 4.000 30.630 4.280 ;
        RECT 31.470 4.000 50.870 4.280 ;
        RECT 51.710 4.000 71.110 4.280 ;
        RECT 71.950 4.000 91.350 4.280 ;
        RECT 92.190 4.000 111.590 4.280 ;
        RECT 112.430 4.000 120.880 4.280 ;
      LAYER met3 ;
        RECT 4.000 111.200 119.000 111.685 ;
        RECT 4.000 109.800 118.600 111.200 ;
        RECT 4.000 108.480 119.000 109.800 ;
        RECT 4.000 107.800 118.600 108.480 ;
        RECT 4.400 107.080 118.600 107.800 ;
        RECT 4.400 106.400 119.000 107.080 ;
        RECT 4.000 105.760 119.000 106.400 ;
        RECT 4.000 104.360 118.600 105.760 ;
        RECT 4.000 103.040 119.000 104.360 ;
        RECT 4.000 101.640 118.600 103.040 ;
        RECT 4.000 100.320 119.000 101.640 ;
        RECT 4.000 98.920 118.600 100.320 ;
        RECT 4.000 97.600 119.000 98.920 ;
        RECT 4.000 96.200 118.600 97.600 ;
        RECT 4.000 94.880 119.000 96.200 ;
        RECT 4.000 93.480 118.600 94.880 ;
        RECT 4.000 92.160 119.000 93.480 ;
        RECT 4.000 90.760 118.600 92.160 ;
        RECT 4.000 89.440 119.000 90.760 ;
        RECT 4.000 88.040 118.600 89.440 ;
        RECT 4.000 86.720 119.000 88.040 ;
        RECT 4.000 85.320 118.600 86.720 ;
        RECT 4.000 84.000 119.000 85.320 ;
        RECT 4.000 82.600 118.600 84.000 ;
        RECT 4.000 81.280 119.000 82.600 ;
        RECT 4.000 79.880 118.600 81.280 ;
        RECT 4.000 78.560 119.000 79.880 ;
        RECT 4.000 77.200 118.600 78.560 ;
        RECT 4.400 77.160 118.600 77.200 ;
        RECT 4.400 75.840 119.000 77.160 ;
        RECT 4.400 75.800 118.600 75.840 ;
        RECT 4.000 74.440 118.600 75.800 ;
        RECT 4.000 73.120 119.000 74.440 ;
        RECT 4.000 71.720 118.600 73.120 ;
        RECT 4.000 70.400 119.000 71.720 ;
        RECT 4.000 69.000 118.600 70.400 ;
        RECT 4.000 67.680 119.000 69.000 ;
        RECT 4.000 66.280 118.600 67.680 ;
        RECT 4.000 64.960 119.000 66.280 ;
        RECT 4.000 63.560 118.600 64.960 ;
        RECT 4.000 62.240 119.000 63.560 ;
        RECT 4.000 60.840 118.600 62.240 ;
        RECT 4.000 59.520 119.000 60.840 ;
        RECT 4.000 58.120 118.600 59.520 ;
        RECT 4.000 56.800 119.000 58.120 ;
        RECT 4.000 55.400 118.600 56.800 ;
        RECT 4.000 54.080 119.000 55.400 ;
        RECT 4.000 52.680 118.600 54.080 ;
        RECT 4.000 51.360 119.000 52.680 ;
        RECT 4.000 49.960 118.600 51.360 ;
        RECT 4.000 48.640 119.000 49.960 ;
        RECT 4.000 47.240 118.600 48.640 ;
        RECT 4.000 46.600 119.000 47.240 ;
        RECT 4.400 45.920 119.000 46.600 ;
        RECT 4.400 45.200 118.600 45.920 ;
        RECT 4.000 44.520 118.600 45.200 ;
        RECT 4.000 43.200 119.000 44.520 ;
        RECT 4.000 41.800 118.600 43.200 ;
        RECT 4.000 40.480 119.000 41.800 ;
        RECT 4.000 39.080 118.600 40.480 ;
        RECT 4.000 37.760 119.000 39.080 ;
        RECT 4.000 36.360 118.600 37.760 ;
        RECT 4.000 35.040 119.000 36.360 ;
        RECT 4.000 33.640 118.600 35.040 ;
        RECT 4.000 32.320 119.000 33.640 ;
        RECT 4.000 30.920 118.600 32.320 ;
        RECT 4.000 29.600 119.000 30.920 ;
        RECT 4.000 28.200 118.600 29.600 ;
        RECT 4.000 26.880 119.000 28.200 ;
        RECT 4.000 25.480 118.600 26.880 ;
        RECT 4.000 24.160 119.000 25.480 ;
        RECT 4.000 22.760 118.600 24.160 ;
        RECT 4.000 21.440 119.000 22.760 ;
        RECT 4.000 20.040 118.600 21.440 ;
        RECT 4.000 18.720 119.000 20.040 ;
        RECT 4.000 17.320 118.600 18.720 ;
        RECT 4.000 16.000 119.000 17.320 ;
        RECT 4.400 14.600 118.600 16.000 ;
        RECT 4.000 13.280 119.000 14.600 ;
        RECT 4.000 11.880 118.600 13.280 ;
        RECT 4.000 10.715 119.000 11.880 ;
      LAYER met4 ;
        RECT 69.295 21.935 74.295 110.665 ;
        RECT 76.695 21.935 88.290 110.665 ;
        RECT 90.690 21.935 102.285 110.665 ;
        RECT 104.685 21.935 108.265 110.665 ;
  END
END grid_clb
END LIBRARY

