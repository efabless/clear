magic
tech sky130A
magscale 1 2
timestamp 1679357744
<< obsli1 >>
rect 1104 2159 49864 24497
<< obsm1 >>
rect 934 2128 49864 25560
<< metal2 >>
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26200 4858 27000
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26200 7434 27000
rect 8022 26200 8078 27000
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26200 10010 27000
rect 10598 26200 10654 27000
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26200 13230 27000
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26200 16450 27000
rect 17038 26200 17094 27000
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26200 20314 27000
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26200 23534 27000
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26200 25466 27000
rect 26054 26200 26110 27000
rect 26698 26200 26754 27000
rect 27342 26200 27398 27000
rect 27986 26200 28042 27000
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 37002 26200 37058 27000
rect 37646 26200 37702 27000
rect 38290 26200 38346 27000
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 40866 26200 40922 27000
rect 41510 26200 41566 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 1398 0 1454 800
rect 4066 0 4122 800
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 17406 0 17462 800
rect 20074 0 20130 800
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< obsm2 >>
rect 938 26144 2170 26330
rect 2338 26144 2814 26330
rect 2982 26144 3458 26330
rect 3626 26144 4102 26330
rect 4270 26144 4746 26330
rect 4914 26144 5390 26330
rect 5558 26144 6034 26330
rect 6202 26144 6678 26330
rect 6846 26144 7322 26330
rect 7490 26144 7966 26330
rect 8134 26144 8610 26330
rect 8778 26144 9254 26330
rect 9422 26144 9898 26330
rect 10066 26144 10542 26330
rect 10710 26144 11186 26330
rect 11354 26144 11830 26330
rect 11998 26144 12474 26330
rect 12642 26144 13118 26330
rect 13286 26144 13762 26330
rect 13930 26144 14406 26330
rect 14574 26144 15050 26330
rect 15218 26144 15694 26330
rect 15862 26144 16338 26330
rect 16506 26144 16982 26330
rect 17150 26144 17626 26330
rect 17794 26144 18270 26330
rect 18438 26144 18914 26330
rect 19082 26144 19558 26330
rect 19726 26144 20202 26330
rect 20370 26144 20846 26330
rect 21014 26144 21490 26330
rect 21658 26144 22134 26330
rect 22302 26144 22778 26330
rect 22946 26144 23422 26330
rect 23590 26144 24066 26330
rect 24234 26144 24710 26330
rect 24878 26144 25354 26330
rect 25522 26144 25998 26330
rect 26166 26144 26642 26330
rect 26810 26144 27286 26330
rect 27454 26144 27930 26330
rect 28098 26144 28574 26330
rect 28742 26144 29218 26330
rect 29386 26144 29862 26330
rect 30030 26144 30506 26330
rect 30674 26144 31150 26330
rect 31318 26144 31794 26330
rect 31962 26144 32438 26330
rect 32606 26144 33082 26330
rect 33250 26144 33726 26330
rect 33894 26144 34370 26330
rect 34538 26144 35014 26330
rect 35182 26144 35658 26330
rect 35826 26144 36302 26330
rect 36470 26144 36946 26330
rect 37114 26144 37590 26330
rect 37758 26144 38234 26330
rect 38402 26144 38878 26330
rect 39046 26144 39522 26330
rect 39690 26144 40166 26330
rect 40334 26144 40810 26330
rect 40978 26144 41454 26330
rect 41622 26144 42098 26330
rect 42266 26144 42742 26330
rect 42910 26144 43386 26330
rect 43554 26144 44030 26330
rect 44198 26144 44674 26330
rect 44842 26144 45318 26330
rect 45486 26144 45962 26330
rect 46130 26144 46606 26330
rect 46774 26144 47250 26330
rect 47418 26144 47894 26330
rect 48062 26144 48538 26330
rect 48706 26144 49476 26330
rect 938 856 49476 26144
rect 938 734 1342 856
rect 1510 734 4010 856
rect 4178 734 6678 856
rect 6846 734 9346 856
rect 9514 734 12014 856
rect 12182 734 14682 856
rect 14850 734 17350 856
rect 17518 734 20018 856
rect 20186 734 22686 856
rect 22854 734 25354 856
rect 25522 734 28022 856
rect 28190 734 30690 856
rect 30858 734 33358 856
rect 33526 734 36026 856
rect 36194 734 38694 856
rect 38862 734 41362 856
rect 41530 734 44030 856
rect 44198 734 46698 856
rect 46866 734 49366 856
<< metal3 >>
rect 0 25576 800 25696
rect 0 25168 800 25288
rect 0 24760 800 24880
rect 50200 24760 51000 24880
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 50200 23808 51000 23928
rect 0 23536 800 23656
rect 0 23128 800 23248
rect 0 22720 800 22840
rect 50200 22856 51000 22976
rect 0 22312 800 22432
rect 0 21904 800 22024
rect 50200 21904 51000 22024
rect 0 21496 800 21616
rect 0 21088 800 21208
rect 50200 20952 51000 21072
rect 0 20680 800 20800
rect 0 20272 800 20392
rect 0 19864 800 19984
rect 0 19456 800 19576
rect 0 19048 800 19168
rect 0 18640 800 18760
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17416 800 17536
rect 0 17008 800 17128
rect 0 16600 800 16720
rect 0 16192 800 16312
rect 0 15784 800 15904
rect 0 15376 800 15496
rect 0 14968 800 15088
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 0 13744 800 13864
rect 0 13336 800 13456
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12112 800 12232
rect 0 11704 800 11824
rect 0 11296 800 11416
rect 0 10888 800 11008
rect 0 10480 800 10600
rect 0 10072 800 10192
rect 0 9664 800 9784
rect 0 9256 800 9376
rect 0 8848 800 8968
rect 0 8440 800 8560
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6808 800 6928
rect 0 6400 800 6520
rect 0 5992 800 6112
rect 0 5584 800 5704
rect 0 5176 800 5296
rect 0 4768 800 4888
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 0 3544 800 3664
rect 0 3136 800 3256
rect 0 2728 800 2848
rect 0 2320 800 2440
rect 0 1912 800 2032
rect 0 1504 800 1624
<< obsm3 >>
rect 880 25496 50200 25669
rect 800 25368 50200 25496
rect 880 25088 50200 25368
rect 800 24960 50200 25088
rect 880 24680 50120 24960
rect 800 24552 50200 24680
rect 880 24272 50200 24552
rect 800 24144 50200 24272
rect 880 24008 50200 24144
rect 880 23864 50120 24008
rect 800 23736 50120 23864
rect 880 23728 50120 23736
rect 880 23456 50200 23728
rect 800 23328 50200 23456
rect 880 23056 50200 23328
rect 880 23048 50120 23056
rect 800 22920 50120 23048
rect 880 22776 50120 22920
rect 880 22640 50200 22776
rect 800 22512 50200 22640
rect 880 22232 50200 22512
rect 800 22104 50200 22232
rect 880 21824 50120 22104
rect 800 21696 50200 21824
rect 880 21416 50200 21696
rect 800 21288 50200 21416
rect 880 21152 50200 21288
rect 880 21008 50120 21152
rect 800 20880 50120 21008
rect 880 20872 50120 20880
rect 880 20600 50200 20872
rect 800 20472 50200 20600
rect 880 20192 50200 20472
rect 800 20064 50200 20192
rect 880 19784 50200 20064
rect 800 19656 50200 19784
rect 880 19376 50200 19656
rect 800 19248 50200 19376
rect 880 18968 50200 19248
rect 800 18840 50200 18968
rect 880 18560 50200 18840
rect 800 18432 50200 18560
rect 880 18152 50200 18432
rect 800 18024 50200 18152
rect 880 17744 50200 18024
rect 800 17616 50200 17744
rect 880 17336 50200 17616
rect 800 17208 50200 17336
rect 880 16928 50200 17208
rect 800 16800 50200 16928
rect 880 16520 50200 16800
rect 800 16392 50200 16520
rect 880 16112 50200 16392
rect 800 15984 50200 16112
rect 880 15704 50200 15984
rect 800 15576 50200 15704
rect 880 15296 50200 15576
rect 800 15168 50200 15296
rect 880 14888 50200 15168
rect 800 14760 50200 14888
rect 880 14480 50200 14760
rect 800 14352 50200 14480
rect 880 14072 50200 14352
rect 800 13944 50200 14072
rect 880 13664 50200 13944
rect 800 13536 50200 13664
rect 880 13256 50200 13536
rect 800 13128 50200 13256
rect 880 12848 50200 13128
rect 800 12720 50200 12848
rect 880 12440 50200 12720
rect 800 12312 50200 12440
rect 880 12032 50200 12312
rect 800 11904 50200 12032
rect 880 11624 50200 11904
rect 800 11496 50200 11624
rect 880 11216 50200 11496
rect 800 11088 50200 11216
rect 880 10808 50200 11088
rect 800 10680 50200 10808
rect 880 10400 50200 10680
rect 800 10272 50200 10400
rect 880 9992 50200 10272
rect 800 9864 50200 9992
rect 880 9584 50200 9864
rect 800 9456 50200 9584
rect 880 9176 50200 9456
rect 800 9048 50200 9176
rect 880 8768 50200 9048
rect 800 8640 50200 8768
rect 880 8360 50200 8640
rect 800 8232 50200 8360
rect 880 7952 50200 8232
rect 800 7824 50200 7952
rect 880 7544 50200 7824
rect 800 7416 50200 7544
rect 880 7136 50200 7416
rect 800 7008 50200 7136
rect 880 6728 50200 7008
rect 800 6600 50200 6728
rect 880 6320 50200 6600
rect 800 6192 50200 6320
rect 880 5912 50200 6192
rect 800 5784 50200 5912
rect 880 5504 50200 5784
rect 800 5376 50200 5504
rect 880 5096 50200 5376
rect 800 4968 50200 5096
rect 880 4688 50200 4968
rect 800 4560 50200 4688
rect 880 4280 50200 4560
rect 800 4152 50200 4280
rect 880 3872 50200 4152
rect 800 3744 50200 3872
rect 880 3464 50200 3744
rect 800 3336 50200 3464
rect 880 3056 50200 3336
rect 800 2928 50200 3056
rect 880 2648 50200 2928
rect 800 2520 50200 2648
rect 880 2240 50200 2520
rect 800 2112 50200 2240
rect 880 1832 50200 2112
rect 800 1704 50200 1832
rect 880 1531 50200 1704
<< metal4 >>
rect 2944 2128 3264 24528
rect 7944 2128 8264 24528
rect 12944 2128 13264 24528
rect 17944 2128 18264 24528
rect 22944 2128 23264 24528
rect 27944 2128 28264 24528
rect 32944 2128 33264 24528
rect 37944 2128 38264 24528
rect 42944 2128 43264 24528
rect 47944 2128 48264 24528
<< obsm4 >>
rect 3555 8195 7864 24173
rect 8344 8195 12864 24173
rect 13344 8195 17864 24173
rect 18344 8195 22864 24173
rect 23344 8195 27725 24173
<< labels >>
rlabel metal4 s 7944 2128 8264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 24528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 24528 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 1398 0 1454 800 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 48594 26200 48650 27000 6 ccff_head_1
port 4 nsew signal input
rlabel metal3 s 50200 20952 51000 21072 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 2226 26200 2282 27000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 chanx_left_in[0]
port 7 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[10]
port 8 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[11]
port 9 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[12]
port 10 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[13]
port 11 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[14]
port 12 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[15]
port 13 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[16]
port 14 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 chanx_left_in[17]
port 15 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[18]
port 16 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[19]
port 17 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 chanx_left_in[1]
port 18 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[20]
port 19 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[21]
port 20 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[22]
port 21 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[23]
port 22 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[24]
port 23 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 chanx_left_in[25]
port 24 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[26]
port 25 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[27]
port 26 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[28]
port 27 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 chanx_left_in[29]
port 28 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 chanx_left_in[2]
port 29 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 chanx_left_in[3]
port 30 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 chanx_left_in[4]
port 31 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[5]
port 32 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[6]
port 33 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[7]
port 34 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[8]
port 35 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[9]
port 36 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 37 nsew signal output
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[10]
port 38 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[11]
port 39 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 chanx_left_out[12]
port 40 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 chanx_left_out[13]
port 41 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 chanx_left_out[14]
port 42 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 chanx_left_out[15]
port 43 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[16]
port 44 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[17]
port 45 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[18]
port 46 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 chanx_left_out[19]
port 47 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 48 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 chanx_left_out[20]
port 49 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 chanx_left_out[21]
port 50 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 chanx_left_out[22]
port 51 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 chanx_left_out[23]
port 52 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 chanx_left_out[24]
port 53 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 chanx_left_out[25]
port 54 nsew signal output
rlabel metal3 s 0 24352 800 24472 6 chanx_left_out[26]
port 55 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 chanx_left_out[27]
port 56 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 chanx_left_out[28]
port 57 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 chanx_left_out[29]
port 58 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 59 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 60 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 61 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[5]
port 62 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[6]
port 63 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 chanx_left_out[7]
port 64 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 65 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 66 nsew signal output
rlabel metal2 s 22190 26200 22246 27000 6 chany_top_in[0]
port 67 nsew signal input
rlabel metal2 s 28630 26200 28686 27000 6 chany_top_in[10]
port 68 nsew signal input
rlabel metal2 s 29274 26200 29330 27000 6 chany_top_in[11]
port 69 nsew signal input
rlabel metal2 s 29918 26200 29974 27000 6 chany_top_in[12]
port 70 nsew signal input
rlabel metal2 s 30562 26200 30618 27000 6 chany_top_in[13]
port 71 nsew signal input
rlabel metal2 s 31206 26200 31262 27000 6 chany_top_in[14]
port 72 nsew signal input
rlabel metal2 s 31850 26200 31906 27000 6 chany_top_in[15]
port 73 nsew signal input
rlabel metal2 s 32494 26200 32550 27000 6 chany_top_in[16]
port 74 nsew signal input
rlabel metal2 s 33138 26200 33194 27000 6 chany_top_in[17]
port 75 nsew signal input
rlabel metal2 s 33782 26200 33838 27000 6 chany_top_in[18]
port 76 nsew signal input
rlabel metal2 s 34426 26200 34482 27000 6 chany_top_in[19]
port 77 nsew signal input
rlabel metal2 s 22834 26200 22890 27000 6 chany_top_in[1]
port 78 nsew signal input
rlabel metal2 s 35070 26200 35126 27000 6 chany_top_in[20]
port 79 nsew signal input
rlabel metal2 s 35714 26200 35770 27000 6 chany_top_in[21]
port 80 nsew signal input
rlabel metal2 s 36358 26200 36414 27000 6 chany_top_in[22]
port 81 nsew signal input
rlabel metal2 s 37002 26200 37058 27000 6 chany_top_in[23]
port 82 nsew signal input
rlabel metal2 s 37646 26200 37702 27000 6 chany_top_in[24]
port 83 nsew signal input
rlabel metal2 s 38290 26200 38346 27000 6 chany_top_in[25]
port 84 nsew signal input
rlabel metal2 s 38934 26200 38990 27000 6 chany_top_in[26]
port 85 nsew signal input
rlabel metal2 s 39578 26200 39634 27000 6 chany_top_in[27]
port 86 nsew signal input
rlabel metal2 s 40222 26200 40278 27000 6 chany_top_in[28]
port 87 nsew signal input
rlabel metal2 s 40866 26200 40922 27000 6 chany_top_in[29]
port 88 nsew signal input
rlabel metal2 s 23478 26200 23534 27000 6 chany_top_in[2]
port 89 nsew signal input
rlabel metal2 s 24122 26200 24178 27000 6 chany_top_in[3]
port 90 nsew signal input
rlabel metal2 s 24766 26200 24822 27000 6 chany_top_in[4]
port 91 nsew signal input
rlabel metal2 s 25410 26200 25466 27000 6 chany_top_in[5]
port 92 nsew signal input
rlabel metal2 s 26054 26200 26110 27000 6 chany_top_in[6]
port 93 nsew signal input
rlabel metal2 s 26698 26200 26754 27000 6 chany_top_in[7]
port 94 nsew signal input
rlabel metal2 s 27342 26200 27398 27000 6 chany_top_in[8]
port 95 nsew signal input
rlabel metal2 s 27986 26200 28042 27000 6 chany_top_in[9]
port 96 nsew signal input
rlabel metal2 s 2870 26200 2926 27000 6 chany_top_out[0]
port 97 nsew signal output
rlabel metal2 s 9310 26200 9366 27000 6 chany_top_out[10]
port 98 nsew signal output
rlabel metal2 s 9954 26200 10010 27000 6 chany_top_out[11]
port 99 nsew signal output
rlabel metal2 s 10598 26200 10654 27000 6 chany_top_out[12]
port 100 nsew signal output
rlabel metal2 s 11242 26200 11298 27000 6 chany_top_out[13]
port 101 nsew signal output
rlabel metal2 s 11886 26200 11942 27000 6 chany_top_out[14]
port 102 nsew signal output
rlabel metal2 s 12530 26200 12586 27000 6 chany_top_out[15]
port 103 nsew signal output
rlabel metal2 s 13174 26200 13230 27000 6 chany_top_out[16]
port 104 nsew signal output
rlabel metal2 s 13818 26200 13874 27000 6 chany_top_out[17]
port 105 nsew signal output
rlabel metal2 s 14462 26200 14518 27000 6 chany_top_out[18]
port 106 nsew signal output
rlabel metal2 s 15106 26200 15162 27000 6 chany_top_out[19]
port 107 nsew signal output
rlabel metal2 s 3514 26200 3570 27000 6 chany_top_out[1]
port 108 nsew signal output
rlabel metal2 s 15750 26200 15806 27000 6 chany_top_out[20]
port 109 nsew signal output
rlabel metal2 s 16394 26200 16450 27000 6 chany_top_out[21]
port 110 nsew signal output
rlabel metal2 s 17038 26200 17094 27000 6 chany_top_out[22]
port 111 nsew signal output
rlabel metal2 s 17682 26200 17738 27000 6 chany_top_out[23]
port 112 nsew signal output
rlabel metal2 s 18326 26200 18382 27000 6 chany_top_out[24]
port 113 nsew signal output
rlabel metal2 s 18970 26200 19026 27000 6 chany_top_out[25]
port 114 nsew signal output
rlabel metal2 s 19614 26200 19670 27000 6 chany_top_out[26]
port 115 nsew signal output
rlabel metal2 s 20258 26200 20314 27000 6 chany_top_out[27]
port 116 nsew signal output
rlabel metal2 s 20902 26200 20958 27000 6 chany_top_out[28]
port 117 nsew signal output
rlabel metal2 s 21546 26200 21602 27000 6 chany_top_out[29]
port 118 nsew signal output
rlabel metal2 s 4158 26200 4214 27000 6 chany_top_out[2]
port 119 nsew signal output
rlabel metal2 s 4802 26200 4858 27000 6 chany_top_out[3]
port 120 nsew signal output
rlabel metal2 s 5446 26200 5502 27000 6 chany_top_out[4]
port 121 nsew signal output
rlabel metal2 s 6090 26200 6146 27000 6 chany_top_out[5]
port 122 nsew signal output
rlabel metal2 s 6734 26200 6790 27000 6 chany_top_out[6]
port 123 nsew signal output
rlabel metal2 s 7378 26200 7434 27000 6 chany_top_out[7]
port 124 nsew signal output
rlabel metal2 s 8022 26200 8078 27000 6 chany_top_out[8]
port 125 nsew signal output
rlabel metal2 s 8666 26200 8722 27000 6 chany_top_out[9]
port 126 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 gfpga_pad_io_soc_dir[0]
port 127 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 gfpga_pad_io_soc_dir[1]
port 128 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 gfpga_pad_io_soc_dir[2]
port 129 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 gfpga_pad_io_soc_dir[3]
port 130 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 gfpga_pad_io_soc_in[0]
port 131 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 gfpga_pad_io_soc_in[1]
port 132 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 gfpga_pad_io_soc_in[2]
port 133 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 gfpga_pad_io_soc_in[3]
port 134 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 gfpga_pad_io_soc_out[0]
port 135 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 gfpga_pad_io_soc_out[1]
port 136 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 gfpga_pad_io_soc_out[2]
port 137 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 gfpga_pad_io_soc_out[3]
port 138 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 isol_n
port 139 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 prog_clk
port 140 nsew signal input
rlabel metal2 s 41510 26200 41566 27000 6 prog_reset_top_in
port 141 nsew signal input
rlabel metal2 s 42154 26200 42210 27000 6 reset_top_in
port 142 nsew signal input
rlabel metal2 s 42798 26200 42854 27000 6 test_enable_top_in
port 143 nsew signal input
rlabel metal2 s 44730 26200 44786 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 144 nsew signal input
rlabel metal2 s 45374 26200 45430 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 145 nsew signal input
rlabel metal2 s 46018 26200 46074 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 146 nsew signal input
rlabel metal2 s 46662 26200 46718 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 147 nsew signal input
rlabel metal2 s 47306 26200 47362 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 148 nsew signal input
rlabel metal2 s 47950 26200 48006 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 149 nsew signal input
rlabel metal2 s 43442 26200 43498 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 150 nsew signal input
rlabel metal2 s 44086 26200 44142 27000 6 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 151 nsew signal input
rlabel metal3 s 50200 21904 51000 22024 6 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 152 nsew signal input
rlabel metal3 s 50200 22856 51000 22976 6 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 153 nsew signal input
rlabel metal3 s 50200 23808 51000 23928 6 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 154 nsew signal input
rlabel metal3 s 50200 24760 51000 24880 6 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 155 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 top_width_0_height_0_subtile_0__pin_inpad_0_
port 156 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 top_width_0_height_0_subtile_1__pin_inpad_0_
port 157 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 top_width_0_height_0_subtile_2__pin_inpad_0_
port 158 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 top_width_0_height_0_subtile_3__pin_inpad_0_
port 159 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 51000 27000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2049652
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/bottom_right_tile/runs/23_03_20_17_14/results/signoff/bottom_right_tile.magic.gds
string GDS_START 170702
<< end >>

