magic
tech sky130A
magscale 1 2
timestamp 1656942998
<< viali >>
rect 2697 17289 2731 17323
rect 3433 17289 3467 17323
rect 4353 17289 4387 17323
rect 6653 17289 6687 17323
rect 11621 17289 11655 17323
rect 1685 17221 1719 17255
rect 2421 17221 2455 17255
rect 4721 17221 4755 17255
rect 12173 17221 12207 17255
rect 1961 17153 1995 17187
rect 2237 17153 2271 17187
rect 2881 17153 2915 17187
rect 3249 17153 3283 17187
rect 4077 17153 4111 17187
rect 4169 17153 4203 17187
rect 4537 17153 4571 17187
rect 6837 17153 6871 17187
rect 11805 17153 11839 17187
rect 12449 17153 12483 17187
rect 12817 17153 12851 17187
rect 7389 17085 7423 17119
rect 7665 17085 7699 17119
rect 13737 17085 13771 17119
rect 3893 17017 3927 17051
rect 7113 17017 7147 17051
rect 13829 17017 13863 17051
rect 2053 16949 2087 16983
rect 3157 16949 3191 16983
rect 5273 16949 5307 16983
rect 6101 16949 6135 16983
rect 7205 16949 7239 16983
rect 9965 16949 9999 16983
rect 12633 16949 12667 16983
rect 14197 16949 14231 16983
rect 8033 16745 8067 16779
rect 9781 16745 9815 16779
rect 6745 16677 6779 16711
rect 7757 16677 7791 16711
rect 5641 16609 5675 16643
rect 5733 16609 5767 16643
rect 7113 16609 7147 16643
rect 8493 16609 8527 16643
rect 8677 16609 8711 16643
rect 9505 16609 9539 16643
rect 10241 16609 10275 16643
rect 10333 16609 10367 16643
rect 11069 16609 11103 16643
rect 11161 16609 11195 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 13277 16609 13311 16643
rect 13461 16609 13495 16643
rect 14565 16609 14599 16643
rect 14657 16609 14691 16643
rect 1593 16541 1627 16575
rect 1869 16541 1903 16575
rect 2421 16541 2455 16575
rect 2973 16541 3007 16575
rect 3249 16541 3283 16575
rect 3617 16541 3651 16575
rect 3985 16541 4019 16575
rect 4629 16541 4663 16575
rect 5089 16541 5123 16575
rect 6009 16541 6043 16575
rect 6561 16541 6595 16575
rect 6929 16541 6963 16575
rect 11713 16541 11747 16575
rect 12725 16541 12759 16575
rect 15117 16541 15151 16575
rect 15393 16541 15427 16575
rect 2145 16473 2179 16507
rect 2697 16473 2731 16507
rect 8401 16473 8435 16507
rect 10977 16473 11011 16507
rect 12173 16473 12207 16507
rect 13185 16473 13219 16507
rect 13645 16473 13679 16507
rect 3433 16405 3467 16439
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 4445 16405 4479 16439
rect 4905 16405 4939 16439
rect 5181 16405 5215 16439
rect 5549 16405 5583 16439
rect 6377 16405 6411 16439
rect 7297 16405 7331 16439
rect 7389 16405 7423 16439
rect 7849 16405 7883 16439
rect 8953 16405 8987 16439
rect 9321 16405 9355 16439
rect 9413 16405 9447 16439
rect 10149 16405 10183 16439
rect 10609 16405 10643 16439
rect 11529 16405 11563 16439
rect 11805 16405 11839 16439
rect 12817 16405 12851 16439
rect 14105 16405 14139 16439
rect 14473 16405 14507 16439
rect 15577 16405 15611 16439
rect 4261 16201 4295 16235
rect 5273 16201 5307 16235
rect 5733 16201 5767 16235
rect 6929 16201 6963 16235
rect 7849 16201 7883 16235
rect 9045 16201 9079 16235
rect 10057 16201 10091 16235
rect 11529 16201 11563 16235
rect 11989 16201 12023 16235
rect 13737 16201 13771 16235
rect 14933 16201 14967 16235
rect 3148 16133 3182 16167
rect 8309 16133 8343 16167
rect 12725 16133 12759 16167
rect 12817 16133 12851 16167
rect 2329 16065 2363 16099
rect 5089 16065 5123 16099
rect 5917 16065 5951 16099
rect 6193 16065 6227 16099
rect 6653 16065 6687 16099
rect 7113 16065 7147 16099
rect 8217 16065 8251 16099
rect 9229 16065 9263 16099
rect 9413 16065 9447 16099
rect 10241 16065 10275 16099
rect 11345 16065 11379 16099
rect 11897 16065 11931 16099
rect 13645 16065 13679 16099
rect 14289 16065 14323 16099
rect 14565 16065 14599 16099
rect 2421 15997 2455 16031
rect 2605 15997 2639 16031
rect 2881 15997 2915 16031
rect 8401 15997 8435 16031
rect 9781 15997 9815 16031
rect 12081 15997 12115 16031
rect 13001 15997 13035 16031
rect 13829 15997 13863 16031
rect 4721 15929 4755 15963
rect 6469 15929 6503 15963
rect 7481 15929 7515 15963
rect 11161 15929 11195 15963
rect 13277 15929 13311 15963
rect 14749 15929 14783 15963
rect 1961 15861 1995 15895
rect 4353 15861 4387 15895
rect 4997 15861 5031 15895
rect 5549 15861 5583 15895
rect 7205 15861 7239 15895
rect 7757 15861 7791 15895
rect 8677 15861 8711 15895
rect 10333 15861 10367 15895
rect 12357 15861 12391 15895
rect 2881 15657 2915 15691
rect 12265 15657 12299 15691
rect 12449 15657 12483 15691
rect 12725 15657 12759 15691
rect 13645 15657 13679 15691
rect 11529 15589 11563 15623
rect 3157 15521 3191 15555
rect 11897 15521 11931 15555
rect 13277 15521 13311 15555
rect 13737 15521 13771 15555
rect 2421 15453 2455 15487
rect 4261 15453 4295 15487
rect 5733 15453 5767 15487
rect 7297 15453 7331 15487
rect 8769 15453 8803 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 13093 15453 13127 15487
rect 2145 15385 2179 15419
rect 3065 15385 3099 15419
rect 4506 15385 4540 15419
rect 7030 15385 7064 15419
rect 8502 15385 8536 15419
rect 9566 15385 9600 15419
rect 13185 15385 13219 15419
rect 2513 15317 2547 15351
rect 5641 15317 5675 15351
rect 5917 15317 5951 15351
rect 7389 15317 7423 15351
rect 10701 15317 10735 15351
rect 1685 15113 1719 15147
rect 4353 15113 4387 15147
rect 12909 15113 12943 15147
rect 14013 15113 14047 15147
rect 15669 15113 15703 15147
rect 2421 15045 2455 15079
rect 5948 15045 5982 15079
rect 8370 15045 8404 15079
rect 11805 15045 11839 15079
rect 11897 15045 11931 15079
rect 1777 14977 1811 15011
rect 2697 14977 2731 15011
rect 3994 14977 4028 15011
rect 4261 14977 4295 15011
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6828 14977 6862 15011
rect 8125 14977 8159 15011
rect 10710 14977 10744 15011
rect 10977 14977 11011 15011
rect 11069 14977 11103 15011
rect 13277 14977 13311 15011
rect 14473 14977 14507 15011
rect 1593 14909 1627 14943
rect 11713 14909 11747 14943
rect 13369 14909 13403 14943
rect 13553 14909 13587 14943
rect 12817 14841 12851 14875
rect 2145 14773 2179 14807
rect 2881 14773 2915 14807
rect 4813 14773 4847 14807
rect 7941 14773 7975 14807
rect 9505 14773 9539 14807
rect 9597 14773 9631 14807
rect 12265 14773 12299 14807
rect 14749 14773 14783 14807
rect 3893 14569 3927 14603
rect 7297 14569 7331 14603
rect 13093 14569 13127 14603
rect 14105 14569 14139 14603
rect 13001 14501 13035 14535
rect 11897 14433 11931 14467
rect 13645 14433 13679 14467
rect 14657 14433 14691 14467
rect 15485 14433 15519 14467
rect 2237 14365 2271 14399
rect 6581 14365 6615 14399
rect 6837 14365 6871 14399
rect 6929 14365 6963 14399
rect 8677 14365 8711 14399
rect 9321 14365 9355 14399
rect 9505 14365 9539 14399
rect 15393 14365 15427 14399
rect 2482 14297 2516 14331
rect 8410 14297 8444 14331
rect 9750 14297 9784 14331
rect 12173 14297 12207 14331
rect 13461 14297 13495 14331
rect 14473 14297 14507 14331
rect 3617 14229 3651 14263
rect 5457 14229 5491 14263
rect 7113 14229 7147 14263
rect 10885 14229 10919 14263
rect 12081 14229 12115 14263
rect 12541 14229 12575 14263
rect 13553 14229 13587 14263
rect 14565 14229 14599 14263
rect 14933 14229 14967 14263
rect 15301 14229 15335 14263
rect 4169 14025 4203 14059
rect 4721 14025 4755 14059
rect 9597 14025 9631 14059
rect 11897 14025 11931 14059
rect 12357 14025 12391 14059
rect 12817 14025 12851 14059
rect 13185 14025 13219 14059
rect 13645 14025 13679 14059
rect 14013 14025 14047 14059
rect 14473 14025 14507 14059
rect 14841 14025 14875 14059
rect 15301 14025 15335 14059
rect 3056 13957 3090 13991
rect 12725 13957 12759 13991
rect 15209 13957 15243 13991
rect 1961 13889 1995 13923
rect 2789 13889 2823 13923
rect 4261 13889 4295 13923
rect 4905 13889 4939 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 6929 13889 6963 13923
rect 7205 13889 7239 13923
rect 8033 13889 8067 13923
rect 8217 13889 8251 13923
rect 8484 13889 8518 13923
rect 13553 13889 13587 13923
rect 14381 13889 14415 13923
rect 1685 13821 1719 13855
rect 11253 13821 11287 13855
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 12909 13821 12943 13855
rect 13737 13821 13771 13855
rect 14565 13821 14599 13855
rect 15393 13821 15427 13855
rect 11529 13685 11563 13719
rect 7205 13481 7239 13515
rect 11897 13481 11931 13515
rect 13185 13481 13219 13515
rect 14289 13481 14323 13515
rect 14657 13481 14691 13515
rect 8769 13413 8803 13447
rect 11069 13413 11103 13447
rect 1777 13345 1811 13379
rect 4353 13345 4387 13379
rect 7389 13345 7423 13379
rect 11253 13345 11287 13379
rect 11437 13345 11471 13379
rect 13737 13345 13771 13379
rect 14105 13345 14139 13379
rect 15209 13345 15243 13379
rect 15485 13345 15519 13379
rect 1961 13277 1995 13311
rect 2513 13277 2547 13311
rect 4620 13277 4654 13311
rect 5825 13277 5859 13311
rect 7645 13277 7679 13311
rect 9137 13277 9171 13311
rect 10609 13277 10643 13311
rect 13093 13277 13127 13311
rect 13553 13277 13587 13311
rect 15117 13277 15151 13311
rect 1869 13209 1903 13243
rect 6092 13209 6126 13243
rect 10342 13209 10376 13243
rect 2329 13141 2363 13175
rect 2697 13141 2731 13175
rect 5733 13141 5767 13175
rect 9229 13141 9263 13175
rect 11529 13141 11563 13175
rect 12449 13141 12483 13175
rect 13645 13141 13679 13175
rect 14473 13141 14507 13175
rect 15025 13141 15059 13175
rect 3341 12937 3375 12971
rect 11897 12937 11931 12971
rect 12357 12937 12391 12971
rect 13369 12937 13403 12971
rect 14289 12937 14323 12971
rect 15485 12937 15519 12971
rect 1409 12801 1443 12835
rect 1961 12801 1995 12835
rect 2228 12801 2262 12835
rect 4546 12801 4580 12835
rect 4813 12801 4847 12835
rect 5089 12801 5123 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 6828 12801 6862 12835
rect 10618 12801 10652 12835
rect 11345 12801 11379 12835
rect 11805 12801 11839 12835
rect 13737 12801 13771 12835
rect 14657 12801 14691 12835
rect 15117 12801 15151 12835
rect 1593 12733 1627 12767
rect 5273 12733 5307 12767
rect 6009 12733 6043 12767
rect 10885 12733 10919 12767
rect 11621 12733 11655 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14749 12733 14783 12767
rect 14841 12733 14875 12767
rect 3433 12597 3467 12631
rect 7941 12597 7975 12631
rect 9321 12597 9355 12631
rect 9505 12597 9539 12631
rect 12265 12597 12299 12631
rect 1501 12393 1535 12427
rect 3525 12393 3559 12427
rect 7389 12393 7423 12427
rect 9413 12393 9447 12427
rect 12541 12393 12575 12427
rect 14381 12393 14415 12427
rect 14565 12393 14599 12427
rect 2145 12257 2179 12291
rect 5181 12257 5215 12291
rect 9229 12257 9263 12291
rect 10793 12257 10827 12291
rect 11897 12257 11931 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 15209 12257 15243 12291
rect 4914 12189 4948 12223
rect 6653 12189 6687 12223
rect 6745 12189 6779 12223
rect 7205 12189 7239 12223
rect 8769 12189 8803 12223
rect 1869 12121 1903 12155
rect 6386 12121 6420 12155
rect 8524 12121 8558 12155
rect 10526 12121 10560 12155
rect 12173 12121 12207 12155
rect 12725 12121 12759 12155
rect 13185 12121 13219 12155
rect 15025 12121 15059 12155
rect 1961 12053 1995 12087
rect 3801 12053 3835 12087
rect 5273 12053 5307 12087
rect 12081 12053 12115 12087
rect 12817 12053 12851 12087
rect 14289 12053 14323 12087
rect 14933 12053 14967 12087
rect 1593 11849 1627 11883
rect 2053 11849 2087 11883
rect 12265 11849 12299 11883
rect 5058 11781 5092 11815
rect 6469 11781 6503 11815
rect 6561 11781 6595 11815
rect 11069 11781 11103 11815
rect 11805 11781 11839 11815
rect 13553 11781 13587 11815
rect 1961 11713 1995 11747
rect 3341 11713 3375 11747
rect 3597 11713 3631 11747
rect 4813 11713 4847 11747
rect 7869 11713 7903 11747
rect 8125 11713 8159 11747
rect 11253 11713 11287 11747
rect 11897 11713 11931 11747
rect 13369 11713 13403 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 2237 11645 2271 11679
rect 11621 11645 11655 11679
rect 14197 11645 14231 11679
rect 2513 11509 2547 11543
rect 4721 11509 4755 11543
rect 6193 11509 6227 11543
rect 6745 11509 6779 11543
rect 13645 11509 13679 11543
rect 4445 11305 4479 11339
rect 6009 11305 6043 11339
rect 9505 11305 9539 11339
rect 11437 11305 11471 11339
rect 11805 11305 11839 11339
rect 13553 11305 13587 11339
rect 14657 11305 14691 11339
rect 14381 11237 14415 11271
rect 2329 11169 2363 11203
rect 5825 11169 5859 11203
rect 10885 11169 10919 11203
rect 12357 11169 12391 11203
rect 13277 11169 13311 11203
rect 15209 11169 15243 11203
rect 2053 11101 2087 11135
rect 2973 11101 3007 11135
rect 5558 11101 5592 11135
rect 10629 11101 10663 11135
rect 12173 11101 12207 11135
rect 13001 11101 13035 11135
rect 2697 11033 2731 11067
rect 9413 11033 9447 11067
rect 11713 11033 11747 11067
rect 12265 11033 12299 11067
rect 15025 11033 15059 11067
rect 1685 10965 1719 10999
rect 2145 10965 2179 10999
rect 12633 10965 12667 10999
rect 13093 10965 13127 10999
rect 13829 10965 13863 10999
rect 14565 10965 14599 10999
rect 15117 10965 15151 10999
rect 4077 10761 4111 10795
rect 4813 10761 4847 10795
rect 6377 10761 6411 10795
rect 12725 10761 12759 10795
rect 13093 10761 13127 10795
rect 13553 10761 13587 10795
rect 13921 10761 13955 10795
rect 14289 10761 14323 10795
rect 14381 10761 14415 10795
rect 8300 10693 8334 10727
rect 13461 10693 13495 10727
rect 15209 10693 15243 10727
rect 1501 10625 1535 10659
rect 3626 10625 3660 10659
rect 3893 10625 3927 10659
rect 6561 10625 6595 10659
rect 6828 10625 6862 10659
rect 8033 10625 8067 10659
rect 10618 10625 10652 10659
rect 10885 10625 10919 10659
rect 15117 10625 15151 10659
rect 1685 10557 1719 10591
rect 13645 10557 13679 10591
rect 14473 10557 14507 10591
rect 15301 10557 15335 10591
rect 9413 10489 9447 10523
rect 15577 10489 15611 10523
rect 2513 10421 2547 10455
rect 7941 10421 7975 10455
rect 9505 10421 9539 10455
rect 14749 10421 14783 10455
rect 3893 10217 3927 10251
rect 4353 10217 4387 10251
rect 7297 10217 7331 10251
rect 9505 10217 9539 10251
rect 11437 10217 11471 10251
rect 12265 10217 12299 10251
rect 13829 10217 13863 10251
rect 3617 10081 3651 10115
rect 5917 10081 5951 10115
rect 10885 10081 10919 10115
rect 11989 10081 12023 10115
rect 12817 10081 12851 10115
rect 13185 10081 13219 10115
rect 13369 10081 13403 10115
rect 14197 10081 14231 10115
rect 14473 10081 14507 10115
rect 15117 10081 15151 10115
rect 15025 10013 15059 10047
rect 3372 9945 3406 9979
rect 5825 9945 5859 9979
rect 6184 9945 6218 9979
rect 10618 9945 10652 9979
rect 12633 9945 12667 9979
rect 14933 9945 14967 9979
rect 2237 9877 2271 9911
rect 7849 9877 7883 9911
rect 9137 9877 9171 9911
rect 9321 9877 9355 9911
rect 11805 9877 11839 9911
rect 11897 9877 11931 9911
rect 12725 9877 12759 9911
rect 13461 9877 13495 9911
rect 14565 9877 14599 9911
rect 2881 9673 2915 9707
rect 9597 9673 9631 9707
rect 12725 9673 12759 9707
rect 13001 9673 13035 9707
rect 13185 9673 13219 9707
rect 2513 9605 2547 9639
rect 6009 9605 6043 9639
rect 10802 9605 10836 9639
rect 15117 9605 15151 9639
rect 1777 9537 1811 9571
rect 2237 9537 2271 9571
rect 4005 9537 4039 9571
rect 5569 9537 5603 9571
rect 6644 9537 6678 9571
rect 8033 9537 8067 9571
rect 8300 9537 8334 9571
rect 12357 9537 12391 9571
rect 13553 9537 13587 9571
rect 14013 9537 14047 9571
rect 1501 9469 1535 9503
rect 1685 9469 1719 9503
rect 4261 9469 4295 9503
rect 5825 9469 5859 9503
rect 6377 9469 6411 9503
rect 11069 9469 11103 9503
rect 12173 9469 12207 9503
rect 12265 9469 12299 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 15209 9469 15243 9503
rect 15301 9469 15335 9503
rect 2145 9401 2179 9435
rect 7757 9401 7791 9435
rect 9689 9401 9723 9435
rect 4445 9333 4479 9367
rect 6101 9333 6135 9367
rect 7941 9333 7975 9367
rect 9413 9333 9447 9367
rect 14289 9333 14323 9367
rect 14749 9333 14783 9367
rect 15577 9333 15611 9367
rect 8585 9129 8619 9163
rect 9413 9129 9447 9163
rect 13185 9129 13219 9163
rect 5365 9061 5399 9095
rect 7113 9061 7147 9095
rect 13369 9061 13403 9095
rect 13737 9061 13771 9095
rect 3985 8993 4019 9027
rect 5733 8993 5767 9027
rect 12173 8993 12207 9027
rect 12633 8993 12667 9027
rect 14841 8993 14875 9027
rect 15301 8993 15335 9027
rect 2237 8925 2271 8959
rect 7205 8925 7239 8959
rect 8677 8925 8711 8959
rect 9229 8925 9263 8959
rect 10793 8925 10827 8959
rect 12081 8925 12115 8959
rect 13461 8925 13495 8959
rect 14565 8925 14599 8959
rect 15117 8925 15151 8959
rect 2504 8857 2538 8891
rect 4230 8857 4264 8891
rect 5549 8857 5583 8891
rect 5978 8857 6012 8891
rect 7450 8857 7484 8891
rect 10526 8857 10560 8891
rect 11529 8857 11563 8891
rect 11989 8857 12023 8891
rect 12725 8857 12759 8891
rect 3617 8789 3651 8823
rect 3801 8789 3835 8823
rect 11621 8789 11655 8823
rect 12817 8789 12851 8823
rect 14197 8789 14231 8823
rect 14657 8789 14691 8823
rect 8861 8585 8895 8619
rect 10425 8585 10459 8619
rect 11529 8585 11563 8619
rect 12449 8585 12483 8619
rect 12817 8585 12851 8619
rect 14013 8585 14047 8619
rect 14565 8585 14599 8619
rect 14933 8585 14967 8619
rect 15209 8585 15243 8619
rect 6920 8517 6954 8551
rect 11897 8517 11931 8551
rect 13921 8517 13955 8551
rect 14473 8517 14507 8551
rect 2872 8449 2906 8483
rect 4261 8449 4295 8483
rect 6653 8449 6687 8483
rect 9045 8449 9079 8483
rect 9301 8449 9335 8483
rect 11989 8449 12023 8483
rect 2605 8381 2639 8415
rect 12081 8381 12115 8415
rect 14289 8381 14323 8415
rect 15025 8381 15059 8415
rect 4169 8313 4203 8347
rect 4445 8313 4479 8347
rect 5549 8313 5583 8347
rect 5733 8313 5767 8347
rect 5917 8313 5951 8347
rect 6101 8313 6135 8347
rect 6469 8313 6503 8347
rect 3985 8245 4019 8279
rect 8033 8245 8067 8279
rect 2145 8041 2179 8075
rect 5733 8041 5767 8075
rect 7205 8041 7239 8075
rect 9045 8041 9079 8075
rect 9505 8041 9539 8075
rect 9689 8041 9723 8075
rect 12357 8041 12391 8075
rect 12909 8041 12943 8075
rect 1593 7905 1627 7939
rect 2789 7905 2823 7939
rect 5825 7905 5859 7939
rect 11069 7905 11103 7939
rect 13461 7905 13495 7939
rect 15117 7905 15151 7939
rect 4353 7837 4387 7871
rect 6081 7837 6115 7871
rect 10813 7837 10847 7871
rect 1777 7769 1811 7803
rect 2697 7769 2731 7803
rect 3249 7769 3283 7803
rect 4620 7769 4654 7803
rect 13369 7769 13403 7803
rect 14933 7769 14967 7803
rect 15393 7769 15427 7803
rect 1685 7701 1719 7735
rect 2237 7701 2271 7735
rect 2605 7701 2639 7735
rect 3157 7701 3191 7735
rect 13277 7701 13311 7735
rect 14565 7701 14599 7735
rect 15025 7701 15059 7735
rect 12357 7497 12391 7531
rect 12817 7497 12851 7531
rect 13185 7497 13219 7531
rect 13553 7497 13587 7531
rect 14289 7497 14323 7531
rect 15485 7497 15519 7531
rect 1685 7429 1719 7463
rect 8024 7429 8058 7463
rect 11253 7429 11287 7463
rect 11897 7429 11931 7463
rect 12725 7429 12759 7463
rect 1961 7361 1995 7395
rect 2513 7361 2547 7395
rect 4465 7361 4499 7395
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 5080 7361 5114 7395
rect 9496 7361 9530 7395
rect 14657 7361 14691 7395
rect 2237 7293 2271 7327
rect 6377 7293 6411 7327
rect 6561 7293 6595 7327
rect 7573 7293 7607 7327
rect 7757 7293 7791 7327
rect 9229 7293 9263 7327
rect 11989 7293 12023 7327
rect 12081 7293 12115 7327
rect 12909 7293 12943 7327
rect 13645 7293 13679 7327
rect 13737 7293 13771 7327
rect 14749 7293 14783 7327
rect 14841 7293 14875 7327
rect 3341 7157 3375 7191
rect 6193 7157 6227 7191
rect 9137 7157 9171 7191
rect 10609 7157 10643 7191
rect 11529 7157 11563 7191
rect 15209 7157 15243 7191
rect 6101 6953 6135 6987
rect 6561 6953 6595 6987
rect 8125 6953 8159 6987
rect 8677 6953 8711 6987
rect 10333 6953 10367 6987
rect 14105 6953 14139 6987
rect 14933 6953 14967 6987
rect 2513 6817 2547 6851
rect 2697 6817 2731 6851
rect 6745 6817 6779 6851
rect 8953 6817 8987 6851
rect 11529 6817 11563 6851
rect 11621 6817 11655 6851
rect 12541 6817 12575 6851
rect 13277 6817 13311 6851
rect 13461 6817 13495 6851
rect 13921 6817 13955 6851
rect 14657 6817 14691 6851
rect 15485 6817 15519 6851
rect 2973 6749 3007 6783
rect 4629 6749 4663 6783
rect 4896 6749 4930 6783
rect 9220 6749 9254 6783
rect 11437 6749 11471 6783
rect 13185 6749 13219 6783
rect 14565 6749 14599 6783
rect 15393 6749 15427 6783
rect 2421 6681 2455 6715
rect 3157 6681 3191 6715
rect 4445 6681 4479 6715
rect 7012 6681 7046 6715
rect 13645 6681 13679 6715
rect 14473 6681 14507 6715
rect 2053 6613 2087 6647
rect 3249 6613 3283 6647
rect 6009 6613 6043 6647
rect 11069 6613 11103 6647
rect 11897 6613 11931 6647
rect 12265 6613 12299 6647
rect 12357 6613 12391 6647
rect 12817 6613 12851 6647
rect 15301 6613 15335 6647
rect 4813 6409 4847 6443
rect 5273 6409 5307 6443
rect 6377 6409 6411 6443
rect 7205 6409 7239 6443
rect 8125 6409 8159 6443
rect 8493 6409 8527 6443
rect 8953 6409 8987 6443
rect 12265 6409 12299 6443
rect 12725 6409 12759 6443
rect 14013 6409 14047 6443
rect 14289 6409 14323 6443
rect 15117 6409 15151 6443
rect 15577 6409 15611 6443
rect 1685 6341 1719 6375
rect 2513 6341 2547 6375
rect 1961 6273 1995 6307
rect 2973 6273 3007 6307
rect 3240 6273 3274 6307
rect 8033 6273 8067 6307
rect 8861 6273 8895 6307
rect 9413 6273 9447 6307
rect 11253 6273 11287 6307
rect 11897 6273 11931 6307
rect 14381 6273 14415 6307
rect 15209 6273 15243 6307
rect 2237 6205 2271 6239
rect 2421 6205 2455 6239
rect 4905 6205 4939 6239
rect 5089 6205 5123 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 8217 6205 8251 6239
rect 9045 6205 9079 6239
rect 11069 6205 11103 6239
rect 11621 6205 11655 6239
rect 11805 6205 11839 6239
rect 13461 6205 13495 6239
rect 15301 6205 15335 6239
rect 4353 6137 4387 6171
rect 14749 6137 14783 6171
rect 2881 6069 2915 6103
rect 4445 6069 4479 6103
rect 7573 6069 7607 6103
rect 7665 6069 7699 6103
rect 12909 6069 12943 6103
rect 14657 6069 14691 6103
rect 1501 5865 1535 5899
rect 2605 5865 2639 5899
rect 8125 5865 8159 5899
rect 8401 5865 8435 5899
rect 9689 5865 9723 5899
rect 12265 5865 12299 5899
rect 14105 5865 14139 5899
rect 14933 5865 14967 5899
rect 2421 5797 2455 5831
rect 12173 5797 12207 5831
rect 1961 5729 1995 5763
rect 2145 5729 2179 5763
rect 3249 5729 3283 5763
rect 4721 5729 4755 5763
rect 4905 5729 4939 5763
rect 6101 5729 6135 5763
rect 6837 5729 6871 5763
rect 7389 5729 7423 5763
rect 7573 5729 7607 5763
rect 10241 5729 10275 5763
rect 11069 5729 11103 5763
rect 11529 5729 11563 5763
rect 12909 5729 12943 5763
rect 13645 5729 13679 5763
rect 14657 5729 14691 5763
rect 15485 5729 15519 5763
rect 1869 5661 1903 5695
rect 3525 5661 3559 5695
rect 6745 5661 6779 5695
rect 11713 5661 11747 5695
rect 13553 5661 13587 5695
rect 15301 5661 15335 5695
rect 2973 5593 3007 5627
rect 3801 5593 3835 5627
rect 5825 5593 5859 5627
rect 6653 5593 6687 5627
rect 7665 5593 7699 5627
rect 10057 5593 10091 5627
rect 11805 5593 11839 5627
rect 12725 5593 12759 5627
rect 13461 5593 13495 5627
rect 3065 5525 3099 5559
rect 4261 5525 4295 5559
rect 4629 5525 4663 5559
rect 5457 5525 5491 5559
rect 5917 5525 5951 5559
rect 6285 5525 6319 5559
rect 7205 5525 7239 5559
rect 8033 5525 8067 5559
rect 10149 5525 10183 5559
rect 10517 5525 10551 5559
rect 10885 5525 10919 5559
rect 10977 5525 11011 5559
rect 12633 5525 12667 5559
rect 13093 5525 13127 5559
rect 14473 5525 14507 5559
rect 14565 5525 14599 5559
rect 15393 5525 15427 5559
rect 3801 5321 3835 5355
rect 4629 5321 4663 5355
rect 5549 5321 5583 5355
rect 6009 5321 6043 5355
rect 6837 5321 6871 5355
rect 7481 5321 7515 5355
rect 7941 5321 7975 5355
rect 8493 5321 8527 5355
rect 9689 5321 9723 5355
rect 10057 5321 10091 5355
rect 10425 5321 10459 5355
rect 10517 5321 10551 5355
rect 10885 5321 10919 5355
rect 11621 5321 11655 5355
rect 11897 5321 11931 5355
rect 12081 5321 12115 5355
rect 12725 5321 12759 5355
rect 13369 5321 13403 5355
rect 13921 5321 13955 5355
rect 14473 5321 14507 5355
rect 14657 5321 14691 5355
rect 15025 5321 15059 5355
rect 2697 5253 2731 5287
rect 3985 5253 4019 5287
rect 6745 5253 6779 5287
rect 8953 5253 8987 5287
rect 9597 5253 9631 5287
rect 14197 5253 14231 5287
rect 2973 5185 3007 5219
rect 3433 5185 3467 5219
rect 4537 5185 4571 5219
rect 5641 5185 5675 5219
rect 7849 5185 7883 5219
rect 8309 5185 8343 5219
rect 8861 5185 8895 5219
rect 10977 5185 11011 5219
rect 14381 5185 14415 5219
rect 3249 5117 3283 5151
rect 3341 5117 3375 5151
rect 4813 5117 4847 5151
rect 5365 5117 5399 5151
rect 6929 5117 6963 5151
rect 7297 5117 7331 5151
rect 8125 5117 8159 5151
rect 9045 5117 9079 5151
rect 9413 5117 9447 5151
rect 10241 5117 10275 5151
rect 13461 5117 13495 5151
rect 13553 5117 13587 5151
rect 15117 5117 15151 5151
rect 15209 5117 15243 5151
rect 15485 5117 15519 5151
rect 11253 5049 11287 5083
rect 13001 5049 13035 5083
rect 4169 4981 4203 5015
rect 6377 4981 6411 5015
rect 4169 4777 4203 4811
rect 5181 4777 5215 4811
rect 5457 4777 5491 4811
rect 6377 4777 6411 4811
rect 8493 4777 8527 4811
rect 9321 4777 9355 4811
rect 9873 4777 9907 4811
rect 10701 4777 10735 4811
rect 13645 4777 13679 4811
rect 3985 4709 4019 4743
rect 8677 4709 8711 4743
rect 10793 4709 10827 4743
rect 13461 4709 13495 4743
rect 3249 4641 3283 4675
rect 3341 4641 3375 4675
rect 4905 4641 4939 4675
rect 6101 4641 6135 4675
rect 7849 4641 7883 4675
rect 7941 4641 7975 4675
rect 8401 4641 8435 4675
rect 10057 4641 10091 4675
rect 11345 4641 11379 4675
rect 12173 4641 12207 4675
rect 13001 4641 13035 4675
rect 14657 4641 14691 4675
rect 15485 4641 15519 4675
rect 2145 4573 2179 4607
rect 4721 4573 4755 4607
rect 5825 4573 5859 4607
rect 7757 4573 7791 4607
rect 9137 4573 9171 4607
rect 10333 4573 10367 4607
rect 11161 4573 11195 4607
rect 12909 4573 12943 4607
rect 14565 4573 14599 4607
rect 15301 4573 15335 4607
rect 15393 4573 15427 4607
rect 1869 4505 1903 4539
rect 11989 4505 12023 4539
rect 12817 4505 12851 4539
rect 13921 4505 13955 4539
rect 14473 4505 14507 4539
rect 2789 4437 2823 4471
rect 3157 4437 3191 4471
rect 4353 4437 4387 4471
rect 4813 4437 4847 4471
rect 5917 4437 5951 4471
rect 6469 4437 6503 4471
rect 7389 4437 7423 4471
rect 10241 4437 10275 4471
rect 11253 4437 11287 4471
rect 11621 4437 11655 4471
rect 12081 4437 12115 4471
rect 12449 4437 12483 4471
rect 14105 4437 14139 4471
rect 14933 4437 14967 4471
rect 1961 4233 1995 4267
rect 2881 4233 2915 4267
rect 3249 4233 3283 4267
rect 4077 4233 4111 4267
rect 5273 4233 5307 4267
rect 6469 4233 6503 4267
rect 8033 4233 8067 4267
rect 8493 4233 8527 4267
rect 8953 4233 8987 4267
rect 9505 4233 9539 4267
rect 9873 4233 9907 4267
rect 10333 4233 10367 4267
rect 11805 4233 11839 4267
rect 13093 4233 13127 4267
rect 13461 4233 13495 4267
rect 15669 4233 15703 4267
rect 5641 4165 5675 4199
rect 8861 4165 8895 4199
rect 10609 4165 10643 4199
rect 12173 4165 12207 4199
rect 14565 4165 14599 4199
rect 15025 4165 15059 4199
rect 1593 4097 1627 4131
rect 1869 4097 1903 4131
rect 2329 4097 2363 4131
rect 2421 4097 2455 4131
rect 3985 4097 4019 4131
rect 8125 4097 8159 4131
rect 9321 4097 9355 4131
rect 9965 4097 9999 4131
rect 10977 4097 11011 4131
rect 11713 4097 11747 4131
rect 12265 4097 12299 4131
rect 12909 4097 12943 4131
rect 13553 4097 13587 4131
rect 15485 4097 15519 4131
rect 2605 4029 2639 4063
rect 3341 4029 3375 4063
rect 3525 4029 3559 4063
rect 3801 4029 3835 4063
rect 4721 4029 4755 4063
rect 5733 4029 5767 4063
rect 5825 4029 5859 4063
rect 8217 4029 8251 4063
rect 9137 4029 9171 4063
rect 10057 4029 10091 4063
rect 12357 4029 12391 4063
rect 13645 4029 13679 4063
rect 14657 4029 14691 4063
rect 14749 4029 14783 4063
rect 4445 3961 4479 3995
rect 7665 3961 7699 3995
rect 10793 3961 10827 3995
rect 14197 3961 14231 3995
rect 4537 3893 4571 3927
rect 4905 3893 4939 3927
rect 12633 3893 12667 3927
rect 13921 3893 13955 3927
rect 15301 3893 15335 3927
rect 2697 3689 2731 3723
rect 3985 3689 4019 3723
rect 4905 3689 4939 3723
rect 5273 3689 5307 3723
rect 8033 3689 8067 3723
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 10149 3689 10183 3723
rect 12357 3689 12391 3723
rect 12449 3689 12483 3723
rect 12725 3689 12759 3723
rect 12909 3689 12943 3723
rect 14105 3689 14139 3723
rect 15669 3689 15703 3723
rect 6193 3621 6227 3655
rect 7849 3621 7883 3655
rect 9965 3621 9999 3655
rect 13093 3621 13127 3655
rect 4353 3553 4387 3587
rect 5917 3553 5951 3587
rect 6745 3553 6779 3587
rect 7573 3553 7607 3587
rect 9505 3553 9539 3587
rect 10701 3553 10735 3587
rect 11713 3553 11747 3587
rect 13737 3553 13771 3587
rect 14565 3553 14599 3587
rect 15209 3553 15243 3587
rect 15301 3553 15335 3587
rect 2145 3485 2179 3519
rect 2513 3485 2547 3519
rect 5733 3485 5767 3519
rect 7389 3485 7423 3519
rect 7481 3485 7515 3519
rect 11529 3485 11563 3519
rect 13553 3485 13587 3519
rect 1869 3417 1903 3451
rect 3249 3417 3283 3451
rect 4445 3417 4479 3451
rect 8769 3417 8803 3451
rect 9321 3417 9355 3451
rect 9413 3417 9447 3451
rect 10517 3417 10551 3451
rect 10977 3417 11011 3451
rect 11897 3417 11931 3451
rect 13645 3417 13679 3451
rect 2329 3349 2363 3383
rect 2881 3349 2915 3383
rect 3525 3349 3559 3383
rect 4537 3349 4571 3383
rect 4997 3349 5031 3383
rect 5365 3349 5399 3383
rect 5825 3349 5859 3383
rect 6561 3349 6595 3383
rect 6653 3349 6687 3383
rect 7021 3349 7055 3383
rect 10609 3349 10643 3383
rect 11345 3349 11379 3383
rect 11989 3349 12023 3383
rect 13185 3349 13219 3383
rect 14381 3349 14415 3383
rect 14749 3349 14783 3383
rect 15117 3349 15151 3383
rect 2881 3145 2915 3179
rect 4261 3145 4295 3179
rect 5365 3145 5399 3179
rect 6009 3145 6043 3179
rect 6193 3145 6227 3179
rect 6377 3145 6411 3179
rect 6745 3145 6779 3179
rect 8033 3145 8067 3179
rect 8309 3145 8343 3179
rect 8677 3145 8711 3179
rect 9137 3145 9171 3179
rect 9597 3145 9631 3179
rect 10885 3145 10919 3179
rect 11253 3145 11287 3179
rect 11621 3145 11655 3179
rect 11989 3145 12023 3179
rect 12449 3145 12483 3179
rect 12817 3145 12851 3179
rect 13277 3145 13311 3179
rect 2329 3077 2363 3111
rect 4629 3077 4663 3111
rect 12357 3077 12391 3111
rect 13185 3077 13219 3111
rect 15025 3077 15059 3111
rect 2053 3009 2087 3043
rect 2605 3009 2639 3043
rect 3065 3009 3099 3043
rect 3433 3009 3467 3043
rect 3801 3009 3835 3043
rect 4169 3009 4203 3043
rect 5457 3009 5491 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7849 3009 7883 3043
rect 8217 3009 8251 3043
rect 9505 3009 9539 3043
rect 10241 3009 10275 3043
rect 10793 3009 10827 3043
rect 11805 3009 11839 3043
rect 13645 3009 13679 3043
rect 14197 3009 14231 3043
rect 14749 3009 14783 3043
rect 15577 3009 15611 3043
rect 1777 2941 1811 2975
rect 4721 2941 4755 2975
rect 4905 2941 4939 2975
rect 5181 2941 5215 2975
rect 7389 2941 7423 2975
rect 8769 2941 8803 2975
rect 8861 2941 8895 2975
rect 9781 2941 9815 2975
rect 10977 2941 11011 2975
rect 12633 2941 12667 2975
rect 13369 2941 13403 2975
rect 13921 2941 13955 2975
rect 14473 2941 14507 2975
rect 3617 2873 3651 2907
rect 3985 2873 4019 2907
rect 7665 2873 7699 2907
rect 10425 2873 10459 2907
rect 15393 2873 15427 2907
rect 3249 2805 3283 2839
rect 5825 2805 5859 2839
rect 10057 2805 10091 2839
rect 3985 2601 4019 2635
rect 4813 2601 4847 2635
rect 4997 2601 5031 2635
rect 10701 2601 10735 2635
rect 11529 2601 11563 2635
rect 12449 2601 12483 2635
rect 12909 2601 12943 2635
rect 13093 2601 13127 2635
rect 13737 2601 13771 2635
rect 14565 2601 14599 2635
rect 2697 2533 2731 2567
rect 3249 2533 3283 2567
rect 7665 2533 7699 2567
rect 8033 2533 8067 2567
rect 10241 2533 10275 2567
rect 2145 2465 2179 2499
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 5641 2465 5675 2499
rect 7205 2465 7239 2499
rect 8769 2465 8803 2499
rect 9597 2465 9631 2499
rect 11345 2465 11379 2499
rect 13369 2465 13403 2499
rect 1961 2397 1995 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 3433 2397 3467 2431
rect 4445 2397 4479 2431
rect 5457 2397 5491 2431
rect 9229 2397 9263 2431
rect 10149 2397 10183 2431
rect 10425 2397 10459 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 13921 2397 13955 2431
rect 14381 2397 14415 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 4353 2329 4387 2363
rect 8309 2329 8343 2363
rect 12725 2329 12759 2363
rect 14933 2329 14967 2363
rect 15485 2329 15519 2363
rect 2329 2261 2363 2295
rect 3617 2261 3651 2295
rect 5089 2261 5123 2295
rect 9045 2261 9079 2295
rect 9321 2261 9355 2295
rect 9965 2261 9999 2295
rect 11161 2261 11195 2295
rect 11805 2261 11839 2295
rect 12173 2261 12207 2295
rect 13461 2261 13495 2295
rect 14197 2261 14231 2295
<< metal1 >>
rect 658 17484 664 17536
rect 716 17524 722 17536
rect 12066 17524 12072 17536
rect 716 17496 12072 17524
rect 716 17484 722 17496
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 2498 17280 2504 17332
rect 2556 17320 2562 17332
rect 2685 17323 2743 17329
rect 2685 17320 2697 17323
rect 2556 17292 2697 17320
rect 2556 17280 2562 17292
rect 2685 17289 2697 17292
rect 2731 17289 2743 17323
rect 2685 17283 2743 17289
rect 3421 17323 3479 17329
rect 3421 17289 3433 17323
rect 3467 17320 3479 17323
rect 3602 17320 3608 17332
rect 3467 17292 3608 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 4338 17320 4344 17332
rect 4299 17292 4344 17320
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 7650 17320 7656 17332
rect 6687 17292 7656 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 8904 17292 11621 17320
rect 8904 17280 8910 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 16482 17320 16488 17332
rect 12032 17292 16488 17320
rect 12032 17280 12038 17292
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 1394 17212 1400 17264
rect 1452 17252 1458 17264
rect 1673 17255 1731 17261
rect 1673 17252 1685 17255
rect 1452 17224 1685 17252
rect 1452 17212 1458 17224
rect 1673 17221 1685 17224
rect 1719 17221 1731 17255
rect 1673 17215 1731 17221
rect 2409 17255 2467 17261
rect 2409 17221 2421 17255
rect 2455 17252 2467 17255
rect 2590 17252 2596 17264
rect 2455 17224 2596 17252
rect 2455 17221 2467 17224
rect 2409 17215 2467 17221
rect 2590 17212 2596 17224
rect 2648 17252 2654 17264
rect 4709 17255 4767 17261
rect 4709 17252 4721 17255
rect 2648 17224 2912 17252
rect 2648 17212 2654 17224
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17184 2007 17187
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1995 17156 2237 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 2225 17153 2237 17156
rect 2271 17184 2283 17187
rect 2774 17184 2780 17196
rect 2271 17156 2780 17184
rect 2271 17153 2283 17156
rect 2225 17147 2283 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 2884 17193 2912 17224
rect 4080 17224 4721 17252
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 3142 17144 3148 17196
rect 3200 17184 3206 17196
rect 3237 17187 3295 17193
rect 3237 17184 3249 17187
rect 3200 17156 3249 17184
rect 3200 17144 3206 17156
rect 3237 17153 3249 17156
rect 3283 17153 3295 17187
rect 3237 17147 3295 17153
rect 3326 17144 3332 17196
rect 3384 17184 3390 17196
rect 4080 17193 4108 17224
rect 4709 17221 4721 17224
rect 4755 17221 4767 17255
rect 4709 17215 4767 17221
rect 12066 17212 12072 17264
rect 12124 17252 12130 17264
rect 12161 17255 12219 17261
rect 12161 17252 12173 17255
rect 12124 17224 12173 17252
rect 12124 17212 12130 17224
rect 12161 17221 12173 17224
rect 12207 17221 12219 17255
rect 12161 17215 12219 17221
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3384 17156 4077 17184
rect 3384 17144 3390 17156
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4212 17156 4537 17184
rect 4212 17144 4218 17156
rect 4525 17153 4537 17156
rect 4571 17153 4583 17187
rect 4525 17147 4583 17153
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 11793 17187 11851 17193
rect 6871 17156 7696 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 2792 17116 2820 17144
rect 4246 17116 4252 17128
rect 2792 17088 4252 17116
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 6362 17076 6368 17128
rect 6420 17116 6426 17128
rect 7668 17125 7696 17156
rect 11793 17153 11805 17187
rect 11839 17184 11851 17187
rect 12437 17187 12495 17193
rect 11839 17156 12388 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6420 17088 7389 17116
rect 6420 17076 6426 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 7653 17119 7711 17125
rect 7653 17085 7665 17119
rect 7699 17116 7711 17119
rect 10042 17116 10048 17128
rect 7699 17088 10048 17116
rect 7699 17085 7711 17088
rect 7653 17079 7711 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 12360 17116 12388 17156
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 12483 17156 12817 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12805 17153 12817 17156
rect 12851 17184 12863 17187
rect 15562 17184 15568 17196
rect 12851 17156 15568 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 12618 17116 12624 17128
rect 12360 17088 12624 17116
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13725 17119 13783 17125
rect 13725 17116 13737 17119
rect 13412 17088 13737 17116
rect 13412 17076 13418 17088
rect 13725 17085 13737 17088
rect 13771 17116 13783 17119
rect 16114 17116 16120 17128
rect 13771 17088 16120 17116
rect 13771 17085 13783 17088
rect 13725 17079 13783 17085
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 2866 17008 2872 17060
rect 2924 17048 2930 17060
rect 3881 17051 3939 17057
rect 3881 17048 3893 17051
rect 2924 17020 3893 17048
rect 2924 17008 2930 17020
rect 3881 17017 3893 17020
rect 3927 17017 3939 17051
rect 3881 17011 3939 17017
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7101 17051 7159 17057
rect 7101 17048 7113 17051
rect 7064 17020 7113 17048
rect 7064 17008 7070 17020
rect 7101 17017 7113 17020
rect 7147 17048 7159 17051
rect 7926 17048 7932 17060
rect 7147 17020 7932 17048
rect 7147 17017 7159 17020
rect 7101 17011 7159 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 13630 17048 13636 17060
rect 11020 17020 13636 17048
rect 11020 17008 11026 17020
rect 13630 17008 13636 17020
rect 13688 17048 13694 17060
rect 13817 17051 13875 17057
rect 13817 17048 13829 17051
rect 13688 17020 13829 17048
rect 13688 17008 13694 17020
rect 13817 17017 13829 17020
rect 13863 17048 13875 17051
rect 14550 17048 14556 17060
rect 13863 17020 14556 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 2038 16980 2044 16992
rect 1999 16952 2044 16980
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 3142 16980 3148 16992
rect 3055 16952 3148 16980
rect 3142 16940 3148 16952
rect 3200 16980 3206 16992
rect 3786 16980 3792 16992
rect 3200 16952 3792 16980
rect 3200 16940 3206 16952
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 6086 16980 6092 16992
rect 6047 16952 6092 16980
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 7190 16980 7196 16992
rect 7151 16952 7196 16980
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9916 16952 9965 16980
rect 9916 16940 9922 16952
rect 9953 16949 9965 16952
rect 9999 16980 10011 16983
rect 10594 16980 10600 16992
rect 9999 16952 10600 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 12618 16980 12624 16992
rect 12579 16952 12624 16980
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 14185 16983 14243 16989
rect 14185 16949 14197 16983
rect 14231 16980 14243 16983
rect 14734 16980 14740 16992
rect 14231 16952 14740 16980
rect 14231 16949 14243 16952
rect 14185 16943 14243 16949
rect 14734 16940 14740 16952
rect 14792 16940 14798 16992
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 5644 16748 8033 16776
rect 5644 16649 5672 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 9398 16776 9404 16788
rect 8444 16748 9404 16776
rect 8444 16736 8450 16748
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 9640 16748 9781 16776
rect 9640 16736 9646 16748
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 13170 16776 13176 16788
rect 9769 16739 9827 16745
rect 10244 16748 13176 16776
rect 6730 16708 6736 16720
rect 6691 16680 6736 16708
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 7745 16711 7803 16717
rect 7116 16680 7696 16708
rect 5629 16643 5687 16649
rect 2056 16612 2728 16640
rect 2056 16584 2084 16612
rect 1578 16572 1584 16584
rect 1539 16544 1584 16572
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 2038 16572 2044 16584
rect 1903 16544 2044 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2590 16572 2596 16584
rect 2455 16544 2596 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2590 16532 2596 16544
rect 2648 16532 2654 16584
rect 2700 16572 2728 16612
rect 5629 16609 5641 16643
rect 5675 16609 5687 16643
rect 5629 16603 5687 16609
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 7006 16640 7012 16652
rect 5776 16612 5821 16640
rect 6932 16612 7012 16640
rect 5776 16600 5782 16612
rect 2961 16575 3019 16581
rect 2961 16572 2973 16575
rect 2700 16544 2973 16572
rect 2961 16541 2973 16544
rect 3007 16541 3019 16575
rect 2961 16535 3019 16541
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 3602 16572 3608 16584
rect 3283 16544 3608 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 2130 16504 2136 16516
rect 2091 16476 2136 16504
rect 2130 16464 2136 16476
rect 2188 16464 2194 16516
rect 2222 16464 2228 16516
rect 2280 16504 2286 16516
rect 2685 16507 2743 16513
rect 2685 16504 2697 16507
rect 2280 16476 2697 16504
rect 2280 16464 2286 16476
rect 2685 16473 2697 16476
rect 2731 16473 2743 16507
rect 2685 16467 2743 16473
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 3252 16504 3280 16535
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3804 16544 3985 16572
rect 2832 16476 3280 16504
rect 2832 16464 2838 16476
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3292 16408 3433 16436
rect 3292 16396 3298 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 3694 16396 3700 16448
rect 3752 16436 3758 16448
rect 3804 16445 3832 16544
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 4614 16572 4620 16584
rect 4575 16544 4620 16572
rect 3973 16535 4031 16541
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16572 5135 16575
rect 5258 16572 5264 16584
rect 5123 16544 5264 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5592 16544 6009 16572
rect 5592 16532 5598 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6932 16581 6960 16612
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7116 16649 7144 16680
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7668 16640 7696 16680
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 7791 16680 8524 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 8386 16640 8392 16652
rect 7668 16612 8392 16640
rect 7101 16603 7159 16609
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 8496 16649 8524 16680
rect 9048 16680 10180 16708
rect 9048 16652 9076 16680
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 8665 16643 8723 16649
rect 8665 16609 8677 16643
rect 8711 16640 8723 16643
rect 9030 16640 9036 16652
rect 8711 16612 9036 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9456 16612 9505 16640
rect 9456 16600 9462 16612
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6420 16544 6561 16572
rect 6420 16532 6426 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16541 6975 16575
rect 9582 16572 9588 16584
rect 6917 16535 6975 16541
rect 7033 16544 9588 16572
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 7033 16504 7061 16544
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10152 16572 10180 16680
rect 10244 16649 10272 16748
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 12710 16708 12716 16720
rect 11072 16680 12716 16708
rect 11072 16649 11100 16680
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13354 16708 13360 16720
rect 13280 16680 13360 16708
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 11057 16603 11115 16609
rect 11149 16643 11207 16649
rect 11149 16609 11161 16643
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 10336 16572 10364 16603
rect 10152 16544 10364 16572
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 11164 16572 11192 16603
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 12124 16612 12265 16640
rect 12124 16600 12130 16612
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12986 16640 12992 16652
rect 12391 16612 12992 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 13280 16649 13308 16680
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13464 16680 14688 16708
rect 13464 16652 13492 16680
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13265 16603 13323 16609
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 14550 16640 14556 16652
rect 14511 16612 14556 16640
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 14660 16649 14688 16680
rect 14645 16643 14703 16649
rect 14645 16609 14657 16643
rect 14691 16609 14703 16643
rect 14645 16603 14703 16609
rect 10836 16544 11192 16572
rect 11701 16575 11759 16581
rect 10836 16532 10842 16544
rect 11701 16541 11713 16575
rect 11747 16572 11759 16575
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 11747 16544 12725 16572
rect 11747 16541 11759 16544
rect 11701 16535 11759 16541
rect 12713 16541 12725 16544
rect 12759 16572 12771 16575
rect 12894 16572 12900 16584
rect 12759 16544 12900 16572
rect 12759 16541 12771 16544
rect 12713 16535 12771 16541
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 15102 16572 15108 16584
rect 15063 16544 15108 16572
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16572 15439 16575
rect 15427 16544 15608 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 4120 16476 4476 16504
rect 4120 16464 4126 16476
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3752 16408 3801 16436
rect 3752 16396 3758 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16436 4215 16439
rect 4338 16436 4344 16448
rect 4203 16408 4344 16436
rect 4203 16405 4215 16408
rect 4157 16399 4215 16405
rect 4338 16396 4344 16408
rect 4396 16396 4402 16448
rect 4448 16445 4476 16476
rect 5552 16476 7061 16504
rect 8389 16507 8447 16513
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16405 4491 16439
rect 4433 16399 4491 16405
rect 4893 16439 4951 16445
rect 4893 16405 4905 16439
rect 4939 16436 4951 16439
rect 5074 16436 5080 16448
rect 4939 16408 5080 16436
rect 4939 16405 4951 16408
rect 4893 16399 4951 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5166 16396 5172 16448
rect 5224 16436 5230 16448
rect 5552 16445 5580 16476
rect 8389 16473 8401 16507
rect 8435 16504 8447 16507
rect 8435 16476 8984 16504
rect 8435 16473 8447 16476
rect 8389 16467 8447 16473
rect 5537 16439 5595 16445
rect 5224 16408 5269 16436
rect 5224 16396 5230 16408
rect 5537 16405 5549 16439
rect 5583 16405 5595 16439
rect 5537 16399 5595 16405
rect 6365 16439 6423 16445
rect 6365 16405 6377 16439
rect 6411 16436 6423 16439
rect 6454 16436 6460 16448
rect 6411 16408 6460 16436
rect 6411 16405 6423 16408
rect 6365 16399 6423 16405
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 7282 16436 7288 16448
rect 7243 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 8956 16445 8984 16476
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 10965 16507 11023 16513
rect 9180 16476 10732 16504
rect 9180 16464 9186 16476
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 7432 16408 7849 16436
rect 7432 16396 7438 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8941 16439 8999 16445
rect 8941 16405 8953 16439
rect 8987 16405 8999 16439
rect 9306 16436 9312 16448
rect 9267 16408 9312 16436
rect 8941 16399 8999 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9858 16436 9864 16448
rect 9447 16408 9864 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 10134 16436 10140 16448
rect 10095 16408 10140 16436
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10594 16436 10600 16448
rect 10555 16408 10600 16436
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 10704 16436 10732 16476
rect 10965 16473 10977 16507
rect 11011 16504 11023 16507
rect 12161 16507 12219 16513
rect 11011 16476 11836 16504
rect 11011 16473 11023 16476
rect 10965 16467 11023 16473
rect 11808 16445 11836 16476
rect 12161 16473 12173 16507
rect 12207 16504 12219 16507
rect 13173 16507 13231 16513
rect 12207 16476 12848 16504
rect 12207 16473 12219 16476
rect 12161 16467 12219 16473
rect 12820 16445 12848 16476
rect 13173 16473 13185 16507
rect 13219 16504 13231 16507
rect 13633 16507 13691 16513
rect 13633 16504 13645 16507
rect 13219 16476 13645 16504
rect 13219 16473 13231 16476
rect 13173 16467 13231 16473
rect 13633 16473 13645 16476
rect 13679 16473 13691 16507
rect 13633 16467 13691 16473
rect 11517 16439 11575 16445
rect 11517 16436 11529 16439
rect 10704 16408 11529 16436
rect 11517 16405 11529 16408
rect 11563 16405 11575 16439
rect 11517 16399 11575 16405
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16405 11851 16439
rect 11793 16399 11851 16405
rect 12805 16439 12863 16445
rect 12805 16405 12817 16439
rect 12851 16405 12863 16439
rect 12805 16399 12863 16405
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 14093 16439 14151 16445
rect 14093 16436 14105 16439
rect 13412 16408 14105 16436
rect 13412 16396 13418 16408
rect 14093 16405 14105 16408
rect 14139 16405 14151 16439
rect 14093 16399 14151 16405
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 14734 16436 14740 16448
rect 14507 16408 14740 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 15580 16445 15608 16544
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 15838 16436 15844 16448
rect 15611 16408 15844 16436
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 4249 16235 4307 16241
rect 4249 16201 4261 16235
rect 4295 16232 4307 16235
rect 4522 16232 4528 16244
rect 4295 16204 4528 16232
rect 4295 16201 4307 16204
rect 4249 16195 4307 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5442 16232 5448 16244
rect 5307 16204 5448 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 6178 16232 6184 16244
rect 5767 16204 6184 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7340 16204 7849 16232
rect 7340 16192 7346 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 8018 16192 8024 16244
rect 8076 16232 8082 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8076 16204 9045 16232
rect 8076 16192 8082 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 9033 16195 9091 16201
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9950 16232 9956 16244
rect 9732 16204 9956 16232
rect 9732 16192 9738 16204
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16201 10103 16235
rect 10045 16195 10103 16201
rect 3142 16173 3148 16176
rect 3136 16127 3148 16173
rect 3200 16164 3206 16176
rect 3200 16136 3236 16164
rect 3142 16124 3148 16127
rect 3200 16124 3206 16136
rect 3602 16124 3608 16176
rect 3660 16164 3666 16176
rect 7374 16164 7380 16176
rect 3660 16136 7380 16164
rect 3660 16124 3666 16136
rect 7374 16124 7380 16136
rect 7432 16124 7438 16176
rect 7742 16124 7748 16176
rect 7800 16164 7806 16176
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 7800 16136 8309 16164
rect 7800 16124 7806 16136
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 8297 16127 8355 16133
rect 8386 16124 8392 16176
rect 8444 16164 8450 16176
rect 10060 16164 10088 16195
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10192 16204 11529 16232
rect 10192 16192 10198 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11974 16232 11980 16244
rect 11935 16204 11980 16232
rect 11517 16195 11575 16201
rect 11974 16192 11980 16204
rect 12032 16232 12038 16244
rect 12434 16232 12440 16244
rect 12032 16204 12440 16232
rect 12032 16192 12038 16204
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 13722 16232 13728 16244
rect 13635 16204 13728 16232
rect 13722 16192 13728 16204
rect 13780 16232 13786 16244
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 13780 16204 14933 16232
rect 13780 16192 13786 16204
rect 14921 16201 14933 16204
rect 14967 16232 14979 16235
rect 15746 16232 15752 16244
rect 14967 16204 15752 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 12250 16164 12256 16176
rect 8444 16136 10088 16164
rect 10336 16136 12256 16164
rect 8444 16124 8450 16136
rect 10336 16108 10364 16136
rect 12250 16124 12256 16136
rect 12308 16164 12314 16176
rect 12713 16167 12771 16173
rect 12713 16164 12725 16167
rect 12308 16136 12725 16164
rect 12308 16124 12314 16136
rect 12713 16133 12725 16136
rect 12759 16133 12771 16167
rect 12713 16127 12771 16133
rect 12805 16167 12863 16173
rect 12805 16133 12817 16167
rect 12851 16164 12863 16167
rect 14458 16164 14464 16176
rect 12851 16136 14464 16164
rect 12851 16133 12863 16136
rect 12805 16127 12863 16133
rect 14458 16124 14464 16136
rect 14516 16124 14522 16176
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2682 16096 2688 16108
rect 2516 16068 2688 16096
rect 2516 16040 2544 16068
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2792 16068 3924 16096
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 16028 2467 16031
rect 2498 16028 2504 16040
rect 2455 16000 2504 16028
rect 2455 15997 2467 16000
rect 2409 15991 2467 15997
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2608 15892 2636 15991
rect 2792 15892 2820 16068
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 15997 2927 16031
rect 3896 16028 3924 16068
rect 4982 16056 4988 16108
rect 5040 16096 5046 16108
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 5040 16068 5089 16096
rect 5040 16056 5046 16068
rect 5077 16065 5089 16068
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 5905 16099 5963 16105
rect 5905 16065 5917 16099
rect 5951 16065 5963 16099
rect 5905 16059 5963 16065
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6454 16096 6460 16108
rect 6227 16068 6460 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 5920 16028 5948 16059
rect 6454 16056 6460 16068
rect 6512 16096 6518 16108
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 6512 16068 6653 16096
rect 6512 16056 6518 16068
rect 6641 16065 6653 16068
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16096 7159 16099
rect 7190 16096 7196 16108
rect 7147 16068 7196 16096
rect 7147 16065 7159 16068
rect 7101 16059 7159 16065
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 8168 16068 8217 16096
rect 8168 16056 8174 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 9217 16099 9275 16105
rect 8205 16059 8263 16065
rect 8312 16068 8524 16096
rect 6086 16028 6092 16040
rect 3896 16000 5120 16028
rect 5920 16000 6092 16028
rect 2869 15991 2927 15997
rect 2608 15864 2820 15892
rect 2884 15892 2912 15991
rect 5092 15972 5120 16000
rect 6086 15988 6092 16000
rect 6144 16028 6150 16040
rect 7834 16028 7840 16040
rect 6144 16000 7840 16028
rect 6144 15988 6150 16000
rect 7834 15988 7840 16000
rect 7892 16028 7898 16040
rect 8312 16028 8340 16068
rect 7892 16000 8340 16028
rect 8389 16031 8447 16037
rect 7892 15988 7898 16000
rect 8389 15997 8401 16031
rect 8435 15997 8447 16031
rect 8496 16028 8524 16068
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 9398 16096 9404 16108
rect 9263 16068 9404 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10229 16099 10287 16105
rect 9732 16068 9904 16096
rect 9732 16056 9738 16068
rect 9306 16028 9312 16040
rect 8496 16000 9312 16028
rect 8389 15991 8447 15997
rect 4430 15920 4436 15972
rect 4488 15960 4494 15972
rect 4614 15960 4620 15972
rect 4488 15932 4620 15960
rect 4488 15920 4494 15932
rect 4614 15920 4620 15932
rect 4672 15960 4678 15972
rect 4709 15963 4767 15969
rect 4709 15960 4721 15963
rect 4672 15932 4721 15960
rect 4672 15920 4678 15932
rect 4709 15929 4721 15932
rect 4755 15929 4767 15963
rect 4709 15923 4767 15929
rect 5074 15920 5080 15972
rect 5132 15920 5138 15972
rect 5810 15920 5816 15972
rect 5868 15960 5874 15972
rect 6457 15963 6515 15969
rect 6457 15960 6469 15963
rect 5868 15932 6469 15960
rect 5868 15920 5874 15932
rect 6457 15929 6469 15932
rect 6503 15929 6515 15963
rect 7469 15963 7527 15969
rect 6457 15923 6515 15929
rect 6564 15932 7328 15960
rect 4338 15892 4344 15904
rect 2884 15864 4344 15892
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4982 15892 4988 15904
rect 4943 15864 4988 15892
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6564 15892 6592 15932
rect 7190 15892 7196 15904
rect 6236 15864 6592 15892
rect 7151 15864 7196 15892
rect 6236 15852 6242 15864
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7300 15892 7328 15932
rect 7469 15929 7481 15963
rect 7515 15960 7527 15963
rect 7515 15932 7880 15960
rect 7515 15929 7527 15932
rect 7469 15923 7527 15929
rect 7742 15892 7748 15904
rect 7300 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 7852 15892 7880 15932
rect 8110 15920 8116 15972
rect 8168 15960 8174 15972
rect 8404 15960 8432 15991
rect 9306 15988 9312 16000
rect 9364 16028 9370 16040
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9364 16000 9781 16028
rect 9364 15988 9370 16000
rect 9769 15997 9781 16000
rect 9815 15997 9827 16031
rect 9876 16028 9904 16068
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10318 16096 10324 16108
rect 10275 16068 10324 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16096 11391 16099
rect 11698 16096 11704 16108
rect 11379 16068 11704 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 11882 16096 11888 16108
rect 11843 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12158 16056 12164 16108
rect 12216 16096 12222 16108
rect 13630 16096 13636 16108
rect 12216 16068 13032 16096
rect 13591 16068 13636 16096
rect 12216 16056 12222 16068
rect 9876 16000 11284 16028
rect 9769 15991 9827 15997
rect 8168 15932 8432 15960
rect 8168 15920 8174 15932
rect 9490 15920 9496 15972
rect 9548 15960 9554 15972
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 9548 15932 11161 15960
rect 9548 15920 9554 15932
rect 11149 15929 11161 15932
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 8294 15892 8300 15904
rect 7852 15864 8300 15892
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8444 15864 8677 15892
rect 8444 15852 8450 15864
rect 8665 15861 8677 15864
rect 8711 15892 8723 15895
rect 9674 15892 9680 15904
rect 8711 15864 9680 15892
rect 8711 15861 8723 15864
rect 8665 15855 8723 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 9766 15852 9772 15904
rect 9824 15892 9830 15904
rect 10318 15892 10324 15904
rect 9824 15864 10324 15892
rect 9824 15852 9830 15864
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11256 15892 11284 16000
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11572 16000 12081 16028
rect 11572 15988 11578 16000
rect 12069 15997 12081 16000
rect 12115 16028 12127 16031
rect 12342 16028 12348 16040
rect 12115 16000 12348 16028
rect 12115 15997 12127 16000
rect 12069 15991 12127 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 13004 16037 13032 16068
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14274 16096 14280 16108
rect 14235 16068 14280 16096
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 14599 16068 14780 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 16028 13047 16031
rect 13817 16031 13875 16037
rect 13035 16000 13400 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 13265 15963 13323 15969
rect 13265 15960 13277 15963
rect 12032 15932 13277 15960
rect 12032 15920 12038 15932
rect 13265 15929 13277 15932
rect 13311 15929 13323 15963
rect 13372 15960 13400 16000
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13832 15960 13860 15991
rect 14752 15969 14780 16068
rect 13372 15932 13860 15960
rect 14737 15963 14795 15969
rect 13265 15923 13323 15929
rect 14737 15929 14749 15963
rect 14783 15960 14795 15963
rect 16022 15960 16028 15972
rect 14783 15932 16028 15960
rect 14783 15929 14795 15932
rect 14737 15923 14795 15929
rect 16022 15920 16028 15932
rect 16080 15920 16086 15972
rect 11514 15892 11520 15904
rect 11256 15864 11520 15892
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 11848 15864 12357 15892
rect 11848 15852 11854 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12345 15855 12403 15861
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 15930 15892 15936 15904
rect 12584 15864 15936 15892
rect 12584 15852 12590 15864
rect 15930 15852 15936 15864
rect 15988 15852 15994 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 2774 15688 2780 15700
rect 2372 15660 2780 15688
rect 2372 15648 2378 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 6178 15688 6184 15700
rect 2915 15660 6184 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 2038 15512 2044 15564
rect 2096 15552 2102 15564
rect 3145 15555 3203 15561
rect 3145 15552 3157 15555
rect 2096 15524 3157 15552
rect 2096 15512 2102 15524
rect 3145 15521 3157 15524
rect 3191 15521 3203 15555
rect 3145 15515 3203 15521
rect 2406 15484 2412 15496
rect 2367 15456 2412 15484
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 3252 15484 3280 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 10686 15688 10692 15700
rect 6972 15660 10692 15688
rect 6972 15648 6978 15660
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 12308 15660 12353 15688
rect 12308 15648 12314 15660
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12710 15688 12716 15700
rect 12492 15660 12537 15688
rect 12671 15660 12716 15688
rect 12492 15648 12498 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 13814 15688 13820 15700
rect 13679 15660 13820 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13814 15648 13820 15660
rect 13872 15688 13878 15700
rect 14458 15688 14464 15700
rect 13872 15660 14464 15688
rect 13872 15648 13878 15660
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 11517 15623 11575 15629
rect 11517 15589 11529 15623
rect 11563 15620 11575 15623
rect 11698 15620 11704 15632
rect 11563 15592 11704 15620
rect 11563 15589 11575 15592
rect 11517 15583 11575 15589
rect 11698 15580 11704 15592
rect 11756 15620 11762 15632
rect 14826 15620 14832 15632
rect 11756 15592 14832 15620
rect 11756 15580 11762 15592
rect 14826 15580 14832 15592
rect 14884 15580 14890 15632
rect 4154 15552 4160 15564
rect 2556 15456 3280 15484
rect 3344 15524 4160 15552
rect 2556 15444 2562 15456
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 2133 15419 2191 15425
rect 2133 15416 2145 15419
rect 1452 15388 2145 15416
rect 1452 15376 1458 15388
rect 2133 15385 2145 15388
rect 2179 15385 2191 15419
rect 2133 15379 2191 15385
rect 2774 15376 2780 15428
rect 2832 15416 2838 15428
rect 3053 15419 3111 15425
rect 3053 15416 3065 15419
rect 2832 15388 3065 15416
rect 2832 15376 2838 15388
rect 3053 15385 3065 15388
rect 3099 15416 3111 15419
rect 3344 15416 3372 15524
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 11882 15552 11888 15564
rect 11843 15524 11888 15552
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 13044 15524 13277 15552
rect 13044 15512 13050 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 13630 15512 13636 15564
rect 13688 15552 13694 15564
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 13688 15524 13737 15552
rect 13688 15512 13694 15524
rect 13725 15521 13737 15524
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4338 15484 4344 15496
rect 4295 15456 4344 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4338 15444 4344 15456
rect 4396 15484 4402 15496
rect 5534 15484 5540 15496
rect 4396 15456 5540 15484
rect 4396 15444 4402 15456
rect 5534 15444 5540 15456
rect 5592 15484 5598 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5592 15456 5733 15484
rect 5592 15444 5598 15456
rect 5721 15453 5733 15456
rect 5767 15484 5779 15487
rect 6178 15484 6184 15496
rect 5767 15456 6184 15484
rect 5767 15453 5779 15456
rect 5721 15447 5779 15453
rect 6178 15444 6184 15456
rect 6236 15484 6242 15496
rect 7190 15484 7196 15496
rect 6236 15456 7196 15484
rect 6236 15444 6242 15456
rect 7190 15444 7196 15456
rect 7248 15484 7254 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7248 15456 7297 15484
rect 7248 15444 7254 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8757 15487 8815 15493
rect 8757 15484 8769 15487
rect 8260 15456 8769 15484
rect 8260 15444 8266 15456
rect 8757 15453 8769 15456
rect 8803 15484 8815 15487
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8803 15456 9137 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9125 15453 9137 15456
rect 9171 15484 9183 15487
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 9171 15456 9321 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 12158 15484 12164 15496
rect 11388 15456 12164 15484
rect 11388 15444 11394 15456
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13354 15484 13360 15496
rect 13127 15456 13360 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 3099 15388 3372 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 4494 15419 4552 15425
rect 4494 15416 4506 15419
rect 4212 15388 4506 15416
rect 4212 15376 4218 15388
rect 4494 15385 4506 15388
rect 4540 15385 4552 15419
rect 7018 15419 7076 15425
rect 7018 15416 7030 15419
rect 4494 15379 4552 15385
rect 5828 15388 7030 15416
rect 5828 15360 5856 15388
rect 7018 15385 7030 15388
rect 7064 15385 7076 15419
rect 7018 15379 7076 15385
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 8490 15419 8548 15425
rect 8490 15416 8502 15419
rect 8352 15388 8502 15416
rect 8352 15376 8358 15388
rect 8490 15385 8502 15388
rect 8536 15385 8548 15419
rect 8490 15379 8548 15385
rect 9490 15376 9496 15428
rect 9548 15425 9554 15428
rect 9548 15419 9612 15425
rect 9548 15385 9566 15419
rect 9600 15385 9612 15419
rect 9548 15379 9612 15385
rect 13173 15419 13231 15425
rect 13173 15385 13185 15419
rect 13219 15416 13231 15419
rect 13906 15416 13912 15428
rect 13219 15388 13912 15416
rect 13219 15385 13231 15388
rect 13173 15379 13231 15385
rect 9548 15376 9554 15379
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 290 15308 296 15360
rect 348 15348 354 15360
rect 2314 15348 2320 15360
rect 348 15320 2320 15348
rect 348 15308 354 15320
rect 2314 15308 2320 15320
rect 2372 15308 2378 15360
rect 2498 15348 2504 15360
rect 2459 15320 2504 15348
rect 2498 15308 2504 15320
rect 2556 15348 2562 15360
rect 2682 15348 2688 15360
rect 2556 15320 2688 15348
rect 2556 15308 2562 15320
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 5166 15348 5172 15360
rect 4120 15320 5172 15348
rect 4120 15308 4126 15320
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5629 15351 5687 15357
rect 5629 15317 5641 15351
rect 5675 15348 5687 15351
rect 5810 15348 5816 15360
rect 5675 15320 5816 15348
rect 5675 15317 5687 15320
rect 5629 15311 5687 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 5905 15351 5963 15357
rect 5905 15317 5917 15351
rect 5951 15348 5963 15351
rect 5994 15348 6000 15360
rect 5951 15320 6000 15348
rect 5951 15317 5963 15320
rect 5905 15311 5963 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 7377 15351 7435 15357
rect 7377 15317 7389 15351
rect 7423 15348 7435 15351
rect 7466 15348 7472 15360
rect 7423 15320 7472 15348
rect 7423 15317 7435 15320
rect 7377 15311 7435 15317
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 10689 15351 10747 15357
rect 10689 15317 10701 15351
rect 10735 15348 10747 15351
rect 10962 15348 10968 15360
rect 10735 15320 10968 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 1673 15147 1731 15153
rect 1673 15113 1685 15147
rect 1719 15144 1731 15147
rect 1946 15144 1952 15156
rect 1719 15116 1952 15144
rect 1719 15113 1731 15116
rect 1673 15107 1731 15113
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 2590 15104 2596 15156
rect 2648 15144 2654 15156
rect 4338 15144 4344 15156
rect 2648 15116 4200 15144
rect 4299 15116 4344 15144
rect 2648 15104 2654 15116
rect 2406 15076 2412 15088
rect 2367 15048 2412 15076
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 4062 15076 4068 15088
rect 2700 15048 4068 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2498 15008 2504 15020
rect 1811 14980 2504 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 2700 15017 2728 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 3982 15011 4040 15017
rect 3982 15008 3994 15011
rect 3660 14980 3994 15008
rect 3660 14968 3666 14980
rect 3982 14977 3994 14980
rect 4028 14977 4040 15011
rect 3982 14971 4040 14977
rect 1578 14940 1584 14952
rect 1539 14912 1584 14940
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 4172 14940 4200 15116
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 4448 15116 12909 15144
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 4356 15008 4384 15104
rect 4295 14980 4384 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4448 14940 4476 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 12897 15107 12955 15113
rect 13538 15104 13544 15156
rect 13596 15144 13602 15156
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 13596 15116 14013 15144
rect 13596 15104 13602 15116
rect 14001 15113 14013 15116
rect 14047 15113 14059 15147
rect 15654 15144 15660 15156
rect 15567 15116 15660 15144
rect 14001 15107 14059 15113
rect 15654 15104 15660 15116
rect 15712 15144 15718 15156
rect 16850 15144 16856 15156
rect 15712 15116 16856 15144
rect 15712 15104 15718 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 5994 15085 6000 15088
rect 5936 15079 6000 15085
rect 5936 15045 5948 15079
rect 5982 15045 6000 15079
rect 5936 15039 6000 15045
rect 5994 15036 6000 15039
rect 6052 15036 6058 15088
rect 6104 15048 7328 15076
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 6104 15008 6132 15048
rect 5408 14980 6132 15008
rect 5408 14968 5414 14980
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 6236 14980 6377 15008
rect 6236 14968 6242 14980
rect 6365 14977 6377 14980
rect 6411 15008 6423 15011
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6411 14980 6561 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6816 15011 6874 15017
rect 6816 14977 6828 15011
rect 6862 15008 6874 15011
rect 7190 15008 7196 15020
rect 6862 14980 7196 15008
rect 6862 14977 6874 14980
rect 6816 14971 6874 14977
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7300 15008 7328 15048
rect 7466 15036 7472 15088
rect 7524 15076 7530 15088
rect 8358 15079 8416 15085
rect 8358 15076 8370 15079
rect 7524 15048 8370 15076
rect 7524 15036 7530 15048
rect 8358 15045 8370 15048
rect 8404 15045 8416 15079
rect 8358 15039 8416 15045
rect 10318 15036 10324 15088
rect 10376 15076 10382 15088
rect 11790 15076 11796 15088
rect 10376 15048 11652 15076
rect 11751 15048 11796 15076
rect 10376 15036 10382 15048
rect 8113 15011 8171 15017
rect 7300 14980 8064 15008
rect 4172 14912 4476 14940
rect 2682 14832 2688 14884
rect 2740 14872 2746 14884
rect 2740 14844 3372 14872
rect 2740 14832 2746 14844
rect 2130 14804 2136 14816
rect 2091 14776 2136 14804
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 2869 14807 2927 14813
rect 2869 14773 2881 14807
rect 2915 14804 2927 14807
rect 3142 14804 3148 14816
rect 2915 14776 3148 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 3344 14804 3372 14844
rect 4801 14807 4859 14813
rect 4801 14804 4813 14807
rect 3344 14776 4813 14804
rect 4801 14773 4813 14776
rect 4847 14773 4859 14807
rect 7926 14804 7932 14816
rect 7887 14776 7932 14804
rect 4801 14767 4859 14773
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 8036 14804 8064 14980
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8202 15008 8208 15020
rect 8159 14980 8208 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 10686 14968 10692 15020
rect 10744 15017 10750 15020
rect 10744 15008 10756 15017
rect 10744 14980 10789 15008
rect 10744 14971 10756 14980
rect 10744 14968 10750 14971
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10928 14980 10977 15008
rect 10928 14968 10934 14980
rect 10965 14977 10977 14980
rect 11011 15008 11023 15011
rect 11057 15011 11115 15017
rect 11057 15008 11069 15011
rect 11011 14980 11069 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11057 14977 11069 14980
rect 11103 14977 11115 15011
rect 11624 15008 11652 15048
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 11885 15079 11943 15085
rect 11885 15045 11897 15079
rect 11931 15076 11943 15079
rect 11974 15076 11980 15088
rect 11931 15048 11980 15076
rect 11931 15045 11943 15048
rect 11885 15039 11943 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 13096 15048 13400 15076
rect 13096 15008 13124 15048
rect 13262 15008 13268 15020
rect 11624 14980 13124 15008
rect 13223 14980 13268 15008
rect 11057 14971 11115 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13372 15008 13400 15048
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 13630 15076 13636 15088
rect 13504 15048 13636 15076
rect 13504 15036 13510 15048
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 13372 14980 14473 15008
rect 14461 14977 14473 14980
rect 14507 15008 14519 15011
rect 14642 15008 14648 15020
rect 14507 14980 14648 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 11701 14943 11759 14949
rect 9140 14912 9628 14940
rect 9140 14804 9168 14912
rect 8036 14776 9168 14804
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9600 14813 9628 14912
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 11882 14940 11888 14952
rect 11747 14912 11888 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 13136 14912 13369 14940
rect 13136 14900 13142 14912
rect 13357 14909 13369 14912
rect 13403 14909 13415 14943
rect 13357 14903 13415 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 16298 14940 16304 14952
rect 13587 14912 16304 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 11020 14844 12817 14872
rect 11020 14832 11026 14844
rect 12805 14841 12817 14844
rect 12851 14872 12863 14875
rect 13556 14872 13584 14903
rect 16298 14900 16304 14912
rect 16356 14900 16362 14952
rect 12851 14844 13584 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 9493 14807 9551 14813
rect 9493 14804 9505 14807
rect 9364 14776 9505 14804
rect 9364 14764 9370 14776
rect 9493 14773 9505 14776
rect 9539 14773 9551 14807
rect 9493 14767 9551 14773
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14773 9643 14807
rect 9585 14767 9643 14773
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 12618 14804 12624 14816
rect 12299 14776 12624 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13814 14804 13820 14816
rect 12768 14776 13820 14804
rect 12768 14764 12774 14776
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 14737 14807 14795 14813
rect 14737 14773 14749 14807
rect 14783 14804 14795 14807
rect 15010 14804 15016 14816
rect 14783 14776 15016 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 3881 14603 3939 14609
rect 3881 14600 3893 14603
rect 2924 14572 3893 14600
rect 2924 14560 2930 14572
rect 3881 14569 3893 14572
rect 3927 14600 3939 14603
rect 4062 14600 4068 14612
rect 3927 14572 4068 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4062 14560 4068 14572
rect 4120 14600 4126 14612
rect 4338 14600 4344 14612
rect 4120 14572 4344 14600
rect 4120 14560 4126 14572
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 5500 14572 7297 14600
rect 5500 14560 5506 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 9306 14600 9312 14612
rect 7285 14563 7343 14569
rect 7668 14572 9312 14600
rect 7668 14464 7696 14572
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 13078 14600 13084 14612
rect 9548 14572 12434 14600
rect 13039 14572 13084 14600
rect 9548 14560 9554 14572
rect 6748 14436 7696 14464
rect 1946 14356 1952 14408
rect 2004 14396 2010 14408
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 2004 14368 2237 14396
rect 2004 14356 2010 14368
rect 2225 14365 2237 14368
rect 2271 14396 2283 14399
rect 2866 14396 2872 14408
rect 2271 14368 2872 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 6569 14399 6627 14405
rect 6569 14365 6581 14399
rect 6615 14396 6627 14399
rect 6748 14396 6776 14436
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 11882 14464 11888 14476
rect 8996 14436 9628 14464
rect 11795 14436 11888 14464
rect 8996 14424 9002 14436
rect 6615 14368 6776 14396
rect 6615 14365 6627 14368
rect 6569 14359 6627 14365
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 6880 14368 6929 14396
rect 6880 14356 6886 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 1762 14288 1768 14340
rect 1820 14328 1826 14340
rect 2470 14331 2528 14337
rect 2470 14328 2482 14331
rect 1820 14300 2482 14328
rect 1820 14288 1826 14300
rect 2470 14297 2482 14300
rect 2516 14328 2528 14331
rect 2682 14328 2688 14340
rect 2516 14300 2688 14328
rect 2516 14297 2528 14300
rect 2470 14291 2528 14297
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 3602 14260 3608 14272
rect 3563 14232 3608 14260
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 5350 14260 5356 14272
rect 4212 14232 5356 14260
rect 4212 14220 4218 14232
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5810 14260 5816 14272
rect 5491 14232 5816 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6932 14260 6960 14359
rect 7098 14356 7104 14408
rect 7156 14356 7162 14408
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8220 14368 8677 14396
rect 7116 14328 7144 14356
rect 8220 14340 8248 14368
rect 8665 14365 8677 14368
rect 8711 14396 8723 14399
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8711 14368 9321 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 9309 14365 9321 14368
rect 9355 14396 9367 14399
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 9355 14368 9505 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 9600 14396 9628 14436
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12406 14464 12434 14572
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13320 14572 14105 14600
rect 13320 14560 13326 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 12989 14535 13047 14541
rect 12989 14532 13001 14535
rect 12952 14504 13001 14532
rect 12952 14492 12958 14504
rect 12989 14501 13001 14504
rect 13035 14532 13047 14535
rect 13446 14532 13452 14544
rect 13035 14504 13452 14532
rect 13035 14501 13047 14504
rect 12989 14495 13047 14501
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 13633 14467 13691 14473
rect 13633 14464 13645 14467
rect 12406 14436 13645 14464
rect 13633 14433 13645 14436
rect 13679 14464 13691 14467
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 13679 14436 14657 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 15252 14436 15485 14464
rect 15252 14424 15258 14436
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 11900 14396 11928 14424
rect 9600 14368 11928 14396
rect 15381 14399 15439 14405
rect 9493 14359 9551 14365
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15654 14396 15660 14408
rect 15427 14368 15660 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 7926 14328 7932 14340
rect 7116 14300 7932 14328
rect 7926 14288 7932 14300
rect 7984 14328 7990 14340
rect 7984 14300 8156 14328
rect 7984 14288 7990 14300
rect 7101 14263 7159 14269
rect 7101 14260 7113 14263
rect 6932 14232 7113 14260
rect 7101 14229 7113 14232
rect 7147 14229 7159 14263
rect 8128 14260 8156 14300
rect 8202 14288 8208 14340
rect 8260 14288 8266 14340
rect 8398 14331 8456 14337
rect 8398 14328 8410 14331
rect 8312 14300 8410 14328
rect 8312 14260 8340 14300
rect 8398 14297 8410 14300
rect 8444 14297 8456 14331
rect 8398 14291 8456 14297
rect 8128 14232 8340 14260
rect 9508 14260 9536 14359
rect 15488 14340 15516 14368
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 9738 14331 9796 14337
rect 9738 14328 9750 14331
rect 9640 14300 9750 14328
rect 9640 14288 9646 14300
rect 9738 14297 9750 14300
rect 9784 14297 9796 14331
rect 9738 14291 9796 14297
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 11940 14300 12173 14328
rect 11940 14288 11946 14300
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12161 14291 12219 14297
rect 13449 14331 13507 14337
rect 13449 14297 13461 14331
rect 13495 14328 13507 14331
rect 13814 14328 13820 14340
rect 13495 14300 13820 14328
rect 13495 14297 13507 14300
rect 13449 14291 13507 14297
rect 13814 14288 13820 14300
rect 13872 14288 13878 14340
rect 14461 14331 14519 14337
rect 14461 14297 14473 14331
rect 14507 14328 14519 14331
rect 14507 14300 14964 14328
rect 14507 14297 14519 14300
rect 14461 14291 14519 14297
rect 9858 14260 9864 14272
rect 9508 14232 9864 14260
rect 7101 14223 7159 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10744 14232 10885 14260
rect 10744 14220 10750 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 12066 14260 12072 14272
rect 12027 14232 12072 14260
rect 10873 14223 10931 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12802 14260 12808 14272
rect 12575 14232 12808 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13541 14263 13599 14269
rect 13541 14260 13553 14263
rect 13320 14232 13553 14260
rect 13320 14220 13326 14232
rect 13541 14229 13553 14232
rect 13587 14229 13599 14263
rect 14550 14260 14556 14272
rect 14511 14232 14556 14260
rect 13541 14223 13599 14229
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 14936 14269 14964 14300
rect 15470 14288 15476 14340
rect 15528 14288 15534 14340
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14229 14979 14263
rect 15286 14260 15292 14272
rect 15247 14232 15292 14260
rect 14921 14223 14979 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4304 14028 4721 14056
rect 4304 14016 4310 14028
rect 4709 14025 4721 14028
rect 4755 14056 4767 14059
rect 5074 14056 5080 14068
rect 4755 14028 5080 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9398 14056 9404 14068
rect 9180 14028 9404 14056
rect 9180 14016 9186 14028
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 9548 14028 9597 14056
rect 9548 14016 9554 14028
rect 9585 14025 9597 14028
rect 9631 14025 9643 14059
rect 9585 14019 9643 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 11664 14028 11897 14056
rect 11664 14016 11670 14028
rect 11885 14025 11897 14028
rect 11931 14056 11943 14059
rect 12250 14056 12256 14068
rect 11931 14028 12256 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14025 12403 14059
rect 12802 14056 12808 14068
rect 12763 14028 12808 14056
rect 12345 14019 12403 14025
rect 2866 13988 2872 14000
rect 2792 13960 2872 13988
rect 2792 13929 2820 13960
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 3044 13991 3102 13997
rect 3044 13957 3056 13991
rect 3090 13988 3102 13991
rect 3510 13988 3516 14000
rect 3090 13960 3516 13988
rect 3090 13957 3102 13960
rect 3044 13951 3102 13957
rect 3510 13948 3516 13960
rect 3568 13948 3574 14000
rect 12360 13988 12388 14019
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 13630 14056 13636 14068
rect 13320 14028 13636 14056
rect 13320 14016 13326 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13964 14028 14013 14056
rect 13964 14016 13970 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14001 14019 14059 14025
rect 14461 14059 14519 14065
rect 14461 14025 14473 14059
rect 14507 14056 14519 14059
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 14507 14028 14841 14056
rect 14507 14025 14519 14028
rect 14461 14019 14519 14025
rect 14829 14025 14841 14028
rect 14875 14025 14887 14059
rect 14829 14019 14887 14025
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15289 14059 15347 14065
rect 15289 14056 15301 14059
rect 15068 14028 15301 14056
rect 15068 14016 15074 14028
rect 15289 14025 15301 14028
rect 15335 14056 15347 14059
rect 15746 14056 15752 14068
rect 15335 14028 15752 14056
rect 15335 14025 15347 14028
rect 15289 14019 15347 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 8312 13960 12388 13988
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 2884 13892 3832 13920
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 1964 13852 1992 13883
rect 2884 13852 2912 13892
rect 1964 13824 2912 13852
rect 3804 13852 3832 13892
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 4120 13892 4261 13920
rect 4120 13880 4126 13892
rect 4249 13889 4261 13892
rect 4295 13920 4307 13923
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4295 13892 4905 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 4893 13889 4905 13892
rect 4939 13920 4951 13923
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 4939 13892 5641 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5629 13889 5641 13892
rect 5675 13920 5687 13923
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5675 13892 5825 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 5902 13920 5908 13932
rect 5859 13892 5908 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 5902 13880 5908 13892
rect 5960 13920 5966 13932
rect 6822 13920 6828 13932
rect 5960 13892 6828 13920
rect 5960 13880 5966 13892
rect 6822 13880 6828 13892
rect 6880 13920 6886 13932
rect 6917 13923 6975 13929
rect 6917 13920 6929 13923
rect 6880 13892 6929 13920
rect 6880 13880 6886 13892
rect 6917 13889 6929 13892
rect 6963 13920 6975 13923
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6963 13892 7205 13920
rect 6963 13889 6975 13892
rect 6917 13883 6975 13889
rect 7193 13889 7205 13892
rect 7239 13920 7251 13923
rect 7374 13920 7380 13932
rect 7239 13892 7380 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7374 13880 7380 13892
rect 7432 13920 7438 13932
rect 8021 13923 8079 13929
rect 8021 13920 8033 13923
rect 7432 13892 8033 13920
rect 7432 13880 7438 13892
rect 8021 13889 8033 13892
rect 8067 13920 8079 13923
rect 8202 13920 8208 13932
rect 8067 13892 8208 13920
rect 8067 13889 8079 13892
rect 8021 13883 8079 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8312 13852 8340 13960
rect 12618 13948 12624 14000
rect 12676 13988 12682 14000
rect 12713 13991 12771 13997
rect 12713 13988 12725 13991
rect 12676 13960 12725 13988
rect 12676 13948 12682 13960
rect 12713 13957 12725 13960
rect 12759 13957 12771 13991
rect 12713 13951 12771 13957
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 14642 13988 14648 14000
rect 13136 13960 14648 13988
rect 13136 13948 13142 13960
rect 14642 13948 14648 13960
rect 14700 13988 14706 14000
rect 15197 13991 15255 13997
rect 15197 13988 15209 13991
rect 14700 13960 15209 13988
rect 14700 13948 14706 13960
rect 15197 13957 15209 13960
rect 15243 13957 15255 13991
rect 15197 13951 15255 13957
rect 8472 13923 8530 13929
rect 8472 13889 8484 13923
rect 8518 13920 8530 13923
rect 8846 13920 8852 13932
rect 8518 13892 8852 13920
rect 8518 13889 8530 13892
rect 8472 13883 8530 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 11146 13920 11152 13932
rect 9364 13892 11152 13920
rect 9364 13880 9370 13892
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12584 13892 13032 13920
rect 12584 13880 12590 13892
rect 3804 13824 8340 13852
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 11112 13824 11253 13852
rect 11112 13812 11118 13824
rect 11241 13821 11253 13824
rect 11287 13852 11299 13855
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11287 13824 11989 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 13004 13852 13032 13892
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13504 13892 13553 13920
rect 13504 13880 13510 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 13964 13892 14381 13920
rect 13964 13880 13970 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 14516 13892 15424 13920
rect 14516 13880 14522 13892
rect 15396 13861 15424 13892
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13004 13824 13737 13852
rect 12897 13815 12955 13821
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 15381 13855 15439 13861
rect 15381 13821 15393 13855
rect 15427 13821 15439 13855
rect 15381 13815 15439 13821
rect 6178 13784 6184 13796
rect 4356 13756 6184 13784
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 4356 13716 4384 13756
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 9824 13756 11744 13784
rect 9824 13744 9830 13756
rect 3568 13688 4384 13716
rect 3568 13676 3574 13688
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 6270 13716 6276 13728
rect 4488 13688 6276 13716
rect 4488 13676 4494 13688
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 11514 13716 11520 13728
rect 11475 13688 11520 13716
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11716 13716 11744 13756
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12084 13784 12112 13815
rect 12912 13784 12940 13815
rect 11848 13756 12112 13784
rect 12406 13756 12940 13784
rect 11848 13744 11854 13756
rect 12406 13716 12434 13756
rect 11716 13688 12434 13716
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 14568 13716 14596 13815
rect 13780 13688 14596 13716
rect 13780 13676 13786 13688
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 5258 13512 5264 13524
rect 4212 13484 5264 13512
rect 4212 13472 4218 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 7190 13512 7196 13524
rect 7151 13484 7196 13512
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7558 13472 7564 13524
rect 7616 13512 7622 13524
rect 11882 13512 11888 13524
rect 7616 13484 11284 13512
rect 11843 13484 11888 13512
rect 7616 13472 7622 13484
rect 8757 13447 8815 13453
rect 8757 13413 8769 13447
rect 8803 13444 8815 13447
rect 8938 13444 8944 13456
rect 8803 13416 8944 13444
rect 8803 13413 8815 13416
rect 8757 13407 8815 13413
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 11054 13444 11060 13456
rect 11015 13416 11060 13444
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 1765 13379 1823 13385
rect 1765 13376 1777 13379
rect 1636 13348 1777 13376
rect 1636 13336 1642 13348
rect 1765 13345 1777 13348
rect 1811 13376 1823 13379
rect 2590 13376 2596 13388
rect 1811 13348 2596 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4246 13376 4252 13388
rect 4120 13348 4252 13376
rect 4120 13336 4126 13348
rect 4246 13336 4252 13348
rect 4304 13376 4310 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 4304 13348 4353 13376
rect 4304 13336 4310 13348
rect 4341 13345 4353 13348
rect 4387 13345 4399 13379
rect 7374 13376 7380 13388
rect 7335 13348 7380 13376
rect 4341 13339 4399 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 11256 13385 11284 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 12032 13484 13185 13512
rect 12032 13472 12038 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13630 13512 13636 13524
rect 13412 13484 13636 13512
rect 13412 13472 13418 13484
rect 13630 13472 13636 13484
rect 13688 13512 13694 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 13688 13484 14289 13512
rect 13688 13472 13694 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 14645 13515 14703 13521
rect 14645 13512 14657 13515
rect 14608 13484 14657 13512
rect 14608 13472 14614 13484
rect 14645 13481 14657 13484
rect 14691 13481 14703 13515
rect 14645 13475 14703 13481
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11330 13376 11336 13388
rect 11287 13348 11336 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13376 11483 13379
rect 11514 13376 11520 13388
rect 11471 13348 11520 13376
rect 11471 13345 11483 13348
rect 11425 13339 11483 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 13722 13376 13728 13388
rect 13412 13348 13728 13376
rect 13412 13336 13418 13348
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 14090 13376 14096 13388
rect 14051 13348 14096 13376
rect 14090 13336 14096 13348
rect 14148 13376 14154 13388
rect 14734 13376 14740 13388
rect 14148 13348 14740 13376
rect 14148 13336 14154 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15194 13376 15200 13388
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 15344 13348 15485 13376
rect 15344 13336 15350 13348
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 1995 13280 2513 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2501 13277 2513 13280
rect 2547 13308 2559 13311
rect 2682 13308 2688 13320
rect 2547 13280 2688 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2682 13268 2688 13280
rect 2740 13308 2746 13320
rect 3694 13308 3700 13320
rect 2740 13280 3700 13308
rect 2740 13268 2746 13280
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 4608 13311 4666 13317
rect 4608 13277 4620 13311
rect 4654 13277 4666 13311
rect 4608 13271 4666 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13308 5871 13311
rect 5902 13308 5908 13320
rect 5859 13280 5908 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 1857 13243 1915 13249
rect 1857 13209 1869 13243
rect 1903 13240 1915 13243
rect 1903 13212 2728 13240
rect 1903 13209 1915 13212
rect 1857 13203 1915 13209
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2700 13181 2728 13212
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 4632 13240 4660 13271
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7633 13311 7691 13317
rect 7633 13308 7645 13311
rect 7340 13280 7645 13308
rect 7340 13268 7346 13280
rect 7633 13277 7645 13280
rect 7679 13277 7691 13311
rect 7633 13271 7691 13277
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 9125 13311 9183 13317
rect 7984 13280 8984 13308
rect 7984 13268 7990 13280
rect 4580 13212 4660 13240
rect 6080 13243 6138 13249
rect 4580 13200 4586 13212
rect 6080 13209 6092 13243
rect 6126 13240 6138 13243
rect 7098 13240 7104 13252
rect 6126 13212 7104 13240
rect 6126 13209 6138 13212
rect 6080 13203 6138 13209
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 8846 13240 8852 13252
rect 8680 13212 8852 13240
rect 2685 13175 2743 13181
rect 2685 13141 2697 13175
rect 2731 13172 2743 13175
rect 4430 13172 4436 13184
rect 2731 13144 4436 13172
rect 2731 13141 2743 13144
rect 2685 13135 2743 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 5721 13175 5779 13181
rect 5721 13141 5733 13175
rect 5767 13172 5779 13175
rect 8680 13172 8708 13212
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 5767 13144 8708 13172
rect 8956 13172 8984 13280
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9858 13308 9864 13320
rect 9171 13280 9864 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 9858 13268 9864 13280
rect 9916 13308 9922 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 9916 13280 10609 13308
rect 9916 13268 9922 13280
rect 10597 13277 10609 13280
rect 10643 13308 10655 13311
rect 10870 13308 10876 13320
rect 10643 13280 10876 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12952 13280 13093 13308
rect 12952 13268 12958 13280
rect 13081 13277 13093 13280
rect 13127 13308 13139 13311
rect 13541 13311 13599 13317
rect 13541 13308 13553 13311
rect 13127 13280 13553 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13541 13277 13553 13280
rect 13587 13308 13599 13311
rect 13998 13308 14004 13320
rect 13587 13280 14004 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 13998 13268 14004 13280
rect 14056 13268 14062 13320
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15378 13308 15384 13320
rect 15151 13280 15384 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 10042 13200 10048 13252
rect 10100 13240 10106 13252
rect 10330 13243 10388 13249
rect 10330 13240 10342 13243
rect 10100 13212 10342 13240
rect 10100 13200 10106 13212
rect 10330 13209 10342 13212
rect 10376 13209 10388 13243
rect 10330 13203 10388 13209
rect 11422 13200 11428 13252
rect 11480 13240 11486 13252
rect 11698 13240 11704 13252
rect 11480 13212 11704 13240
rect 11480 13200 11486 13212
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 9217 13175 9275 13181
rect 9217 13172 9229 13175
rect 8956 13144 9229 13172
rect 5767 13141 5779 13144
rect 5721 13135 5779 13141
rect 9217 13141 9229 13144
rect 9263 13141 9275 13175
rect 9217 13135 9275 13141
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11112 13144 11529 13172
rect 11112 13132 11118 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 11606 13132 11612 13184
rect 11664 13172 11670 13184
rect 11790 13172 11796 13184
rect 11664 13144 11796 13172
rect 11664 13132 11670 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12250 13172 12256 13184
rect 12032 13144 12256 13172
rect 12032 13132 12038 13144
rect 12250 13132 12256 13144
rect 12308 13172 12314 13184
rect 12437 13175 12495 13181
rect 12437 13172 12449 13175
rect 12308 13144 12449 13172
rect 12308 13132 12314 13144
rect 12437 13141 12449 13144
rect 12483 13141 12495 13175
rect 12437 13135 12495 13141
rect 13630 13132 13636 13184
rect 13688 13172 13694 13184
rect 13688 13144 13733 13172
rect 13688 13132 13694 13144
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 13964 13144 14473 13172
rect 13964 13132 13970 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15010 13172 15016 13184
rect 14884 13144 15016 13172
rect 14884 13132 14890 13144
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 3329 12971 3387 12977
rect 3329 12937 3341 12971
rect 3375 12968 3387 12971
rect 4062 12968 4068 12980
rect 3375 12940 4068 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 4798 12968 4804 12980
rect 4304 12940 4804 12968
rect 4304 12928 4310 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5902 12968 5908 12980
rect 5552 12940 5908 12968
rect 5552 12900 5580 12940
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 10134 12968 10140 12980
rect 8772 12940 10140 12968
rect 8772 12900 8800 12940
rect 10134 12928 10140 12940
rect 10192 12968 10198 12980
rect 11422 12968 11428 12980
rect 10192 12940 11428 12968
rect 10192 12928 10198 12940
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11756 12940 11897 12968
rect 11756 12928 11762 12940
rect 11885 12937 11897 12940
rect 11931 12968 11943 12971
rect 12345 12971 12403 12977
rect 12345 12968 12357 12971
rect 11931 12940 12357 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12345 12937 12357 12940
rect 12391 12937 12403 12971
rect 12345 12931 12403 12937
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 13538 12968 13544 12980
rect 13403 12940 13544 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 13872 12940 14289 12968
rect 13872 12928 13878 12940
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 14277 12931 14335 12937
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15378 12968 15384 12980
rect 15252 12940 15384 12968
rect 15252 12928 15258 12940
rect 15378 12928 15384 12940
rect 15436 12968 15442 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 15436 12940 15485 12968
rect 15436 12928 15442 12940
rect 15473 12937 15485 12940
rect 15519 12937 15531 12971
rect 15473 12931 15531 12937
rect 2746 12872 5580 12900
rect 6656 12872 8800 12900
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2216 12835 2274 12841
rect 2216 12801 2228 12835
rect 2262 12832 2274 12835
rect 2746 12832 2774 12872
rect 2262 12804 2774 12832
rect 2262 12801 2274 12804
rect 2216 12795 2274 12801
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4534 12835 4592 12841
rect 4534 12832 4546 12835
rect 4212 12804 4546 12832
rect 4212 12792 4218 12804
rect 4534 12801 4546 12804
rect 4580 12832 4592 12835
rect 4706 12832 4712 12844
rect 4580 12804 4712 12832
rect 4580 12801 4592 12804
rect 4534 12795 4592 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5074 12832 5080 12844
rect 4856 12804 4901 12832
rect 5035 12804 5080 12832
rect 4856 12792 4862 12804
rect 5074 12792 5080 12804
rect 5132 12832 5138 12844
rect 6086 12832 6092 12844
rect 5132 12804 6092 12832
rect 5132 12792 5138 12804
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6187 12804 6377 12832
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 4816 12764 4844 12792
rect 5166 12764 5172 12776
rect 4816 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12764 5230 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 5224 12736 5273 12764
rect 5224 12724 5230 12736
rect 5261 12733 5273 12736
rect 5307 12764 5319 12767
rect 5997 12767 6055 12773
rect 5997 12764 6009 12767
rect 5307 12736 6009 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 5997 12733 6009 12736
rect 6043 12764 6055 12767
rect 6187 12764 6215 12804
rect 6365 12801 6377 12804
rect 6411 12832 6423 12835
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6411 12804 6561 12832
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6043 12736 6215 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 6270 12724 6276 12776
rect 6328 12764 6334 12776
rect 6656 12764 6684 12872
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 14734 12900 14740 12912
rect 8904 12872 13952 12900
rect 8904 12860 8910 12872
rect 6822 12841 6828 12844
rect 6816 12795 6828 12841
rect 6880 12832 6886 12844
rect 6880 12804 6916 12832
rect 6822 12792 6828 12795
rect 6880 12792 6886 12804
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10606 12835 10664 12841
rect 10606 12832 10618 12835
rect 10192 12804 10618 12832
rect 10192 12792 10198 12804
rect 10606 12801 10618 12804
rect 10652 12801 10664 12835
rect 10606 12795 10664 12801
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11296 12804 11345 12832
rect 11296 12792 11302 12804
rect 11333 12801 11345 12804
rect 11379 12832 11391 12835
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11379 12804 11805 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 13354 12832 13360 12844
rect 11793 12795 11851 12801
rect 12406 12804 13360 12832
rect 7926 12764 7932 12776
rect 6328 12736 6684 12764
rect 7576 12736 7932 12764
rect 6328 12724 6334 12736
rect 5902 12656 5908 12708
rect 5960 12696 5966 12708
rect 6454 12696 6460 12708
rect 5960 12668 6460 12696
rect 5960 12656 5966 12668
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 4154 12628 4160 12640
rect 3467 12600 4160 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 7576 12628 7604 12736
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 10870 12764 10876 12776
rect 10831 12736 10876 12764
rect 10870 12724 10876 12736
rect 10928 12724 10934 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11204 12736 11621 12764
rect 11204 12724 11210 12736
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 12406 12696 12434 12804
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 13924 12773 13952 12872
rect 14660 12872 14740 12900
rect 14660 12841 14688 12872
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 15068 12804 15117 12832
rect 15068 12792 15074 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 13596 12736 13829 12764
rect 13596 12724 13602 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 14734 12764 14740 12776
rect 14695 12736 14740 12764
rect 13909 12727 13967 12733
rect 7708 12668 9628 12696
rect 7708 12656 7714 12668
rect 4948 12600 7604 12628
rect 7929 12631 7987 12637
rect 4948 12588 4954 12600
rect 7929 12597 7941 12631
rect 7975 12628 7987 12631
rect 8754 12628 8760 12640
rect 7975 12600 8760 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9490 12628 9496 12640
rect 9451 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9600 12628 9628 12668
rect 10888 12668 12434 12696
rect 13924 12696 13952 12727
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15286 12764 15292 12776
rect 14875 12736 15292 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 14844 12696 14872 12727
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 13924 12668 14872 12696
rect 10888 12628 10916 12668
rect 12250 12628 12256 12640
rect 9600 12600 10916 12628
rect 12211 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 15010 12628 15016 12640
rect 14056 12600 15016 12628
rect 14056 12588 14062 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 1394 12384 1400 12436
rect 1452 12424 1458 12436
rect 1489 12427 1547 12433
rect 1489 12424 1501 12427
rect 1452 12396 1501 12424
rect 1452 12384 1458 12396
rect 1489 12393 1501 12396
rect 1535 12393 1547 12427
rect 1489 12387 1547 12393
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 4246 12424 4252 12436
rect 3559 12396 4252 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 3528 12356 3556 12387
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 5684 12396 7389 12424
rect 5684 12384 5690 12396
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 10778 12424 10784 12436
rect 9447 12396 10784 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 12066 12384 12072 12436
rect 12124 12424 12130 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12124 12396 12541 12424
rect 12124 12384 12130 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 14090 12424 14096 12436
rect 13964 12396 14096 12424
rect 13964 12384 13970 12396
rect 14090 12384 14096 12396
rect 14148 12424 14154 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14148 12396 14381 12424
rect 14148 12384 14154 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14553 12427 14611 12433
rect 14553 12393 14565 12427
rect 14599 12424 14611 12427
rect 14826 12424 14832 12436
rect 14599 12396 14832 12424
rect 14599 12393 14611 12396
rect 14553 12387 14611 12393
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 14918 12384 14924 12436
rect 14976 12384 14982 12436
rect 3384 12328 3556 12356
rect 3384 12316 3390 12328
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 14182 12356 14188 12368
rect 11204 12328 14188 12356
rect 11204 12316 11210 12328
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2222 12288 2228 12300
rect 2179 12260 2228 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 9217 12291 9275 12297
rect 9217 12288 9229 12291
rect 8772 12260 9229 12288
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4890 12220 4896 12232
rect 4948 12229 4954 12232
rect 3752 12192 4896 12220
rect 3752 12180 3758 12192
rect 4890 12180 4896 12192
rect 4948 12220 4960 12229
rect 5184 12220 5212 12248
rect 5994 12220 6000 12232
rect 4948 12192 4993 12220
rect 5184 12192 6000 12220
rect 4948 12183 4960 12192
rect 4948 12180 4954 12183
rect 5994 12180 6000 12192
rect 6052 12220 6058 12232
rect 6546 12220 6552 12232
rect 6052 12192 6552 12220
rect 6052 12180 6058 12192
rect 6546 12180 6552 12192
rect 6604 12220 6610 12232
rect 8772 12229 8800 12260
rect 9217 12257 9229 12260
rect 9263 12288 9275 12291
rect 9306 12288 9312 12300
rect 9263 12260 9312 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 10870 12288 10876 12300
rect 10827 12260 10876 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11330 12248 11336 12300
rect 11388 12288 11394 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11388 12260 11897 12288
rect 11388 12248 11394 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 12308 12260 13277 12288
rect 12308 12248 12314 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13412 12260 13457 12288
rect 13412 12248 13418 12260
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 6604 12192 6653 12220
rect 6604 12180 6610 12192
rect 6641 12189 6653 12192
rect 6687 12220 6699 12223
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6687 12192 6745 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6733 12189 6745 12192
rect 6779 12220 6791 12223
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6779 12192 7205 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7193 12189 7205 12192
rect 7239 12220 7251 12223
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 7239 12192 8769 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 8757 12189 8769 12192
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 9398 12220 9404 12232
rect 8996 12192 9404 12220
rect 8996 12180 9002 12192
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 12986 12220 12992 12232
rect 11164 12192 12992 12220
rect 1857 12155 1915 12161
rect 1857 12121 1869 12155
rect 1903 12152 1915 12155
rect 4062 12152 4068 12164
rect 1903 12124 4068 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 6374 12155 6432 12161
rect 6374 12152 6386 12155
rect 5132 12124 6386 12152
rect 5132 12112 5138 12124
rect 6374 12121 6386 12124
rect 6420 12121 6432 12155
rect 6374 12115 6432 12121
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 8110 12152 8116 12164
rect 6972 12124 8116 12152
rect 6972 12112 6978 12124
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 8512 12155 8570 12161
rect 8512 12121 8524 12155
rect 8558 12152 8570 12155
rect 9030 12152 9036 12164
rect 8558 12124 9036 12152
rect 8558 12121 8570 12124
rect 8512 12115 8570 12121
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 10514 12155 10572 12161
rect 10514 12152 10526 12155
rect 10008 12124 10526 12152
rect 10008 12112 10014 12124
rect 10514 12121 10526 12124
rect 10560 12152 10572 12155
rect 11164 12152 11192 12192
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14936 12220 14964 12384
rect 15194 12288 15200 12300
rect 15155 12260 15200 12288
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 13964 12192 14964 12220
rect 13964 12180 13970 12192
rect 10560 12124 11192 12152
rect 10560 12121 10572 12124
rect 10514 12115 10572 12121
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 11848 12124 12173 12152
rect 11848 12112 11854 12124
rect 12161 12121 12173 12124
rect 12207 12121 12219 12155
rect 12161 12115 12219 12121
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 12308 12124 12725 12152
rect 12308 12112 12314 12124
rect 12713 12121 12725 12124
rect 12759 12152 12771 12155
rect 13173 12155 13231 12161
rect 13173 12152 13185 12155
rect 12759 12124 13185 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 13173 12121 13185 12124
rect 13219 12121 13231 12155
rect 13173 12115 13231 12121
rect 14090 12112 14096 12164
rect 14148 12152 14154 12164
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 14148 12124 15025 12152
rect 14148 12112 14154 12124
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2004 12056 2049 12084
rect 2004 12044 2010 12056
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3660 12056 3801 12084
rect 3660 12044 3666 12056
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 5258 12084 5264 12096
rect 5219 12056 5264 12084
rect 3789 12047 3847 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 9674 12084 9680 12096
rect 6512 12056 9680 12084
rect 6512 12044 6518 12056
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 12066 12084 12072 12096
rect 12027 12056 12072 12084
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 12986 12084 12992 12096
rect 12851 12056 12992 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 13688 12056 14289 12084
rect 13688 12044 13694 12056
rect 14277 12053 14289 12056
rect 14323 12084 14335 12087
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14323 12056 14933 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 1946 11880 1952 11892
rect 1627 11852 1952 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 1946 11840 1952 11852
rect 2004 11840 2010 11892
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 2130 11880 2136 11892
rect 2087 11852 2136 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 7466 11880 7472 11892
rect 2280 11852 7472 11880
rect 2280 11840 2286 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7616 11852 12020 11880
rect 7616 11840 7622 11852
rect 4246 11772 4252 11824
rect 4304 11772 4310 11824
rect 4430 11772 4436 11824
rect 4488 11812 4494 11824
rect 5046 11815 5104 11821
rect 5046 11812 5058 11815
rect 4488 11784 5058 11812
rect 4488 11772 4494 11784
rect 5046 11781 5058 11784
rect 5092 11812 5104 11815
rect 5442 11812 5448 11824
rect 5092 11784 5448 11812
rect 5092 11781 5104 11784
rect 5046 11775 5104 11781
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 6457 11815 6515 11821
rect 6457 11781 6469 11815
rect 6503 11812 6515 11815
rect 6546 11812 6552 11824
rect 6503 11784 6552 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 6546 11772 6552 11784
rect 6604 11812 6610 11824
rect 6604 11784 8156 11812
rect 6604 11772 6610 11784
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2314 11744 2320 11756
rect 1995 11716 2320 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3585 11747 3643 11753
rect 3585 11744 3597 11747
rect 3436 11716 3597 11744
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2271 11648 2544 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2516 11549 2544 11648
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3436 11676 3464 11716
rect 3585 11713 3597 11716
rect 3631 11713 3643 11747
rect 4264 11744 4292 11772
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4264 11716 4813 11744
rect 3585 11707 3643 11713
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 7558 11744 7564 11756
rect 4948 11716 7564 11744
rect 4948 11704 4954 11716
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8128 11753 8156 11784
rect 10226 11772 10232 11824
rect 10284 11812 10290 11824
rect 10962 11812 10968 11824
rect 10284 11784 10968 11812
rect 10284 11772 10290 11784
rect 10962 11772 10968 11784
rect 11020 11772 11026 11824
rect 11057 11815 11115 11821
rect 11057 11781 11069 11815
rect 11103 11812 11115 11815
rect 11793 11815 11851 11821
rect 11793 11812 11805 11815
rect 11103 11784 11805 11812
rect 11103 11781 11115 11784
rect 11057 11775 11115 11781
rect 11793 11781 11805 11784
rect 11839 11781 11851 11815
rect 11793 11775 11851 11781
rect 7857 11747 7915 11753
rect 7857 11713 7869 11747
rect 7903 11744 7915 11747
rect 8113 11747 8171 11753
rect 7903 11716 8064 11744
rect 7903 11713 7915 11716
rect 7857 11707 7915 11713
rect 2648 11648 3464 11676
rect 8036 11676 8064 11716
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 11072 11744 11100 11775
rect 8536 11716 11100 11744
rect 8536 11704 8542 11716
rect 11146 11704 11152 11756
rect 11204 11744 11210 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 11204 11716 11253 11744
rect 11204 11704 11210 11716
rect 11241 11713 11253 11716
rect 11287 11744 11299 11747
rect 11514 11744 11520 11756
rect 11287 11716 11520 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 11514 11704 11520 11716
rect 11572 11744 11578 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11572 11716 11897 11744
rect 11572 11704 11578 11716
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 9490 11676 9496 11688
rect 8036 11648 9496 11676
rect 2648 11636 2654 11648
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 11606 11676 11612 11688
rect 9732 11648 11612 11676
rect 9732 11636 9738 11648
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 11992 11676 12020 11852
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 12124 11852 12265 11880
rect 12124 11840 12130 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 13170 11840 13176 11892
rect 13228 11880 13234 11892
rect 13630 11880 13636 11892
rect 13228 11852 13636 11880
rect 13228 11840 13234 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 13541 11815 13599 11821
rect 13541 11781 13553 11815
rect 13587 11812 13599 11815
rect 13814 11812 13820 11824
rect 13587 11784 13820 11812
rect 13587 11781 13599 11784
rect 13541 11775 13599 11781
rect 13814 11772 13820 11784
rect 13872 11812 13878 11824
rect 13872 11784 14136 11812
rect 13872 11772 13878 11784
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13630 11744 13636 11756
rect 13403 11716 13636 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 13998 11744 14004 11756
rect 13959 11716 14004 11744
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14108 11753 14136 11784
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14550 11744 14556 11756
rect 14139 11716 14556 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 11992 11648 13952 11676
rect 6104 11580 7236 11608
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 4706 11540 4712 11552
rect 2547 11512 4712 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 6104 11540 6132 11580
rect 5500 11512 6132 11540
rect 5500 11500 5506 11512
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 6236 11512 6281 11540
rect 6236 11500 6242 11512
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6733 11543 6791 11549
rect 6733 11540 6745 11543
rect 6512 11512 6745 11540
rect 6512 11500 6518 11512
rect 6733 11509 6745 11512
rect 6779 11509 6791 11543
rect 7208 11540 7236 11580
rect 8110 11568 8116 11620
rect 8168 11608 8174 11620
rect 11514 11608 11520 11620
rect 8168 11580 11520 11608
rect 8168 11568 8174 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 13924 11608 13952 11648
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14458 11676 14464 11688
rect 14240 11648 14464 11676
rect 14240 11636 14246 11648
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 15194 11608 15200 11620
rect 13924 11580 15200 11608
rect 15194 11568 15200 11580
rect 15252 11568 15258 11620
rect 11422 11540 11428 11552
rect 7208 11512 11428 11540
rect 6733 11503 6791 11509
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2498 11336 2504 11348
rect 2372 11308 2504 11336
rect 2372 11296 2378 11308
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 4522 11336 4528 11348
rect 4479 11308 4528 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 4522 11296 4528 11308
rect 4580 11336 4586 11348
rect 4890 11336 4896 11348
rect 4580 11308 4896 11336
rect 4580 11296 4586 11308
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5994 11336 6000 11348
rect 5955 11308 6000 11336
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 8260 11308 9505 11336
rect 8260 11296 8266 11308
rect 9493 11305 9505 11308
rect 9539 11336 9551 11339
rect 10134 11336 10140 11348
rect 9539 11308 10140 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11112 11308 11437 11336
rect 11112 11296 11118 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11425 11299 11483 11305
rect 6012 11268 6040 11296
rect 5828 11240 6040 11268
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 3694 11200 3700 11212
rect 2363 11172 3700 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 5828 11209 5856 11240
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 8478 11268 8484 11280
rect 7800 11240 8484 11268
rect 7800 11228 7806 11240
rect 8220 11212 8248 11240
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6454 11200 6460 11212
rect 6328 11172 6460 11200
rect 6328 11160 6334 11172
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 8202 11160 8208 11212
rect 8260 11160 8266 11212
rect 10870 11200 10876 11212
rect 10831 11172 10876 11200
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2087 11104 2912 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 1946 11024 1952 11076
rect 2004 11064 2010 11076
rect 2685 11067 2743 11073
rect 2685 11064 2697 11067
rect 2004 11036 2697 11064
rect 2004 11024 2010 11036
rect 2685 11033 2697 11036
rect 2731 11033 2743 11067
rect 2884 11064 2912 11104
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3016 11104 3061 11132
rect 3016 11092 3022 11104
rect 5534 11092 5540 11144
rect 5592 11141 5598 11144
rect 5592 11132 5604 11141
rect 10617 11135 10675 11141
rect 5592 11104 5637 11132
rect 8404 11104 10548 11132
rect 5592 11095 5604 11104
rect 5592 11092 5598 11095
rect 5442 11064 5448 11076
rect 2884 11036 5448 11064
rect 2685 11027 2743 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 8404 11064 8432 11104
rect 5736 11036 8432 11064
rect 9401 11067 9459 11073
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1673 10999 1731 11005
rect 1673 10996 1685 10999
rect 1544 10968 1685 10996
rect 1544 10956 1550 10968
rect 1673 10965 1685 10968
rect 1719 10965 1731 10999
rect 1673 10959 1731 10965
rect 2133 10999 2191 11005
rect 2133 10965 2145 10999
rect 2179 10996 2191 10999
rect 5736 10996 5764 11036
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9674 11064 9680 11076
rect 9447 11036 9680 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10520 11064 10548 11104
rect 10617 11101 10629 11135
rect 10663 11132 10675 11135
rect 10778 11132 10784 11144
rect 10663 11104 10784 11132
rect 10663 11101 10675 11104
rect 10617 11095 10675 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11440 11132 11468 11299
rect 11514 11296 11520 11348
rect 11572 11296 11578 11348
rect 11790 11336 11796 11348
rect 11751 11308 11796 11336
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13136 11308 13553 11336
rect 13136 11296 13142 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 13541 11299 13599 11305
rect 11532 11268 11560 11296
rect 13556 11268 13584 11299
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 13780 11308 14657 11336
rect 13780 11296 13786 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 14645 11299 14703 11305
rect 14090 11268 14096 11280
rect 11532 11240 13308 11268
rect 13556 11240 14096 11268
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 13280 11209 13308 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14366 11268 14372 11280
rect 14327 11240 14372 11268
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 11664 11172 12357 11200
rect 11664 11160 11670 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11169 13323 11203
rect 15194 11200 15200 11212
rect 15155 11172 15200 11200
rect 13265 11163 13323 11169
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 11440 11104 12173 11132
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12161 11095 12219 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13280 11132 13308 11163
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15286 11132 15292 11144
rect 13280 11104 15292 11132
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 11422 11064 11428 11076
rect 10520 11036 11428 11064
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11701 11067 11759 11073
rect 11701 11033 11713 11067
rect 11747 11064 11759 11067
rect 12066 11064 12072 11076
rect 11747 11036 12072 11064
rect 11747 11033 11759 11036
rect 11701 11027 11759 11033
rect 12066 11024 12072 11036
rect 12124 11064 12130 11076
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 12124 11036 12265 11064
rect 12124 11024 12130 11036
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14240 11036 15025 11064
rect 14240 11024 14246 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15013 11027 15071 11033
rect 2179 10968 5764 10996
rect 2179 10965 2191 10968
rect 2133 10959 2191 10965
rect 5810 10956 5816 11008
rect 5868 10996 5874 11008
rect 6454 10996 6460 11008
rect 5868 10968 6460 10996
rect 5868 10956 5874 10968
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 11238 10996 11244 11008
rect 6696 10968 11244 10996
rect 6696 10956 6702 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12618 10996 12624 11008
rect 12579 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 13817 10999 13875 11005
rect 13136 10968 13181 10996
rect 13136 10956 13142 10968
rect 13817 10965 13829 10999
rect 13863 10996 13875 10999
rect 14366 10996 14372 11008
rect 13863 10968 14372 10996
rect 13863 10965 13875 10968
rect 13817 10959 13875 10965
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 15105 10999 15163 11005
rect 15105 10996 15117 10999
rect 14608 10968 15117 10996
rect 14608 10956 14614 10968
rect 15105 10965 15117 10968
rect 15151 10996 15163 10999
rect 15654 10996 15660 11008
rect 15151 10968 15660 10996
rect 15151 10965 15163 10968
rect 15105 10959 15163 10965
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 2682 10792 2688 10804
rect 2280 10764 2688 10792
rect 2280 10752 2286 10764
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4246 10792 4252 10804
rect 4111 10764 4252 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 1486 10656 1492 10668
rect 1447 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 3602 10616 3608 10668
rect 3660 10665 3666 10668
rect 3660 10656 3672 10665
rect 3878 10656 3884 10668
rect 3660 10628 3705 10656
rect 3791 10628 3884 10656
rect 3660 10619 3672 10628
rect 3660 10616 3666 10619
rect 3878 10616 3884 10628
rect 3936 10656 3942 10668
rect 4080 10656 4108 10755
rect 4246 10752 4252 10764
rect 4304 10792 4310 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4304 10764 4813 10792
rect 4304 10752 4310 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6052 10764 6377 10792
rect 6052 10752 6058 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 6178 10724 6184 10736
rect 5592 10696 6184 10724
rect 5592 10684 5598 10696
rect 6178 10684 6184 10696
rect 6236 10684 6242 10736
rect 6380 10724 6408 10755
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6512 10764 8984 10792
rect 6512 10752 6518 10764
rect 8288 10727 8346 10733
rect 6380 10696 8064 10724
rect 3936 10628 4108 10656
rect 6380 10656 6408 10696
rect 8036 10665 8064 10696
rect 8288 10693 8300 10727
rect 8334 10724 8346 10727
rect 8846 10724 8852 10736
rect 8334 10696 8852 10724
rect 8334 10693 8346 10696
rect 8288 10687 8346 10693
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 8956 10724 8984 10764
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10962 10792 10968 10804
rect 10284 10764 10968 10792
rect 10284 10752 10290 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12342 10792 12348 10804
rect 12032 10764 12348 10792
rect 12032 10752 12038 10764
rect 12342 10752 12348 10764
rect 12400 10792 12406 10804
rect 12713 10795 12771 10801
rect 12713 10792 12725 10795
rect 12400 10764 12725 10792
rect 12400 10752 12406 10764
rect 12713 10761 12725 10764
rect 12759 10761 12771 10795
rect 13078 10792 13084 10804
rect 13039 10764 13084 10792
rect 12713 10755 12771 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13587 10764 13921 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 14090 10792 14096 10804
rect 13909 10755 13967 10761
rect 14016 10764 14096 10792
rect 13449 10727 13507 10733
rect 8956 10696 12434 10724
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6380 10628 6561 10656
rect 3936 10616 3942 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6816 10659 6874 10665
rect 6816 10625 6828 10659
rect 6862 10656 6874 10659
rect 8021 10659 8079 10665
rect 6862 10628 7972 10656
rect 6862 10625 6874 10628
rect 6816 10619 6874 10625
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1452 10560 1685 10588
rect 1452 10548 1458 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 7944 10588 7972 10628
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8754 10656 8760 10668
rect 8021 10619 8079 10625
rect 8128 10628 8760 10656
rect 8128 10588 8156 10628
rect 8754 10616 8760 10628
rect 8812 10656 8818 10668
rect 9398 10656 9404 10668
rect 8812 10628 9404 10656
rect 8812 10616 8818 10628
rect 9398 10616 9404 10628
rect 9456 10616 9462 10668
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10606 10659 10664 10665
rect 10606 10656 10618 10659
rect 10284 10628 10618 10656
rect 10284 10616 10290 10628
rect 10606 10625 10618 10628
rect 10652 10625 10664 10659
rect 10870 10656 10876 10668
rect 10831 10628 10876 10656
rect 10606 10619 10664 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 12406 10588 12434 10696
rect 13449 10693 13461 10727
rect 13495 10724 13507 10727
rect 13630 10724 13636 10736
rect 13495 10696 13636 10724
rect 13495 10693 13507 10696
rect 13449 10687 13507 10693
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14016 10724 14044 10764
rect 14090 10752 14096 10764
rect 14148 10792 14154 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 14148 10764 14289 10792
rect 14148 10752 14154 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 14366 10752 14372 10804
rect 14424 10792 14430 10804
rect 15746 10792 15752 10804
rect 14424 10764 15752 10792
rect 14424 10752 14430 10764
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 13872 10696 14044 10724
rect 13872 10684 13878 10696
rect 14550 10684 14556 10736
rect 14608 10724 14614 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 14608 10696 15209 10724
rect 14608 10684 14614 10696
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15197 10687 15255 10693
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14700 10628 15117 10656
rect 14700 10616 14706 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 13354 10588 13360 10600
rect 7944 10560 8156 10588
rect 9048 10560 9904 10588
rect 12406 10560 13360 10588
rect 1673 10551 1731 10557
rect 2498 10452 2504 10464
rect 2459 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10412 2562 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7926 10452 7932 10464
rect 7708 10424 7932 10452
rect 7708 10412 7714 10424
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9048 10452 9076 10560
rect 9401 10523 9459 10529
rect 9401 10489 9413 10523
rect 9447 10520 9459 10523
rect 9766 10520 9772 10532
rect 9447 10492 9772 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 9490 10452 9496 10464
rect 8352 10424 9076 10452
rect 9451 10424 9496 10452
rect 8352 10412 8358 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9876 10452 9904 10560
rect 13354 10548 13360 10560
rect 13412 10588 13418 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13412 10560 13645 10588
rect 13412 10548 13418 10560
rect 13633 10557 13645 10560
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 15289 10591 15347 10597
rect 14516 10560 14561 10588
rect 14516 10548 14522 10560
rect 15289 10557 15301 10591
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 15304 10520 15332 10551
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 12406 10492 15577 10520
rect 12406 10452 12434 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 15565 10483 15623 10489
rect 14734 10452 14740 10464
rect 9876 10424 12434 10452
rect 14695 10424 14740 10452
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 3878 10248 3884 10260
rect 3839 10220 3884 10248
rect 3878 10208 3884 10220
rect 3936 10248 3942 10260
rect 4246 10248 4252 10260
rect 3936 10220 4252 10248
rect 3936 10208 3942 10220
rect 4246 10208 4252 10220
rect 4304 10248 4310 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4304 10220 4353 10248
rect 4304 10208 4310 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 7285 10251 7343 10257
rect 4341 10211 4399 10217
rect 5920 10220 6960 10248
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 3896 10112 3924 10208
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 5920 10180 5948 10220
rect 4120 10152 5948 10180
rect 4120 10140 4126 10152
rect 3651 10084 3924 10112
rect 5905 10115 5963 10121
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 3360 9979 3418 9985
rect 3360 9945 3372 9979
rect 3406 9976 3418 9979
rect 5258 9976 5264 9988
rect 3406 9948 5264 9976
rect 3406 9945 3418 9948
rect 3360 9939 3418 9945
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5813 9979 5871 9985
rect 5813 9945 5825 9979
rect 5859 9976 5871 9979
rect 5920 9976 5948 10075
rect 6932 10044 6960 10220
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 8110 10248 8116 10260
rect 7331 10220 8116 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9272 10220 9505 10248
rect 9272 10208 9278 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 11422 10248 11428 10260
rect 9493 10211 9551 10217
rect 9600 10220 10916 10248
rect 11383 10220 11428 10248
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 9600 10180 9628 10220
rect 7708 10152 9628 10180
rect 10888 10180 10916 10220
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 11664 10220 12265 10248
rect 11664 10208 11670 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12253 10211 12311 10217
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 13817 10251 13875 10257
rect 12400 10220 13400 10248
rect 12400 10208 12406 10220
rect 12360 10180 12388 10208
rect 10888 10152 12388 10180
rect 7708 10140 7714 10152
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7374 10112 7380 10124
rect 7156 10084 7380 10112
rect 7156 10072 7162 10084
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 10870 10112 10876 10124
rect 10831 10084 10876 10112
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11977 10115 12035 10121
rect 11977 10112 11989 10115
rect 11020 10084 11989 10112
rect 11020 10072 11026 10084
rect 11977 10081 11989 10084
rect 12023 10112 12035 10115
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12023 10084 12817 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12805 10081 12817 10084
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13372 10121 13400 10220
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 14550 10248 14556 10260
rect 13863 10220 14556 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 14200 10152 15240 10180
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12952 10084 13185 10112
rect 12952 10072 12958 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14200 10121 14228 10152
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13872 10084 14197 10112
rect 13872 10072 13878 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14458 10112 14464 10124
rect 14419 10084 14464 10112
rect 14185 10075 14243 10081
rect 14458 10072 14464 10084
rect 14516 10112 14522 10124
rect 15102 10112 15108 10124
rect 14516 10084 14872 10112
rect 15063 10084 15108 10112
rect 14516 10072 14522 10084
rect 14734 10044 14740 10056
rect 6932 10016 14740 10044
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 14844 10044 14872 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14844 10016 15025 10044
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 5994 9976 6000 9988
rect 5859 9948 6000 9976
rect 5859 9945 5871 9948
rect 5813 9939 5871 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 6172 9979 6230 9985
rect 6172 9945 6184 9979
rect 6218 9976 6230 9979
rect 6454 9976 6460 9988
rect 6218 9948 6460 9976
rect 6218 9945 6230 9948
rect 6172 9939 6230 9945
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9272 9948 10088 9976
rect 9272 9936 9278 9948
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 2590 9908 2596 9920
rect 2271 9880 2596 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 2590 9868 2596 9880
rect 2648 9908 2654 9920
rect 7190 9908 7196 9920
rect 2648 9880 7196 9908
rect 2648 9868 2654 9880
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9908 7898 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 7892 9880 9137 9908
rect 7892 9868 7898 9880
rect 9125 9877 9137 9880
rect 9171 9908 9183 9911
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9171 9880 9321 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9309 9877 9321 9880
rect 9355 9908 9367 9911
rect 9674 9908 9680 9920
rect 9355 9880 9680 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 10060 9908 10088 9948
rect 10134 9936 10140 9988
rect 10192 9976 10198 9988
rect 10606 9979 10664 9985
rect 10606 9976 10618 9979
rect 10192 9948 10618 9976
rect 10192 9936 10198 9948
rect 10606 9945 10618 9948
rect 10652 9945 10664 9979
rect 10606 9939 10664 9945
rect 12621 9979 12679 9985
rect 12621 9945 12633 9979
rect 12667 9976 12679 9979
rect 13170 9976 13176 9988
rect 12667 9948 13176 9976
rect 12667 9945 12679 9948
rect 12621 9939 12679 9945
rect 13170 9936 13176 9948
rect 13228 9936 13234 9988
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 14921 9979 14979 9985
rect 13596 9948 14596 9976
rect 13596 9936 13602 9948
rect 10502 9908 10508 9920
rect 10060 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 11790 9908 11796 9920
rect 11751 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 11940 9880 11985 9908
rect 11940 9868 11946 9880
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12768 9880 12813 9908
rect 12768 9868 12774 9880
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 14568 9917 14596 9948
rect 14921 9945 14933 9979
rect 14967 9976 14979 9979
rect 15212 9976 15240 10152
rect 15746 9976 15752 9988
rect 14967 9948 15752 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13044 9880 13461 9908
rect 13044 9868 13050 9880
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 14553 9911 14611 9917
rect 14553 9877 14565 9911
rect 14599 9877 14611 9911
rect 14553 9871 14611 9877
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 2869 9707 2927 9713
rect 2869 9673 2881 9707
rect 2915 9673 2927 9707
rect 2869 9667 2927 9673
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2774 9636 2780 9648
rect 2547 9608 2780 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2884 9636 2912 9667
rect 5166 9664 5172 9716
rect 5224 9704 5230 9716
rect 6638 9704 6644 9716
rect 5224 9676 6644 9704
rect 5224 9664 5230 9676
rect 3326 9636 3332 9648
rect 2884 9608 3332 9636
rect 3326 9596 3332 9608
rect 3384 9636 3390 9648
rect 6012 9645 6040 9676
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 9585 9707 9643 9713
rect 7248 9676 9536 9704
rect 7248 9664 7254 9676
rect 5997 9639 6055 9645
rect 3384 9608 5600 9636
rect 3384 9596 3390 9608
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 2148 9540 2237 9568
rect 1489 9503 1547 9509
rect 1489 9469 1501 9503
rect 1535 9469 1547 9503
rect 1670 9500 1676 9512
rect 1631 9472 1676 9500
rect 1489 9463 1547 9469
rect 1504 9364 1532 9463
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2148 9441 2176 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2590 9528 2596 9580
rect 2648 9568 2654 9580
rect 3993 9571 4051 9577
rect 3993 9568 4005 9571
rect 2648 9540 4005 9568
rect 2648 9528 2654 9540
rect 3993 9537 4005 9540
rect 4039 9568 4051 9571
rect 4614 9568 4620 9580
rect 4039 9540 4620 9568
rect 4039 9537 4051 9540
rect 3993 9531 4051 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 5572 9577 5600 9608
rect 5997 9605 6009 9639
rect 6043 9605 6055 9639
rect 7466 9636 7472 9648
rect 5997 9599 6055 9605
rect 6084 9608 7472 9636
rect 5557 9571 5615 9577
rect 5557 9537 5569 9571
rect 5603 9568 5615 9571
rect 6084 9568 6112 9608
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 9508 9636 9536 9676
rect 9585 9673 9597 9707
rect 9631 9704 9643 9707
rect 9674 9704 9680 9716
rect 9631 9676 9680 9704
rect 9631 9673 9643 9676
rect 9585 9667 9643 9673
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 12710 9704 12716 9716
rect 9784 9676 12434 9704
rect 12671 9676 12716 9704
rect 9784 9636 9812 9676
rect 9508 9608 9812 9636
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 10790 9639 10848 9645
rect 10790 9636 10802 9639
rect 10560 9608 10802 9636
rect 10560 9596 10566 9608
rect 10790 9605 10802 9608
rect 10836 9605 10848 9639
rect 12406 9636 12434 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 12986 9704 12992 9716
rect 12947 9676 12992 9704
rect 12986 9664 12992 9676
rect 13044 9664 13050 9716
rect 13170 9704 13176 9716
rect 13131 9676 13176 9704
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 12894 9636 12900 9648
rect 12406 9608 12900 9636
rect 10790 9599 10848 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 13354 9596 13360 9648
rect 13412 9636 13418 9648
rect 15105 9639 15163 9645
rect 13412 9608 15056 9636
rect 13412 9596 13418 9608
rect 6638 9577 6644 9580
rect 6632 9568 6644 9577
rect 5603 9540 6112 9568
rect 6599 9540 6644 9568
rect 5603 9537 5615 9540
rect 5557 9531 5615 9537
rect 6632 9531 6644 9540
rect 6638 9528 6644 9531
rect 6696 9528 6702 9580
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8021 9571 8079 9577
rect 8021 9568 8033 9571
rect 7892 9540 8033 9568
rect 7892 9528 7898 9540
rect 8021 9537 8033 9540
rect 8067 9537 8079 9571
rect 8288 9571 8346 9577
rect 8288 9568 8300 9571
rect 8021 9531 8079 9537
rect 8128 9540 8300 9568
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 5813 9503 5871 9509
rect 5813 9469 5825 9503
rect 5859 9500 5871 9503
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 5859 9472 6377 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 8128 9500 8156 9540
rect 8288 9537 8300 9540
rect 8334 9568 8346 9571
rect 12345 9571 12403 9577
rect 8334 9540 9251 9568
rect 8334 9537 8346 9540
rect 8288 9531 8346 9537
rect 6365 9463 6423 9469
rect 7760 9472 8156 9500
rect 9223 9500 9251 9540
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 13446 9568 13452 9580
rect 12391 9540 13452 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 14001 9571 14059 9577
rect 14001 9568 14013 9571
rect 13587 9540 14013 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 14001 9537 14013 9540
rect 14047 9537 14059 9571
rect 15028 9568 15056 9608
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 15194 9636 15200 9648
rect 15151 9608 15200 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 15028 9540 15332 9568
rect 14001 9531 14059 9537
rect 11054 9500 11060 9512
rect 9223 9472 9812 9500
rect 11015 9472 11060 9500
rect 2133 9435 2191 9441
rect 2133 9401 2145 9435
rect 2179 9401 2191 9435
rect 2133 9395 2191 9401
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 1504 9336 4445 9364
rect 4433 9333 4445 9336
rect 4479 9364 4491 9367
rect 5074 9364 5080 9376
rect 4479 9336 5080 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5828 9364 5856 9463
rect 7760 9441 7788 9472
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9401 7803 9435
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 7745 9395 7803 9401
rect 9600 9404 9689 9432
rect 9600 9376 9628 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 9677 9395 9735 9401
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5500 9336 6101 9364
rect 5500 9324 5506 9336
rect 6089 9333 6101 9336
rect 6135 9364 6147 9367
rect 7834 9364 7840 9376
rect 6135 9336 7840 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 7834 9324 7840 9336
rect 7892 9364 7898 9376
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 7892 9336 7941 9364
rect 7892 9324 7898 9336
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 7929 9327 7987 9333
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9364 9336 9413 9364
rect 9364 9324 9370 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 9582 9324 9588 9376
rect 9640 9324 9646 9376
rect 9784 9364 9812 9472
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 12161 9503 12219 9509
rect 12161 9469 12173 9503
rect 12207 9469 12219 9503
rect 12161 9463 12219 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12526 9500 12532 9512
rect 12299 9472 12532 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12176 9432 12204 9463
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 13630 9500 13636 9512
rect 13591 9472 13636 9500
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 15304 9509 15332 9540
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9469 15347 9503
rect 15289 9463 15347 9469
rect 12710 9432 12716 9444
rect 11756 9404 12716 9432
rect 11756 9392 11762 9404
rect 12710 9392 12716 9404
rect 12768 9432 12774 9444
rect 13740 9432 13768 9463
rect 12768 9404 13768 9432
rect 12768 9392 12774 9404
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 15010 9432 15016 9444
rect 13872 9404 15016 9432
rect 13872 9392 13878 9404
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 12066 9364 12072 9376
rect 9784 9336 12072 9364
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 13688 9336 14289 9364
rect 13688 9324 13694 9336
rect 14277 9333 14289 9336
rect 14323 9364 14335 9367
rect 14458 9364 14464 9376
rect 14323 9336 14464 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14608 9336 14749 9364
rect 14608 9324 14614 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 15212 9364 15240 9463
rect 15378 9364 15384 9376
rect 15212 9336 15384 9364
rect 14737 9327 14795 9333
rect 15378 9324 15384 9336
rect 15436 9364 15442 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15436 9336 15577 9364
rect 15436 9324 15442 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 6052 9132 8585 9160
rect 6052 9120 6058 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 5353 9095 5411 9101
rect 5353 9061 5365 9095
rect 5399 9092 5411 9095
rect 5626 9092 5632 9104
rect 5399 9064 5632 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 7098 9092 7104 9104
rect 7059 9064 7104 9092
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 8588 9092 8616 9123
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 8904 9132 9413 9160
rect 8904 9120 8910 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 13173 9163 13231 9169
rect 9401 9123 9459 9129
rect 9876 9132 12434 9160
rect 9876 9092 9904 9132
rect 8588 9064 9904 9092
rect 10962 9052 10968 9104
rect 11020 9092 11026 9104
rect 12406 9092 12434 9132
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 14642 9160 14648 9172
rect 13219 9132 14648 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15286 9160 15292 9172
rect 14844 9132 15292 9160
rect 13357 9095 13415 9101
rect 11020 9064 12296 9092
rect 12406 9064 13308 9092
rect 11020 9052 11026 9064
rect 3878 8984 3884 9036
rect 3936 9024 3942 9036
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3936 8996 3985 9024
rect 3936 8984 3942 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5500 8996 5733 9024
rect 5500 8984 5506 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9582 9024 9588 9036
rect 9088 8996 9588 9024
rect 9088 8984 9094 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 11974 9024 11980 9036
rect 11164 8996 11980 9024
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2188 8928 2237 8956
rect 2188 8916 2194 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 3620 8928 5672 8956
rect 2492 8891 2550 8897
rect 2492 8857 2504 8891
rect 2538 8888 2550 8891
rect 2682 8888 2688 8900
rect 2538 8860 2688 8888
rect 2538 8857 2550 8860
rect 2492 8851 2550 8857
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 3620 8829 3648 8928
rect 4218 8891 4276 8897
rect 4218 8888 4230 8891
rect 3804 8860 4230 8888
rect 3804 8832 3832 8860
rect 4218 8857 4230 8860
rect 4264 8857 4276 8891
rect 4218 8851 4276 8857
rect 5442 8848 5448 8900
rect 5500 8888 5506 8900
rect 5537 8891 5595 8897
rect 5537 8888 5549 8891
rect 5500 8860 5549 8888
rect 5500 8848 5506 8860
rect 5537 8857 5549 8860
rect 5583 8857 5595 8891
rect 5644 8888 5672 8928
rect 6730 8916 6736 8968
rect 6788 8956 6794 8968
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 6788 8928 7205 8956
rect 6788 8916 6794 8928
rect 7193 8925 7205 8928
rect 7239 8956 7251 8959
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 7239 8928 8677 8956
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 8665 8925 8677 8928
rect 8711 8956 8723 8959
rect 8846 8956 8852 8968
rect 8711 8928 8852 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 8846 8916 8852 8928
rect 8904 8956 8910 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8904 8928 9229 8956
rect 8904 8916 8910 8928
rect 9217 8925 9229 8928
rect 9263 8956 9275 8959
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 9263 8928 10793 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 10781 8925 10793 8928
rect 10827 8956 10839 8959
rect 11054 8956 11060 8968
rect 10827 8928 11060 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 5810 8888 5816 8900
rect 5644 8860 5816 8888
rect 5537 8851 5595 8857
rect 5810 8848 5816 8860
rect 5868 8888 5874 8900
rect 5966 8891 6024 8897
rect 5966 8888 5978 8891
rect 5868 8860 5978 8888
rect 5868 8848 5874 8860
rect 5966 8857 5978 8860
rect 6012 8857 6024 8891
rect 5966 8851 6024 8857
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 7438 8891 7496 8897
rect 7438 8888 7450 8891
rect 6236 8860 7450 8888
rect 6236 8848 6242 8860
rect 7438 8857 7450 8860
rect 7484 8857 7496 8891
rect 7438 8851 7496 8857
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 10514 8891 10572 8897
rect 10514 8888 10526 8891
rect 9824 8860 10526 8888
rect 9824 8848 9830 8860
rect 10514 8857 10526 8860
rect 10560 8857 10572 8891
rect 10514 8851 10572 8857
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8789 3663 8823
rect 3786 8820 3792 8832
rect 3747 8792 3792 8820
rect 3605 8783 3663 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 11164 8820 11192 8996
rect 11974 8984 11980 8996
rect 12032 9024 12038 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 12032 8996 12173 9024
rect 12032 8984 12038 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11296 8928 12081 8956
rect 11296 8916 11302 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11563 8860 11989 8888
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 12268 8888 12296 9064
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 12894 9024 12900 9036
rect 12667 8996 12900 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13280 9024 13308 9064
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 13446 9092 13452 9104
rect 13403 9064 13452 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13722 9092 13728 9104
rect 13683 9064 13728 9092
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 14844 9033 14872 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 15160 9064 15332 9092
rect 15160 9052 15166 9064
rect 15304 9033 15332 9064
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 16390 9092 16396 9104
rect 15528 9064 16396 9092
rect 15528 9052 15534 9064
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 14829 9027 14887 9033
rect 13280 8996 14780 9024
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 12584 8928 13461 8956
rect 12584 8916 12590 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 14550 8956 14556 8968
rect 14511 8928 14556 8956
rect 13449 8919 13507 8925
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14752 8956 14780 8996
rect 14829 8993 14841 9027
rect 14875 8993 14887 9027
rect 15289 9027 15347 9033
rect 14829 8987 14887 8993
rect 15028 8996 15240 9024
rect 15028 8956 15056 8996
rect 14752 8928 15056 8956
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8925 15163 8959
rect 15212 8956 15240 8996
rect 15289 8993 15301 9027
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15470 8956 15476 8968
rect 15212 8928 15476 8956
rect 15105 8919 15163 8925
rect 12713 8891 12771 8897
rect 12713 8888 12725 8891
rect 12268 8860 12725 8888
rect 11977 8851 12035 8857
rect 12713 8857 12725 8860
rect 12759 8888 12771 8891
rect 13722 8888 13728 8900
rect 12759 8860 13728 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 15120 8888 15148 8919
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15286 8888 15292 8900
rect 15120 8860 15292 8888
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 4672 8792 11192 8820
rect 4672 8780 4678 8792
rect 11422 8780 11428 8832
rect 11480 8820 11486 8832
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11480 8792 11621 8820
rect 11480 8780 11486 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 12860 8792 12905 8820
rect 12860 8780 12866 8792
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13630 8820 13636 8832
rect 13136 8792 13636 8820
rect 13136 8780 13142 8792
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14185 8823 14243 8829
rect 14185 8820 14197 8823
rect 13872 8792 14197 8820
rect 13872 8780 13878 8792
rect 14185 8789 14197 8792
rect 14231 8789 14243 8823
rect 14185 8783 14243 8789
rect 14645 8823 14703 8829
rect 14645 8789 14657 8823
rect 14691 8820 14703 8823
rect 14918 8820 14924 8832
rect 14691 8792 14924 8820
rect 14691 8789 14703 8792
rect 14645 8783 14703 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 3142 8616 3148 8628
rect 2740 8588 3148 8616
rect 2740 8576 2746 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 8846 8616 8852 8628
rect 8807 8588 8852 8616
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9324 8588 9904 8616
rect 6908 8551 6966 8557
rect 6908 8517 6920 8551
rect 6954 8548 6966 8551
rect 7098 8548 7104 8560
rect 6954 8520 7104 8548
rect 6954 8517 6966 8520
rect 6908 8511 6966 8517
rect 7098 8508 7104 8520
rect 7156 8508 7162 8560
rect 9324 8548 9352 8588
rect 8772 8520 9352 8548
rect 9876 8548 9904 8588
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10008 8588 10425 8616
rect 10008 8576 10014 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 10413 8579 10471 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12802 8616 12808 8628
rect 12763 8588 12808 8616
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 13998 8576 14004 8588
rect 14056 8616 14062 8628
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14056 8588 14565 8616
rect 14056 8576 14062 8588
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14918 8616 14924 8628
rect 14879 8588 14924 8616
rect 14553 8579 14611 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15194 8616 15200 8628
rect 15155 8588 15200 8616
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 11698 8548 11704 8560
rect 9876 8520 11704 8548
rect 2860 8483 2918 8489
rect 2860 8449 2872 8483
rect 2906 8480 2918 8483
rect 4154 8480 4160 8492
rect 2906 8452 4160 8480
rect 2906 8449 2918 8452
rect 2860 8443 2918 8449
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 4249 8483 4307 8489
rect 4249 8480 4261 8483
rect 4212 8452 4261 8480
rect 4212 8440 4218 8452
rect 4249 8449 4261 8452
rect 4295 8449 4307 8483
rect 6638 8480 6644 8492
rect 6599 8452 6644 8480
rect 4249 8443 4307 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 8772 8480 8800 8520
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 11885 8551 11943 8557
rect 11885 8517 11897 8551
rect 11931 8548 11943 8551
rect 13170 8548 13176 8560
rect 11931 8520 13176 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 13170 8508 13176 8520
rect 13228 8508 13234 8560
rect 13906 8548 13912 8560
rect 13819 8520 13912 8548
rect 13906 8508 13912 8520
rect 13964 8548 13970 8560
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 13964 8520 14473 8548
rect 13964 8508 13970 8520
rect 14461 8517 14473 8520
rect 14507 8548 14519 8551
rect 14826 8548 14832 8560
rect 14507 8520 14832 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 6748 8452 8800 8480
rect 2130 8372 2136 8424
rect 2188 8412 2194 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2188 8384 2605 8412
rect 2188 8372 2194 8384
rect 2593 8381 2605 8384
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 2608 8276 2636 8375
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 6748 8412 6776 8452
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8904 8452 9045 8480
rect 8904 8440 8910 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9289 8483 9347 8489
rect 9289 8480 9301 8483
rect 9033 8443 9091 8449
rect 9140 8452 9301 8480
rect 5868 8384 6776 8412
rect 5868 8372 5874 8384
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 9140 8412 9168 8452
rect 9289 8449 9301 8452
rect 9335 8449 9347 8483
rect 9289 8443 9347 8449
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12894 8480 12900 8492
rect 12023 8452 12900 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 7984 8384 9168 8412
rect 7984 8372 7990 8384
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 10100 8384 12081 8412
rect 10100 8372 10106 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 14277 8415 14335 8421
rect 14277 8412 14289 8415
rect 13412 8384 14289 8412
rect 13412 8372 13418 8384
rect 14277 8381 14289 8384
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 14792 8384 15025 8412
rect 14792 8372 14798 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 15013 8375 15071 8381
rect 3878 8344 3884 8356
rect 3528 8316 3884 8344
rect 3528 8276 3556 8316
rect 3878 8304 3884 8316
rect 3936 8344 3942 8356
rect 4157 8347 4215 8353
rect 4157 8344 4169 8347
rect 3936 8316 4169 8344
rect 3936 8304 3942 8316
rect 4157 8313 4169 8316
rect 4203 8344 4215 8347
rect 4246 8344 4252 8356
rect 4203 8316 4252 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4246 8304 4252 8316
rect 4304 8344 4310 8356
rect 4433 8347 4491 8353
rect 4433 8344 4445 8347
rect 4304 8316 4445 8344
rect 4304 8304 4310 8316
rect 4433 8313 4445 8316
rect 4479 8344 4491 8347
rect 5442 8344 5448 8356
rect 4479 8316 5448 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 5500 8316 5549 8344
rect 5500 8304 5506 8316
rect 5537 8313 5549 8316
rect 5583 8344 5595 8347
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 5583 8316 5733 8344
rect 5583 8313 5595 8316
rect 5537 8307 5595 8313
rect 5721 8313 5733 8316
rect 5767 8344 5779 8347
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5767 8316 5917 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 5905 8313 5917 8316
rect 5951 8344 5963 8347
rect 6089 8347 6147 8353
rect 6089 8344 6101 8347
rect 5951 8316 6101 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6089 8313 6101 8316
rect 6135 8344 6147 8347
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 6135 8316 6469 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 6457 8313 6469 8316
rect 6503 8344 6515 8347
rect 6638 8344 6644 8356
rect 6503 8316 6644 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 11440 8316 11652 8344
rect 2608 8248 3556 8276
rect 3973 8279 4031 8285
rect 3973 8245 3985 8279
rect 4019 8276 4031 8279
rect 5074 8276 5080 8288
rect 4019 8248 5080 8276
rect 4019 8245 4031 8248
rect 3973 8239 4031 8245
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 8018 8276 8024 8288
rect 7979 8248 8024 8276
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 11440 8276 11468 8316
rect 11388 8248 11468 8276
rect 11624 8276 11652 8316
rect 13998 8276 14004 8288
rect 11624 8248 14004 8276
rect 11388 8236 11394 8248
rect 13998 8236 14004 8248
rect 14056 8236 14062 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1728 8044 2145 8072
rect 1728 8032 1734 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 6178 8072 6184 8084
rect 5767 8044 6184 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7374 8072 7380 8084
rect 7239 8044 7380 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8904 8044 9045 8072
rect 8904 8032 8910 8044
rect 9033 8041 9045 8044
rect 9079 8072 9091 8075
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9079 8044 9505 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9674 8072 9680 8084
rect 9635 8044 9680 8072
rect 9493 8035 9551 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 11606 8072 11612 8084
rect 9784 8044 11612 8072
rect 3326 8004 3332 8016
rect 1596 7976 3332 8004
rect 1596 7945 1624 7976
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 9398 7964 9404 8016
rect 9456 8004 9462 8016
rect 9784 8004 9812 8044
rect 11606 8032 11612 8044
rect 11664 8072 11670 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11664 8044 12357 8072
rect 11664 8032 11670 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12345 8035 12403 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 9456 7976 9812 8004
rect 11164 7976 12940 8004
rect 9456 7964 9462 7976
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7905 1639 7939
rect 1581 7899 1639 7905
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2498 7936 2504 7948
rect 2188 7908 2504 7936
rect 2188 7896 2194 7908
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2556 7908 2789 7936
rect 2556 7896 2562 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 2777 7899 2835 7905
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 5500 7908 5825 7936
rect 5500 7896 5506 7908
rect 5813 7905 5825 7908
rect 5859 7905 5871 7939
rect 11054 7936 11060 7948
rect 11015 7908 11060 7936
rect 5813 7899 5871 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4304 7840 4353 7868
rect 4304 7828 4310 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6069 7871 6127 7877
rect 6069 7868 6081 7871
rect 5684 7840 6081 7868
rect 5684 7828 5690 7840
rect 6069 7837 6081 7840
rect 6115 7868 6127 7871
rect 9030 7868 9036 7880
rect 6115 7840 9036 7868
rect 6115 7837 6127 7840
rect 6069 7831 6127 7837
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10801 7871 10859 7877
rect 10801 7868 10813 7871
rect 9180 7840 10813 7868
rect 9180 7828 9186 7840
rect 10801 7837 10813 7840
rect 10847 7868 10859 7871
rect 11164 7868 11192 7976
rect 12912 7948 12940 7976
rect 11238 7896 11244 7948
rect 11296 7896 11302 7948
rect 12894 7896 12900 7948
rect 12952 7896 12958 7948
rect 13446 7936 13452 7948
rect 13407 7908 13452 7936
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 15105 7939 15163 7945
rect 15105 7936 15117 7939
rect 14884 7908 15117 7936
rect 14884 7896 14890 7908
rect 15105 7905 15117 7908
rect 15151 7905 15163 7939
rect 15105 7899 15163 7905
rect 10847 7840 11192 7868
rect 10847 7837 10859 7840
rect 10801 7831 10859 7837
rect 1765 7803 1823 7809
rect 1765 7769 1777 7803
rect 1811 7800 1823 7803
rect 2685 7803 2743 7809
rect 1811 7772 2268 7800
rect 1811 7769 1823 7772
rect 1765 7763 1823 7769
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 2240 7741 2268 7772
rect 2685 7769 2697 7803
rect 2731 7800 2743 7803
rect 3237 7803 3295 7809
rect 3237 7800 3249 7803
rect 2731 7772 3249 7800
rect 2731 7769 2743 7772
rect 2685 7763 2743 7769
rect 3237 7769 3249 7772
rect 3283 7800 3295 7803
rect 3878 7800 3884 7812
rect 3283 7772 3884 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 3878 7760 3884 7772
rect 3936 7760 3942 7812
rect 4614 7809 4620 7812
rect 4608 7800 4620 7809
rect 4575 7772 4620 7800
rect 4608 7763 4620 7772
rect 4614 7760 4620 7763
rect 4672 7760 4678 7812
rect 9766 7800 9772 7812
rect 7116 7772 9772 7800
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7701 2283 7735
rect 2225 7695 2283 7701
rect 2593 7735 2651 7741
rect 2593 7701 2605 7735
rect 2639 7732 2651 7735
rect 3145 7735 3203 7741
rect 3145 7732 3157 7735
rect 2639 7704 3157 7732
rect 2639 7701 2651 7704
rect 2593 7695 2651 7701
rect 3145 7701 3157 7704
rect 3191 7732 3203 7735
rect 3694 7732 3700 7744
rect 3191 7704 3700 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 7116 7732 7144 7772
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11256 7800 11284 7896
rect 12434 7800 12440 7812
rect 11112 7772 12440 7800
rect 11112 7760 11118 7772
rect 12434 7760 12440 7772
rect 12492 7800 12498 7812
rect 12802 7800 12808 7812
rect 12492 7772 12808 7800
rect 12492 7760 12498 7772
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 14274 7800 14280 7812
rect 13403 7772 14280 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7800 14979 7803
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 14967 7772 15393 7800
rect 14967 7769 14979 7772
rect 14921 7763 14979 7769
rect 15381 7769 15393 7772
rect 15427 7769 15439 7803
rect 15381 7763 15439 7769
rect 4212 7704 7144 7732
rect 4212 7692 4218 7704
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 11238 7732 11244 7744
rect 8168 7704 11244 7732
rect 8168 7692 8174 7704
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 13596 7704 14565 7732
rect 13596 7692 13602 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 15013 7735 15071 7741
rect 15013 7701 15025 7735
rect 15059 7732 15071 7735
rect 15194 7732 15200 7744
rect 15059 7704 15200 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 3234 7528 3240 7540
rect 1688 7500 3240 7528
rect 1688 7469 1716 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 4172 7500 12357 7528
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7429 1731 7463
rect 4172 7460 4200 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12676 7500 12817 7528
rect 12676 7488 12682 7500
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 13170 7528 13176 7540
rect 13131 7500 13176 7528
rect 12805 7491 12863 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 13538 7528 13544 7540
rect 13499 7500 13544 7528
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14274 7528 14280 7540
rect 14235 7500 14280 7528
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 15252 7500 15485 7528
rect 15252 7488 15258 7500
rect 15473 7497 15485 7500
rect 15519 7528 15531 7531
rect 16114 7528 16120 7540
rect 15519 7500 16120 7528
rect 15519 7497 15531 7500
rect 15473 7491 15531 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 6270 7460 6276 7472
rect 1673 7423 1731 7429
rect 1964 7432 4200 7460
rect 5000 7432 6276 7460
rect 1964 7401 1992 7432
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 1949 7355 2007 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 4453 7395 4511 7401
rect 4453 7361 4465 7395
rect 4499 7392 4511 7395
rect 4499 7364 4660 7392
rect 4499 7361 4511 7364
rect 4453 7355 4511 7361
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 4632 7324 4660 7364
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 4801 7395 4859 7401
rect 4801 7392 4813 7395
rect 4764 7364 4813 7392
rect 4764 7352 4770 7364
rect 4801 7361 4813 7364
rect 4847 7361 4859 7395
rect 5000 7392 5028 7432
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 8018 7469 8024 7472
rect 8012 7460 8024 7469
rect 7979 7432 8024 7460
rect 8012 7423 8024 7432
rect 8076 7460 8082 7472
rect 9122 7460 9128 7472
rect 8076 7432 9128 7460
rect 8018 7420 8024 7423
rect 8076 7420 8082 7432
rect 9122 7420 9128 7432
rect 9180 7420 9186 7472
rect 11238 7460 11244 7472
rect 11199 7432 11244 7460
rect 11238 7420 11244 7432
rect 11296 7460 11302 7472
rect 11885 7463 11943 7469
rect 11885 7460 11897 7463
rect 11296 7432 11897 7460
rect 11296 7420 11302 7432
rect 11885 7429 11897 7432
rect 11931 7429 11943 7463
rect 11885 7423 11943 7429
rect 11974 7420 11980 7472
rect 12032 7460 12038 7472
rect 12713 7463 12771 7469
rect 12032 7432 12112 7460
rect 12032 7420 12038 7432
rect 5074 7401 5080 7404
rect 4801 7355 4859 7361
rect 4908 7364 5028 7392
rect 4908 7324 4936 7364
rect 5068 7355 5080 7401
rect 5132 7392 5138 7404
rect 5132 7364 5168 7392
rect 5074 7352 5080 7355
rect 5132 7352 5138 7364
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 9484 7395 9542 7401
rect 9484 7392 9496 7395
rect 7892 7364 9496 7392
rect 7892 7352 7898 7364
rect 9484 7361 9496 7364
rect 9530 7392 9542 7395
rect 9530 7364 10272 7392
rect 9530 7361 9542 7364
rect 9484 7355 9542 7361
rect 4632 7296 4936 7324
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 6144 7296 6377 7324
rect 6144 7284 6150 7296
rect 6365 7293 6377 7296
rect 6411 7324 6423 7327
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 6411 7296 6561 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 6549 7293 6561 7296
rect 6595 7324 6607 7327
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 6595 7296 7573 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 7561 7293 7573 7296
rect 7607 7324 7619 7327
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7607 7296 7757 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 7098 7256 7104 7268
rect 6196 7228 7104 7256
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3329 7191 3387 7197
rect 3329 7188 3341 7191
rect 3292 7160 3341 7188
rect 3292 7148 3298 7160
rect 3329 7157 3341 7160
rect 3375 7157 3387 7191
rect 3329 7151 3387 7157
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 6196 7197 6224 7228
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5224 7160 6193 7188
rect 5224 7148 5230 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 7760 7188 7788 7287
rect 9232 7256 9260 7287
rect 8680 7228 9260 7256
rect 10244 7256 10272 7364
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 12084 7333 12112 7432
rect 12713 7429 12725 7463
rect 12759 7460 12771 7463
rect 13814 7460 13820 7472
rect 12759 7432 13820 7460
rect 12759 7429 12771 7432
rect 12713 7423 12771 7429
rect 13814 7420 13820 7432
rect 13872 7420 13878 7472
rect 14642 7392 14648 7404
rect 14603 7364 14648 7392
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11664 7296 11989 7324
rect 11664 7284 11670 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7293 12127 7327
rect 12894 7324 12900 7336
rect 12855 7296 12900 7324
rect 12069 7287 12127 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 13630 7324 13636 7336
rect 13591 7296 13636 7324
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 14734 7324 14740 7336
rect 14695 7296 14740 7324
rect 13725 7287 13783 7293
rect 13446 7256 13452 7268
rect 10244 7228 13452 7256
rect 8680 7200 8708 7228
rect 13446 7216 13452 7228
rect 13504 7256 13510 7268
rect 13740 7256 13768 7287
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 14826 7284 14832 7336
rect 14884 7324 14890 7336
rect 14884 7296 14929 7324
rect 14884 7284 14890 7296
rect 13504 7228 13768 7256
rect 13504 7216 13510 7228
rect 8662 7188 8668 7200
rect 7760 7160 8668 7188
rect 6181 7151 6239 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9125 7191 9183 7197
rect 9125 7157 9137 7191
rect 9171 7188 9183 7191
rect 9214 7188 9220 7200
rect 9171 7160 9220 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10192 7160 10609 7188
rect 10192 7148 10198 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 11514 7188 11520 7200
rect 11475 7160 11520 7188
rect 10597 7151 10655 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7188 15255 7191
rect 15286 7188 15292 7200
rect 15243 7160 15292 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15286 7148 15292 7160
rect 15344 7188 15350 7200
rect 15654 7188 15660 7200
rect 15344 7160 15660 7188
rect 15344 7148 15350 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 4154 6984 4160 6996
rect 2556 6956 4160 6984
rect 2556 6944 2562 6956
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 6086 6984 6092 6996
rect 4856 6956 6092 6984
rect 4856 6944 4862 6956
rect 6086 6944 6092 6956
rect 6144 6984 6150 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6144 6956 6561 6984
rect 6144 6944 6150 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 3602 6848 3608 6860
rect 2731 6820 3608 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2516 6780 2544 6811
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 6564 6848 6592 6947
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 7524 6956 7696 6984
rect 7524 6944 7530 6956
rect 7668 6916 7696 6956
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7892 6956 8125 6984
rect 7892 6944 7898 6956
rect 8113 6953 8125 6956
rect 8159 6953 8171 6987
rect 8662 6984 8668 6996
rect 8623 6956 8668 6984
rect 8113 6947 8171 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10321 6987 10379 6993
rect 10321 6984 10333 6987
rect 10284 6956 10333 6984
rect 10284 6944 10290 6956
rect 10321 6953 10333 6956
rect 10367 6953 10379 6987
rect 10321 6947 10379 6953
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12124 6956 13584 6984
rect 12124 6944 12130 6956
rect 7668 6888 8248 6916
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 6564 6820 6745 6848
rect 6733 6817 6745 6820
rect 6779 6817 6791 6851
rect 6733 6811 6791 6817
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2516 6752 2973 6780
rect 2961 6749 2973 6752
rect 3007 6780 3019 6783
rect 3510 6780 3516 6792
rect 3007 6752 3516 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4448 6752 4629 6780
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 3145 6715 3203 6721
rect 3145 6712 3157 6715
rect 2455 6684 3157 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 3145 6681 3157 6684
rect 3191 6712 3203 6715
rect 3418 6712 3424 6724
rect 3191 6684 3424 6712
rect 3191 6681 3203 6684
rect 3145 6675 3203 6681
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4448 6721 4476 6752
rect 4617 6749 4629 6752
rect 4663 6780 4675 6783
rect 4706 6780 4712 6792
rect 4663 6752 4712 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 4884 6783 4942 6789
rect 4884 6749 4896 6783
rect 4930 6780 4942 6783
rect 5994 6780 6000 6792
rect 4930 6752 6000 6780
rect 4930 6749 4942 6752
rect 4884 6743 4942 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 8220 6780 8248 6888
rect 8680 6848 8708 6944
rect 13556 6916 13584 6956
rect 13630 6944 13636 6996
rect 13688 6984 13694 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13688 6956 14105 6984
rect 13688 6944 13694 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 14700 6956 14933 6984
rect 14700 6944 14706 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 15102 6944 15108 6996
rect 15160 6944 15166 6996
rect 13556 6888 14136 6916
rect 14108 6860 14136 6888
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8680 6820 8953 6848
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 11514 6848 11520 6860
rect 11475 6820 11520 6848
rect 8941 6811 8999 6817
rect 11514 6808 11520 6820
rect 11572 6808 11578 6860
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 9214 6789 9220 6792
rect 9208 6780 9220 6789
rect 6512 6752 8156 6780
rect 8220 6752 9076 6780
rect 9175 6752 9220 6780
rect 6512 6740 6518 6752
rect 7006 6721 7012 6724
rect 4433 6715 4491 6721
rect 4433 6712 4445 6715
rect 4304 6684 4445 6712
rect 4304 6672 4310 6684
rect 4433 6681 4445 6684
rect 4479 6681 4491 6715
rect 7000 6712 7012 6721
rect 4433 6675 4491 6681
rect 6012 6684 7012 6712
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2041 6647 2099 6653
rect 2041 6644 2053 6647
rect 2004 6616 2053 6644
rect 2004 6604 2010 6616
rect 2041 6613 2053 6616
rect 2087 6613 2099 6647
rect 2041 6607 2099 6613
rect 2314 6604 2320 6656
rect 2372 6644 2378 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 2372 6616 3249 6644
rect 2372 6604 2378 6616
rect 3237 6613 3249 6616
rect 3283 6644 3295 6647
rect 5810 6644 5816 6656
rect 3283 6616 5816 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6012 6653 6040 6684
rect 7000 6675 7012 6684
rect 7006 6672 7012 6675
rect 7064 6672 7070 6724
rect 7650 6672 7656 6724
rect 7708 6712 7714 6724
rect 8018 6712 8024 6724
rect 7708 6684 8024 6712
rect 7708 6672 7714 6684
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 8128 6712 8156 6752
rect 9048 6712 9076 6752
rect 9208 6743 9220 6752
rect 9214 6740 9220 6743
rect 9272 6740 9278 6792
rect 11422 6780 11428 6792
rect 11383 6752 11428 6780
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11624 6712 11652 6811
rect 12544 6780 12572 6811
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 13136 6820 13277 6848
rect 13136 6808 13142 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13814 6848 13820 6860
rect 13495 6820 13820 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 13964 6820 14009 6848
rect 13964 6808 13970 6820
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14642 6848 14648 6860
rect 14603 6820 14648 6848
rect 14642 6808 14648 6820
rect 14700 6848 14706 6860
rect 14826 6848 14832 6860
rect 14700 6820 14832 6848
rect 14700 6808 14706 6820
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15120 6848 15148 6944
rect 15470 6848 15476 6860
rect 14936 6820 15148 6848
rect 15431 6820 15476 6848
rect 12710 6780 12716 6792
rect 12544 6752 12716 6780
rect 12544 6712 12572 6752
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 8128 6684 8984 6712
rect 9048 6684 11652 6712
rect 11716 6684 12572 6712
rect 13096 6712 13124 6808
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13354 6780 13360 6792
rect 13219 6752 13360 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13924 6780 13952 6808
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 13924 6752 14565 6780
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13096 6684 13645 6712
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 8202 6644 8208 6656
rect 7524 6616 8208 6644
rect 7524 6604 7530 6616
rect 8202 6604 8208 6616
rect 8260 6644 8266 6656
rect 8846 6644 8852 6656
rect 8260 6616 8852 6644
rect 8260 6604 8266 6616
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 8956 6644 8984 6684
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 8956 6616 11069 6644
rect 11057 6613 11069 6616
rect 11103 6613 11115 6647
rect 11057 6607 11115 6613
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11716 6644 11744 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 14461 6715 14519 6721
rect 14461 6712 14473 6715
rect 14056 6684 14473 6712
rect 14056 6672 14062 6684
rect 14461 6681 14473 6684
rect 14507 6712 14519 6715
rect 14936 6712 14964 6820
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15286 6780 15292 6792
rect 15068 6752 15292 6780
rect 15068 6740 15074 6752
rect 15286 6740 15292 6752
rect 15344 6780 15350 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15344 6752 15393 6780
rect 15344 6740 15350 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 14507 6684 14964 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 11882 6644 11888 6656
rect 11572 6616 11744 6644
rect 11843 6616 11888 6644
rect 11572 6604 11578 6616
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12253 6647 12311 6653
rect 12253 6644 12265 6647
rect 12124 6616 12265 6644
rect 12124 6604 12130 6616
rect 12253 6613 12265 6616
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 12345 6647 12403 6653
rect 12345 6613 12357 6647
rect 12391 6644 12403 6647
rect 12618 6644 12624 6656
rect 12391 6616 12624 6644
rect 12391 6613 12403 6616
rect 12345 6607 12403 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 12894 6644 12900 6656
rect 12851 6616 12900 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 14550 6644 14556 6656
rect 13136 6616 14556 6644
rect 13136 6604 13142 6616
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 14884 6616 15301 6644
rect 14884 6604 14890 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 3970 6440 3976 6452
rect 1964 6412 3976 6440
rect 1578 6332 1584 6384
rect 1636 6372 1642 6384
rect 1673 6375 1731 6381
rect 1673 6372 1685 6375
rect 1636 6344 1685 6372
rect 1636 6332 1642 6344
rect 1673 6341 1685 6344
rect 1719 6341 1731 6375
rect 1673 6335 1731 6341
rect 1964 6313 1992 6412
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4798 6440 4804 6452
rect 4120 6412 4804 6440
rect 4120 6400 4126 6412
rect 4798 6400 4804 6412
rect 4856 6440 4862 6452
rect 5261 6443 5319 6449
rect 5261 6440 5273 6443
rect 4856 6412 5273 6440
rect 4856 6400 4862 6412
rect 5261 6409 5273 6412
rect 5307 6409 5319 6443
rect 5261 6403 5319 6409
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 5994 6440 6000 6452
rect 5868 6412 6000 6440
rect 5868 6400 5874 6412
rect 5994 6400 6000 6412
rect 6052 6440 6058 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 6052 6412 6377 6440
rect 6052 6400 6058 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7742 6440 7748 6452
rect 7239 6412 7748 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8159 6412 8493 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8904 6412 8953 6440
rect 8904 6400 8910 6412
rect 8941 6409 8953 6412
rect 8987 6440 8999 6443
rect 9306 6440 9312 6452
rect 8987 6412 9312 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 11054 6440 11060 6452
rect 9640 6412 11060 6440
rect 9640 6400 9646 6412
rect 11054 6400 11060 6412
rect 11112 6400 11118 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12434 6440 12440 6452
rect 12299 6412 12440 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12710 6440 12716 6452
rect 12623 6412 12716 6440
rect 12710 6400 12716 6412
rect 12768 6440 12774 6452
rect 13354 6440 13360 6452
rect 12768 6412 13360 6440
rect 12768 6400 12774 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14277 6443 14335 6449
rect 14277 6409 14289 6443
rect 14323 6440 14335 6443
rect 14550 6440 14556 6452
rect 14323 6412 14556 6440
rect 14323 6409 14335 6412
rect 14277 6403 14335 6409
rect 14550 6400 14556 6412
rect 14608 6440 14614 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14608 6412 15117 6440
rect 14608 6400 14614 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15344 6412 15577 6440
rect 15344 6400 15350 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 2314 6332 2320 6384
rect 2372 6372 2378 6384
rect 2501 6375 2559 6381
rect 2501 6372 2513 6375
rect 2372 6344 2513 6372
rect 2372 6332 2378 6344
rect 2501 6341 2513 6344
rect 2547 6341 2559 6375
rect 4246 6372 4252 6384
rect 2501 6335 2559 6341
rect 2976 6344 4252 6372
rect 2976 6313 3004 6344
rect 4246 6332 4252 6344
rect 4304 6332 4310 6384
rect 6086 6372 6092 6384
rect 4724 6344 6092 6372
rect 3234 6313 3240 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 3228 6304 3240 6313
rect 3147 6276 3240 6304
rect 2961 6267 3019 6273
rect 3228 6267 3240 6276
rect 3292 6304 3298 6316
rect 4724 6304 4752 6344
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 7006 6332 7012 6384
rect 7064 6372 7070 6384
rect 14642 6372 14648 6384
rect 7064 6344 14648 6372
rect 7064 6332 7070 6344
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 3292 6276 4752 6304
rect 8021 6307 8079 6313
rect 3234 6264 3240 6267
rect 3292 6264 3298 6276
rect 8021 6273 8033 6307
rect 8067 6304 8079 6307
rect 8294 6304 8300 6316
rect 8067 6276 8300 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8846 6304 8852 6316
rect 8759 6276 8852 6304
rect 8846 6264 8852 6276
rect 8904 6304 8910 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 8904 6276 9413 6304
rect 8904 6264 8910 6276
rect 9401 6273 9413 6276
rect 9447 6304 9459 6307
rect 11238 6304 11244 6316
rect 9447 6276 11244 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 11238 6264 11244 6276
rect 11296 6304 11302 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11296 6276 11897 6304
rect 11296 6264 11302 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 12618 6304 12624 6316
rect 12492 6276 12624 6304
rect 12492 6264 12498 6276
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 12802 6264 12808 6316
rect 12860 6304 12866 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 12860 6276 14381 6304
rect 12860 6264 12866 6276
rect 14369 6273 14381 6276
rect 14415 6304 14427 6307
rect 15197 6307 15255 6313
rect 15197 6304 15209 6307
rect 14415 6276 15209 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 15197 6273 15209 6276
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 2225 6239 2283 6245
rect 2225 6236 2237 6239
rect 1544 6208 2237 6236
rect 1544 6196 1550 6208
rect 2225 6205 2237 6208
rect 2271 6205 2283 6239
rect 2225 6199 2283 6205
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2590 6236 2596 6248
rect 2455 6208 2596 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2240 6168 2268 6199
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4120 6208 4905 6236
rect 4120 6196 4126 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5626 6236 5632 6248
rect 5123 6208 5632 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6205 6975 6239
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 6917 6199 6975 6205
rect 2498 6168 2504 6180
rect 2240 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 4614 6168 4620 6180
rect 4387 6140 4620 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 4614 6128 4620 6140
rect 4672 6168 4678 6180
rect 5534 6168 5540 6180
rect 4672 6140 5540 6168
rect 4672 6128 4678 6140
rect 5534 6128 5540 6140
rect 5592 6128 5598 6180
rect 6932 6168 6960 6199
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 7374 6168 7380 6180
rect 6932 6140 7380 6168
rect 7374 6128 7380 6140
rect 7432 6168 7438 6180
rect 8220 6168 8248 6199
rect 9030 6196 9036 6248
rect 9088 6236 9094 6248
rect 9088 6208 9133 6236
rect 9088 6196 9094 6208
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 9364 6208 11069 6236
rect 9364 6196 9370 6208
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 10042 6168 10048 6180
rect 7432 6140 10048 6168
rect 7432 6128 7438 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 11072 6168 11100 6199
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11609 6239 11667 6245
rect 11609 6236 11621 6239
rect 11480 6208 11621 6236
rect 11480 6196 11486 6208
rect 11609 6205 11621 6208
rect 11655 6205 11667 6239
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11609 6199 11667 6205
rect 11716 6208 11805 6236
rect 11716 6168 11744 6208
rect 11793 6205 11805 6208
rect 11839 6205 11851 6239
rect 13446 6236 13452 6248
rect 13407 6208 13452 6236
rect 11793 6199 11851 6205
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13998 6236 14004 6248
rect 13648 6208 14004 6236
rect 13648 6168 13676 6208
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 15102 6236 15108 6248
rect 14148 6208 15108 6236
rect 14148 6196 14154 6208
rect 15102 6196 15108 6208
rect 15160 6236 15166 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 15160 6208 15301 6236
rect 15160 6196 15166 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 11072 6140 11744 6168
rect 11808 6140 13676 6168
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 3234 6100 3240 6112
rect 2915 6072 3240 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 4706 6100 4712 6112
rect 4479 6072 4712 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 7558 6100 7564 6112
rect 7519 6072 7564 6100
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 7708 6072 7753 6100
rect 7708 6060 7714 6072
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 11808 6100 11836 6140
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 13780 6140 14749 6168
rect 13780 6128 13786 6140
rect 14737 6137 14749 6140
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 11756 6072 11836 6100
rect 11756 6060 11762 6072
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12710 6100 12716 6112
rect 11940 6072 12716 6100
rect 11940 6060 11946 6072
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12860 6072 12909 6100
rect 12860 6060 12866 6072
rect 12897 6069 12909 6072
rect 12943 6100 12955 6103
rect 13538 6100 13544 6112
rect 12943 6072 13544 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13538 6060 13544 6072
rect 13596 6060 13602 6112
rect 14645 6103 14703 6109
rect 14645 6069 14657 6103
rect 14691 6100 14703 6103
rect 14826 6100 14832 6112
rect 14691 6072 14832 6100
rect 14691 6069 14703 6072
rect 14645 6063 14703 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1489 5899 1547 5905
rect 1489 5865 1501 5899
rect 1535 5896 1547 5899
rect 1670 5896 1676 5908
rect 1535 5868 1676 5896
rect 1535 5865 1547 5868
rect 1489 5859 1547 5865
rect 1670 5856 1676 5868
rect 1728 5856 1734 5908
rect 2590 5896 2596 5908
rect 2551 5868 2596 5896
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 4798 5896 4804 5908
rect 2746 5868 4804 5896
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 2056 5800 2421 5828
rect 1946 5760 1952 5772
rect 1907 5732 1952 5760
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2056 5692 2084 5800
rect 2409 5797 2421 5800
rect 2455 5828 2467 5831
rect 2746 5828 2774 5868
rect 4798 5856 4804 5868
rect 4856 5896 4862 5908
rect 5074 5896 5080 5908
rect 4856 5868 5080 5896
rect 4856 5856 4862 5868
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 7800 5868 8125 5896
rect 7800 5856 7806 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9306 5896 9312 5908
rect 8435 5868 9312 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5896 9735 5899
rect 9766 5896 9772 5908
rect 9723 5868 9772 5896
rect 9723 5865 9735 5868
rect 9677 5859 9735 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 12124 5868 12265 5896
rect 12124 5856 12130 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13320 5868 14105 5896
rect 13320 5856 13326 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14792 5868 14933 5896
rect 14792 5856 14798 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 5902 5828 5908 5840
rect 2455 5800 2774 5828
rect 3252 5800 5908 5828
rect 2455 5797 2467 5800
rect 2409 5791 2467 5797
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 3252 5769 3280 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 6104 5800 11652 5828
rect 6104 5772 6132 5800
rect 3237 5763 3295 5769
rect 2188 5732 2233 5760
rect 2188 5720 2194 5732
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3237 5723 3295 5729
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4430 5760 4436 5772
rect 3660 5732 4436 5760
rect 3660 5720 3666 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4706 5760 4712 5772
rect 4667 5732 4712 5760
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4893 5763 4951 5769
rect 4893 5729 4905 5763
rect 4939 5760 4951 5763
rect 5350 5760 5356 5772
rect 4939 5732 5356 5760
rect 4939 5729 4951 5732
rect 4893 5723 4951 5729
rect 5350 5720 5356 5732
rect 5408 5760 5414 5772
rect 5810 5760 5816 5772
rect 5408 5732 5816 5760
rect 5408 5720 5414 5732
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 6086 5760 6092 5772
rect 5999 5732 6092 5760
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6328 5732 6837 5760
rect 6328 5720 6334 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7340 5732 7389 5760
rect 7340 5720 7346 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7650 5760 7656 5772
rect 7607 5732 7656 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 1903 5664 2084 5692
rect 3513 5695 3571 5701
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 6733 5695 6791 5701
rect 6733 5692 6745 5695
rect 3559 5664 6745 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2832 5596 2973 5624
rect 2832 5584 2838 5596
rect 2961 5593 2973 5596
rect 3007 5624 3019 5627
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 3007 5596 3801 5624
rect 3007 5593 3019 5596
rect 2961 5587 3019 5593
rect 3789 5593 3801 5596
rect 3835 5593 3847 5627
rect 3789 5587 3847 5593
rect 3053 5559 3111 5565
rect 3053 5525 3065 5559
rect 3099 5556 3111 5559
rect 3896 5556 3924 5664
rect 6733 5661 6745 5664
rect 6779 5692 6791 5695
rect 7392 5692 7420 5723
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 7984 5732 9444 5760
rect 7984 5720 7990 5732
rect 9122 5692 9128 5704
rect 6779 5664 7328 5692
rect 7392 5664 9128 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 5813 5627 5871 5633
rect 5813 5593 5825 5627
rect 5859 5624 5871 5627
rect 5994 5624 6000 5636
rect 5859 5596 6000 5624
rect 5859 5593 5871 5596
rect 5813 5587 5871 5593
rect 5994 5584 6000 5596
rect 6052 5584 6058 5636
rect 6641 5627 6699 5633
rect 6641 5593 6653 5627
rect 6687 5593 6699 5627
rect 7300 5624 7328 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9416 5692 9444 5732
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 9548 5732 10241 5760
rect 9548 5720 9554 5732
rect 10229 5729 10241 5732
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 10318 5720 10324 5772
rect 10376 5760 10382 5772
rect 11057 5763 11115 5769
rect 11057 5760 11069 5763
rect 10376 5732 11069 5760
rect 10376 5720 10382 5732
rect 11057 5729 11069 5732
rect 11103 5760 11115 5763
rect 11330 5760 11336 5772
rect 11103 5732 11336 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11514 5760 11520 5772
rect 11475 5732 11520 5760
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 11624 5760 11652 5800
rect 11790 5788 11796 5840
rect 11848 5828 11854 5840
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 11848 5800 12173 5828
rect 11848 5788 11854 5800
rect 12161 5797 12173 5800
rect 12207 5797 12219 5831
rect 13814 5828 13820 5840
rect 12161 5791 12219 5797
rect 12268 5800 13820 5828
rect 12268 5760 12296 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 11624 5732 12296 5760
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12400 5732 12909 5760
rect 12400 5720 12406 5732
rect 12897 5729 12909 5732
rect 12943 5760 12955 5763
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 12943 5732 13645 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 14642 5760 14648 5772
rect 14603 5732 14648 5760
rect 13633 5723 13691 5729
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 15470 5760 15476 5772
rect 15431 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 9582 5692 9588 5704
rect 9416 5664 9588 5692
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 13538 5692 13544 5704
rect 11747 5664 13124 5692
rect 13499 5664 13544 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 7466 5624 7472 5636
rect 7300 5596 7472 5624
rect 6641 5587 6699 5593
rect 4246 5556 4252 5568
rect 3099 5528 3924 5556
rect 4207 5528 4252 5556
rect 3099 5525 3111 5528
rect 3053 5519 3111 5525
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4614 5556 4620 5568
rect 4575 5528 4620 5556
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 5951 5528 6285 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6273 5525 6285 5528
rect 6319 5525 6331 5559
rect 6273 5519 6331 5525
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6656 5556 6684 5587
rect 7466 5584 7472 5596
rect 7524 5584 7530 5636
rect 7558 5584 7564 5636
rect 7616 5624 7622 5636
rect 7653 5627 7711 5633
rect 7653 5624 7665 5627
rect 7616 5596 7665 5624
rect 7616 5584 7622 5596
rect 7653 5593 7665 5596
rect 7699 5593 7711 5627
rect 8846 5624 8852 5636
rect 7653 5587 7711 5593
rect 7760 5596 8852 5624
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 6420 5528 7205 5556
rect 6420 5516 6426 5528
rect 7193 5525 7205 5528
rect 7239 5556 7251 5559
rect 7760 5556 7788 5596
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 10045 5627 10103 5633
rect 10045 5593 10057 5627
rect 10091 5624 10103 5627
rect 10778 5624 10784 5636
rect 10091 5596 10784 5624
rect 10091 5593 10103 5596
rect 10045 5587 10103 5593
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 11606 5584 11612 5636
rect 11664 5624 11670 5636
rect 11793 5627 11851 5633
rect 11793 5624 11805 5627
rect 11664 5596 11805 5624
rect 11664 5584 11670 5596
rect 11793 5593 11805 5596
rect 11839 5593 11851 5627
rect 11793 5587 11851 5593
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12124 5596 12725 5624
rect 12124 5584 12130 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 12713 5587 12771 5593
rect 7239 5528 7788 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 8021 5559 8079 5565
rect 8021 5556 8033 5559
rect 7892 5528 8033 5556
rect 7892 5516 7898 5528
rect 8021 5525 8033 5528
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 9766 5556 9772 5568
rect 9272 5528 9772 5556
rect 9272 5516 9278 5528
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 10137 5559 10195 5565
rect 10137 5525 10149 5559
rect 10183 5556 10195 5559
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 10183 5528 10517 5556
rect 10183 5525 10195 5528
rect 10137 5519 10195 5525
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 10870 5556 10876 5568
rect 10831 5528 10876 5556
rect 10505 5519 10563 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11020 5528 11065 5556
rect 11020 5516 11026 5528
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 13096 5565 13124 5664
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 14366 5652 14372 5704
rect 14424 5692 14430 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14424 5664 15301 5692
rect 14424 5652 14430 5664
rect 15289 5661 15301 5664
rect 15335 5692 15347 5695
rect 15746 5692 15752 5704
rect 15335 5664 15752 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 13412 5596 13461 5624
rect 13412 5584 13418 5596
rect 13449 5593 13461 5596
rect 13495 5593 13507 5627
rect 13449 5587 13507 5593
rect 13081 5559 13139 5565
rect 12676 5528 12721 5556
rect 12676 5516 12682 5528
rect 13081 5525 13093 5559
rect 13127 5525 13139 5559
rect 13081 5519 13139 5525
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14461 5559 14519 5565
rect 14461 5556 14473 5559
rect 13964 5528 14473 5556
rect 13964 5516 13970 5528
rect 14461 5525 14473 5528
rect 14507 5525 14519 5559
rect 14461 5519 14519 5525
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14608 5528 14653 5556
rect 14608 5516 14614 5528
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15381 5559 15439 5565
rect 15381 5556 15393 5559
rect 15344 5528 15393 5556
rect 15344 5516 15350 5528
rect 15381 5525 15393 5528
rect 15427 5556 15439 5559
rect 16114 5556 16120 5568
rect 15427 5528 16120 5556
rect 15427 5525 15439 5528
rect 15381 5519 15439 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 4062 5352 4068 5364
rect 3835 5324 4068 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4304 5324 4629 5352
rect 4304 5312 4310 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5537 5355 5595 5361
rect 5537 5352 5549 5355
rect 5500 5324 5549 5352
rect 5500 5312 5506 5324
rect 5537 5321 5549 5324
rect 5583 5321 5595 5355
rect 5537 5315 5595 5321
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 6043 5324 6837 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 7156 5324 7481 5352
rect 7156 5312 7162 5324
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7926 5352 7932 5364
rect 7887 5324 7932 5352
rect 7469 5315 7527 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8352 5324 8493 5352
rect 8352 5312 8358 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 8481 5315 8539 5321
rect 8864 5324 9689 5352
rect 2682 5284 2688 5296
rect 2643 5256 2688 5284
rect 2682 5244 2688 5256
rect 2740 5244 2746 5296
rect 3602 5284 3608 5296
rect 3252 5256 3608 5284
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3142 5216 3148 5228
rect 3007 5188 3148 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3252 5157 3280 5256
rect 3602 5244 3608 5256
rect 3660 5244 3666 5296
rect 3973 5287 4031 5293
rect 3973 5253 3985 5287
rect 4019 5284 4031 5287
rect 6730 5284 6736 5296
rect 4019 5256 5764 5284
rect 6691 5256 6736 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 3988 5216 4016 5247
rect 3476 5188 4016 5216
rect 4525 5219 4583 5225
rect 3476 5176 3482 5188
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4706 5216 4712 5228
rect 4571 5188 4712 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5500 5188 5641 5216
rect 5500 5176 5506 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5736 5216 5764 5256
rect 6730 5244 6736 5256
rect 6788 5244 6794 5296
rect 8864 5284 8892 5324
rect 9677 5321 9689 5324
rect 9723 5352 9735 5355
rect 10045 5355 10103 5361
rect 9723 5324 9996 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 6831 5256 8892 5284
rect 8941 5287 8999 5293
rect 6831 5216 6859 5256
rect 8941 5253 8953 5287
rect 8987 5284 8999 5287
rect 9306 5284 9312 5296
rect 8987 5256 9312 5284
rect 8987 5253 8999 5256
rect 8941 5247 8999 5253
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 9582 5284 9588 5296
rect 9543 5256 9588 5284
rect 9582 5244 9588 5256
rect 9640 5244 9646 5296
rect 9968 5284 9996 5324
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10091 5324 10425 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10873 5355 10931 5361
rect 10560 5324 10605 5352
rect 10560 5312 10566 5324
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 10962 5352 10968 5364
rect 10919 5324 10968 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11606 5352 11612 5364
rect 11567 5324 11612 5352
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 11882 5352 11888 5364
rect 11843 5324 11888 5352
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12710 5352 12716 5364
rect 12671 5324 12716 5352
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 13446 5352 13452 5364
rect 13403 5324 13452 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 13906 5352 13912 5364
rect 13867 5324 13912 5352
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 14424 5324 14473 5352
rect 14424 5312 14430 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14645 5355 14703 5361
rect 14645 5352 14657 5355
rect 14608 5324 14657 5352
rect 14608 5312 14614 5324
rect 14645 5321 14657 5324
rect 14691 5321 14703 5355
rect 15010 5352 15016 5364
rect 14923 5324 15016 5352
rect 14645 5315 14703 5321
rect 15010 5312 15016 5324
rect 15068 5352 15074 5364
rect 15930 5352 15936 5364
rect 15068 5324 15936 5352
rect 15068 5312 15074 5324
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 10134 5284 10140 5296
rect 9968 5256 10140 5284
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 13538 5244 13544 5296
rect 13596 5284 13602 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13596 5256 14197 5284
rect 13596 5244 13602 5256
rect 14185 5253 14197 5256
rect 14231 5284 14243 5287
rect 15194 5284 15200 5296
rect 14231 5256 15200 5284
rect 14231 5253 14243 5256
rect 14185 5247 14243 5253
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 15470 5244 15476 5296
rect 15528 5244 15534 5296
rect 5736 5188 6859 5216
rect 5629 5179 5687 5185
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7064 5188 7849 5216
rect 7064 5176 7070 5188
rect 7837 5185 7849 5188
rect 7883 5216 7895 5219
rect 8202 5216 8208 5228
rect 7883 5188 8208 5216
rect 7883 5185 7895 5188
rect 7837 5179 7895 5185
rect 8202 5176 8208 5188
rect 8260 5216 8266 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8260 5188 8309 5216
rect 8260 5176 8266 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8846 5216 8852 5228
rect 8807 5188 8852 5216
rect 8297 5179 8355 5185
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10560 5188 10977 5216
rect 10560 5176 10566 5188
rect 10965 5185 10977 5188
rect 11011 5216 11023 5219
rect 11606 5216 11612 5228
rect 11011 5188 11612 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 14274 5216 14280 5228
rect 12124 5188 14280 5216
rect 12124 5176 12130 5188
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14734 5216 14740 5228
rect 14415 5188 14740 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14734 5176 14740 5188
rect 14792 5216 14798 5228
rect 15010 5216 15016 5228
rect 14792 5188 15016 5216
rect 14792 5176 14798 5188
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15488 5216 15516 5244
rect 15212 5188 15516 5216
rect 3237 5151 3295 5157
rect 3237 5117 3249 5151
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3344 5012 3372 5111
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 4801 5151 4859 5157
rect 4028 5120 4292 5148
rect 4028 5108 4034 5120
rect 3510 5012 3516 5024
rect 3344 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 5012 3574 5024
rect 3970 5012 3976 5024
rect 3568 4984 3976 5012
rect 3568 4972 3574 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4120 4984 4169 5012
rect 4120 4972 4126 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 4264 5012 4292 5120
rect 4801 5117 4813 5151
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5534 5148 5540 5160
rect 5399 5120 5540 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 4816 5080 4844 5111
rect 5534 5108 5540 5120
rect 5592 5148 5598 5160
rect 5902 5148 5908 5160
rect 5592 5120 5908 5148
rect 5592 5108 5598 5120
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6236 5120 6929 5148
rect 6236 5108 6242 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7466 5148 7472 5160
rect 7331 5120 7472 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 5718 5080 5724 5092
rect 4816 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 8128 5080 8156 5111
rect 9030 5108 9036 5160
rect 9088 5148 9094 5160
rect 9398 5148 9404 5160
rect 9088 5120 9133 5148
rect 9359 5120 9404 5148
rect 9088 5108 9094 5120
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9824 5120 10241 5148
rect 9824 5108 9830 5120
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 11790 5148 11796 5160
rect 10275 5120 11796 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 11790 5108 11796 5120
rect 11848 5148 11854 5160
rect 13446 5148 13452 5160
rect 11848 5120 12756 5148
rect 13407 5120 13452 5148
rect 11848 5108 11854 5120
rect 9048 5080 9076 5108
rect 6052 5052 8055 5080
rect 8128 5052 9076 5080
rect 6052 5040 6058 5052
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 4264 4984 6377 5012
rect 4157 4975 4215 4981
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 8027 5012 8055 5052
rect 10134 5040 10140 5092
rect 10192 5080 10198 5092
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 10192 5052 11253 5080
rect 10192 5040 10198 5052
rect 11241 5049 11253 5052
rect 11287 5080 11299 5083
rect 12066 5080 12072 5092
rect 11287 5052 12072 5080
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 12066 5040 12072 5052
rect 12124 5040 12130 5092
rect 8386 5012 8392 5024
rect 8027 4984 8392 5012
rect 6365 4975 6423 4981
rect 8386 4972 8392 4984
rect 8444 5012 8450 5024
rect 9306 5012 9312 5024
rect 8444 4984 9312 5012
rect 8444 4972 8450 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12618 5012 12624 5024
rect 12032 4984 12624 5012
rect 12032 4972 12038 4984
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 12728 5012 12756 5120
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 12860 5052 13001 5080
rect 12860 5040 12866 5052
rect 12989 5049 13001 5052
rect 13035 5049 13047 5083
rect 12989 5043 13047 5049
rect 13556 5012 13584 5111
rect 13630 5108 13636 5160
rect 13688 5148 13694 5160
rect 15212 5157 15240 5188
rect 15105 5151 15163 5157
rect 15105 5148 15117 5151
rect 13688 5120 15117 5148
rect 13688 5108 13694 5120
rect 15105 5117 15117 5120
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5117 15255 5151
rect 15197 5111 15255 5117
rect 15286 5108 15292 5160
rect 15344 5148 15350 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15344 5120 15485 5148
rect 15344 5108 15350 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 12728 4984 13584 5012
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 4154 4808 4160 4820
rect 4115 4780 4160 4808
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 5132 4780 5181 4808
rect 5132 4768 5138 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5442 4808 5448 4820
rect 5403 4780 5448 4808
rect 5169 4771 5227 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 6365 4811 6423 4817
rect 6365 4808 6377 4811
rect 6104 4780 6377 4808
rect 3970 4740 3976 4752
rect 3931 4712 3976 4740
rect 3970 4700 3976 4712
rect 4028 4700 4034 4752
rect 6104 4740 6132 4780
rect 6365 4777 6377 4780
rect 6411 4808 6423 4811
rect 7742 4808 7748 4820
rect 6411 4780 7748 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8202 4808 8208 4820
rect 7984 4780 8208 4808
rect 7984 4768 7990 4780
rect 8202 4768 8208 4780
rect 8260 4808 8266 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8260 4780 8493 4808
rect 8260 4768 8266 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 8904 4780 9321 4808
rect 8904 4768 8910 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 9309 4771 9367 4777
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 10870 4808 10876 4820
rect 10735 4780 10876 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 13630 4808 13636 4820
rect 12452 4780 13492 4808
rect 13591 4780 13636 4808
rect 5920 4712 6132 4740
rect 3234 4672 3240 4684
rect 3195 4644 3240 4672
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 3384 4644 3429 4672
rect 3384 4632 3390 4644
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4212 4644 4905 4672
rect 4212 4632 4218 4644
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 5920 4672 5948 4712
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 6972 4712 7972 4740
rect 6972 4700 6978 4712
rect 6086 4672 6092 4684
rect 4893 4635 4951 4641
rect 5828 4644 5948 4672
rect 6047 4644 6092 4672
rect 2130 4604 2136 4616
rect 2091 4576 2136 4604
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 4246 4604 4252 4616
rect 3200 4576 4252 4604
rect 3200 4564 3206 4576
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 5074 4604 5080 4616
rect 4755 4576 5080 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5828 4613 5856 4644
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 7834 4672 7840 4684
rect 7795 4644 7840 4672
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 7944 4681 7972 4712
rect 8110 4700 8116 4752
rect 8168 4740 8174 4752
rect 8665 4743 8723 4749
rect 8665 4740 8677 4743
rect 8168 4712 8677 4740
rect 8168 4700 8174 4712
rect 8665 4709 8677 4712
rect 8711 4740 8723 4743
rect 10318 4740 10324 4752
rect 8711 4712 10324 4740
rect 8711 4709 8723 4712
rect 8665 4703 8723 4709
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 10778 4740 10784 4752
rect 10739 4712 10784 4740
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 11974 4700 11980 4752
rect 12032 4740 12038 4752
rect 12452 4740 12480 4780
rect 12032 4712 12480 4740
rect 12032 4700 12038 4712
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 13078 4740 13084 4752
rect 12584 4712 13084 4740
rect 12584 4700 12590 4712
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 13464 4749 13492 4780
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13449 4743 13507 4749
rect 13449 4709 13461 4743
rect 13495 4740 13507 4743
rect 13495 4712 15608 4740
rect 13495 4709 13507 4712
rect 13449 4703 13507 4709
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4641 7987 4675
rect 8386 4672 8392 4684
rect 8347 4644 8392 4672
rect 7929 4635 7987 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9272 4644 10057 4672
rect 9272 4632 9278 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 10045 4635 10103 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 12158 4672 12164 4684
rect 12119 4644 12164 4672
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12406 4644 13001 4672
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 7745 4607 7803 4613
rect 5960 4576 7512 4604
rect 5960 4564 5966 4576
rect 1854 4536 1860 4548
rect 1815 4508 1860 4536
rect 1854 4496 1860 4508
rect 1912 4496 1918 4548
rect 2222 4496 2228 4548
rect 2280 4536 2286 4548
rect 7484 4536 7512 4576
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8294 4604 8300 4616
rect 7791 4576 8300 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 9088 4576 9137 4604
rect 9088 4564 9094 4576
rect 9125 4573 9137 4576
rect 9171 4604 9183 4607
rect 9582 4604 9588 4616
rect 9171 4576 9588 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9858 4564 9864 4616
rect 9916 4604 9922 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 9916 4576 10333 4604
rect 9916 4564 9922 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4604 11207 4607
rect 11238 4604 11244 4616
rect 11195 4576 11244 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 12406 4604 12434 4644
rect 12989 4641 13001 4644
rect 13035 4641 13047 4675
rect 12989 4635 13047 4641
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 13872 4644 14657 4672
rect 13872 4632 13878 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15160 4644 15485 4672
rect 15160 4632 15166 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15473 4635 15531 4641
rect 12894 4604 12900 4616
rect 11348 4576 12434 4604
rect 12855 4576 12900 4604
rect 11348 4536 11376 4576
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 14550 4604 14556 4616
rect 14511 4576 14556 4604
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15580 4604 15608 4712
rect 15654 4604 15660 4616
rect 15427 4576 15660 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15654 4564 15660 4576
rect 15712 4604 15718 4616
rect 16390 4604 16396 4616
rect 15712 4576 16396 4604
rect 15712 4564 15718 4576
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 2280 4508 7420 4536
rect 7484 4508 11376 4536
rect 11977 4539 12035 4545
rect 2280 4496 2286 4508
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3142 4468 3148 4480
rect 2832 4440 2877 4468
rect 3103 4440 3148 4468
rect 2832 4428 2838 4440
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 4341 4471 4399 4477
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 4430 4468 4436 4480
rect 4387 4440 4436 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 4706 4468 4712 4480
rect 4580 4440 4712 4468
rect 4580 4428 4586 4440
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 5074 4468 5080 4480
rect 4847 4440 5080 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5905 4471 5963 4477
rect 5905 4437 5917 4471
rect 5951 4468 5963 4471
rect 6270 4468 6276 4480
rect 5951 4440 6276 4468
rect 5951 4437 5963 4440
rect 5905 4431 5963 4437
rect 6270 4428 6276 4440
rect 6328 4468 6334 4480
rect 7392 4477 7420 4508
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12710 4536 12716 4548
rect 12023 4508 12716 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 12805 4539 12863 4545
rect 12805 4505 12817 4539
rect 12851 4536 12863 4539
rect 13909 4539 13967 4545
rect 12851 4508 13676 4536
rect 12851 4505 12863 4508
rect 12805 4499 12863 4505
rect 6457 4471 6515 4477
rect 6457 4468 6469 4471
rect 6328 4440 6469 4468
rect 6328 4428 6334 4440
rect 6457 4437 6469 4440
rect 6503 4437 6515 4471
rect 6457 4431 6515 4437
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4437 7435 4471
rect 7377 4431 7435 4437
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 9030 4468 9036 4480
rect 7708 4440 9036 4468
rect 7708 4428 7714 4440
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9858 4428 9864 4480
rect 9916 4468 9922 4480
rect 10229 4471 10287 4477
rect 10229 4468 10241 4471
rect 9916 4440 10241 4468
rect 9916 4428 9922 4440
rect 10229 4437 10241 4440
rect 10275 4437 10287 4471
rect 10229 4431 10287 4437
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 11606 4468 11612 4480
rect 11296 4440 11341 4468
rect 11567 4440 11612 4468
rect 11296 4428 11302 4440
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 13648 4468 13676 4508
rect 13909 4505 13921 4539
rect 13955 4536 13967 4539
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 13955 4508 14473 4536
rect 13955 4505 13967 4508
rect 13909 4499 13967 4505
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 14461 4499 14519 4505
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 12492 4440 12537 4468
rect 13648 4440 14105 4468
rect 12492 4428 12498 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14918 4468 14924 4480
rect 14879 4440 14924 4468
rect 14093 4431 14151 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1949 4267 2007 4273
rect 1949 4233 1961 4267
rect 1995 4264 2007 4267
rect 2130 4264 2136 4276
rect 1995 4236 2136 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 2869 4267 2927 4273
rect 2869 4233 2881 4267
rect 2915 4264 2927 4267
rect 3142 4264 3148 4276
rect 2915 4236 3148 4264
rect 2915 4233 2927 4236
rect 2869 4227 2927 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3292 4236 3337 4264
rect 3292 4224 3298 4236
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3970 4264 3976 4276
rect 3752 4236 3976 4264
rect 3752 4224 3758 4236
rect 3970 4224 3976 4236
rect 4028 4264 4034 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 4028 4236 4077 4264
rect 4028 4224 4034 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 4065 4227 4123 4233
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 4580 4236 5273 4264
rect 4580 4224 4586 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 6328 4236 6469 4264
rect 6328 4224 6334 4236
rect 6457 4233 6469 4236
rect 6503 4264 6515 4267
rect 7190 4264 7196 4276
rect 6503 4236 7196 4264
rect 6503 4233 6515 4236
rect 6457 4227 6515 4233
rect 7190 4224 7196 4236
rect 7248 4264 7254 4276
rect 7466 4264 7472 4276
rect 7248 4236 7472 4264
rect 7248 4224 7254 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4264 8079 4267
rect 8110 4264 8116 4276
rect 8067 4236 8116 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8352 4236 8493 4264
rect 8352 4224 8358 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 8941 4267 8999 4273
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 9493 4267 9551 4273
rect 9493 4264 9505 4267
rect 8987 4236 9505 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9493 4233 9505 4236
rect 9539 4233 9551 4267
rect 9493 4227 9551 4233
rect 9861 4267 9919 4273
rect 9861 4233 9873 4267
rect 9907 4264 9919 4267
rect 9950 4264 9956 4276
rect 9907 4236 9956 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 9950 4224 9956 4236
rect 10008 4264 10014 4276
rect 10321 4267 10379 4273
rect 10321 4264 10333 4267
rect 10008 4236 10333 4264
rect 10008 4224 10014 4236
rect 10321 4233 10333 4236
rect 10367 4264 10379 4267
rect 10962 4264 10968 4276
rect 10367 4236 10968 4264
rect 10367 4233 10379 4236
rect 10321 4227 10379 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 11296 4236 11805 4264
rect 11296 4224 11302 4236
rect 11793 4233 11805 4236
rect 11839 4233 11851 4267
rect 11793 4227 11851 4233
rect 11900 4236 12388 4264
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 2556 4168 3403 4196
rect 2556 4156 2562 4168
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2130 4128 2136 4140
rect 1903 4100 2136 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2774 4128 2780 4140
rect 2455 4100 2780 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3375 4128 3403 4168
rect 3804 4168 4108 4196
rect 3375 4100 3556 4128
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3528 4069 3556 4100
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3694 4060 3700 4072
rect 3559 4032 3700 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3804 4069 3832 4168
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 4080 4128 4108 4168
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 4982 4196 4988 4208
rect 4212 4168 4988 4196
rect 4212 4156 4218 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 8754 4196 8760 4208
rect 5675 4168 8760 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 8849 4199 8907 4205
rect 8849 4165 8861 4199
rect 8895 4196 8907 4199
rect 10134 4196 10140 4208
rect 8895 4168 10140 4196
rect 8895 4165 8907 4168
rect 8849 4159 8907 4165
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 10597 4199 10655 4205
rect 10597 4165 10609 4199
rect 10643 4196 10655 4199
rect 10778 4196 10784 4208
rect 10643 4168 10784 4196
rect 10643 4165 10655 4168
rect 10597 4159 10655 4165
rect 4080 4100 6040 4128
rect 3973 4091 4031 4097
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4029 3847 4063
rect 3988 4060 4016 4091
rect 5644 4072 5672 4100
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 3988 4032 4721 4060
rect 3789 4023 3847 4029
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5350 4060 5356 4072
rect 4948 4032 5356 4060
rect 4948 4020 4954 4032
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5626 4020 5632 4072
rect 5684 4020 5690 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 4433 3995 4491 4001
rect 4433 3961 4445 3995
rect 4479 3992 4491 3995
rect 4614 3992 4620 4004
rect 4479 3964 4620 3992
rect 4479 3961 4491 3964
rect 4433 3955 4491 3961
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5736 3992 5764 4023
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 6012 4060 6040 4100
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 6144 4100 8125 4128
rect 6144 4088 6150 4100
rect 8113 4097 8125 4100
rect 8159 4128 8171 4131
rect 9306 4128 9312 4140
rect 8159 4100 9312 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 10612 4128 10640 4159
rect 10778 4156 10784 4168
rect 10836 4196 10842 4208
rect 11900 4196 11928 4236
rect 10836 4168 11928 4196
rect 10836 4156 10842 4168
rect 12158 4156 12164 4208
rect 12216 4196 12222 4208
rect 12360 4196 12388 4236
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 13081 4267 13139 4273
rect 13081 4264 13093 4267
rect 12768 4236 13093 4264
rect 12768 4224 12774 4236
rect 13081 4233 13093 4236
rect 13127 4233 13139 4267
rect 13081 4227 13139 4233
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 14918 4264 14924 4276
rect 13495 4236 14924 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 14918 4224 14924 4236
rect 14976 4224 14982 4276
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 15252 4236 15669 4264
rect 15252 4224 15258 4236
rect 15657 4233 15669 4236
rect 15703 4264 15715 4267
rect 16114 4264 16120 4276
rect 15703 4236 16120 4264
rect 15703 4233 15715 4236
rect 15657 4227 15715 4233
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 13170 4196 13176 4208
rect 12216 4168 12261 4196
rect 12360 4168 13176 4196
rect 12216 4156 12222 4168
rect 13170 4156 13176 4168
rect 13228 4156 13234 4208
rect 14458 4156 14464 4208
rect 14516 4196 14522 4208
rect 14553 4199 14611 4205
rect 14553 4196 14565 4199
rect 14516 4168 14565 4196
rect 14516 4156 14522 4168
rect 14553 4165 14565 4168
rect 14599 4165 14611 4199
rect 14553 4159 14611 4165
rect 9999 4100 10640 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10744 4100 10977 4128
rect 10744 4088 10750 4100
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 11974 4128 11980 4140
rect 11747 4100 11980 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12434 4128 12440 4140
rect 12299 4100 12440 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12434 4088 12440 4100
rect 12492 4128 12498 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12492 4100 12909 4128
rect 12492 4088 12498 4100
rect 12897 4097 12909 4100
rect 12943 4128 12955 4131
rect 13262 4128 13268 4140
rect 12943 4100 13268 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13722 4128 13728 4140
rect 13587 4100 13728 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 14568 4128 14596 4159
rect 14642 4156 14648 4208
rect 14700 4196 14706 4208
rect 15013 4199 15071 4205
rect 15013 4196 15025 4199
rect 14700 4168 15025 4196
rect 14700 4156 14706 4168
rect 15013 4165 15025 4168
rect 15059 4165 15071 4199
rect 15013 4159 15071 4165
rect 14826 4128 14832 4140
rect 14568 4100 14832 4128
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15470 4128 15476 4140
rect 15431 4100 15476 4128
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 8202 4060 8208 4072
rect 5868 4032 5913 4060
rect 6012 4032 8208 4060
rect 5868 4020 5874 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 9122 4060 9128 4072
rect 9083 4032 9128 4060
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 10042 4060 10048 4072
rect 10003 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 11848 4032 12357 4060
rect 11848 4020 11854 4032
rect 12345 4029 12357 4032
rect 12391 4029 12403 4063
rect 12345 4023 12403 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 7653 3995 7711 4001
rect 7653 3992 7665 3995
rect 4856 3964 5028 3992
rect 5736 3964 7665 3992
rect 4856 3952 4862 3964
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4154 3924 4160 3936
rect 4028 3896 4160 3924
rect 4028 3884 4034 3896
rect 4154 3884 4160 3896
rect 4212 3924 4218 3936
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4212 3896 4537 3924
rect 4212 3884 4218 3896
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4764 3896 4905 3924
rect 4764 3884 4770 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 5000 3924 5028 3964
rect 7653 3961 7665 3964
rect 7699 3961 7711 3995
rect 7653 3955 7711 3961
rect 9858 3952 9864 4004
rect 9916 3992 9922 4004
rect 10781 3995 10839 4001
rect 10781 3992 10793 3995
rect 9916 3964 10793 3992
rect 9916 3952 9922 3964
rect 10781 3961 10793 3964
rect 10827 3992 10839 3995
rect 10827 3964 11192 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 6178 3924 6184 3936
rect 5000 3896 6184 3924
rect 4893 3887 4951 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 11054 3924 11060 3936
rect 9456 3896 11060 3924
rect 9456 3884 9462 3896
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11164 3924 11192 3964
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 13648 3992 13676 4023
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14550 4060 14556 4072
rect 14424 4032 14556 4060
rect 14424 4020 14430 4032
rect 14550 4020 14556 4032
rect 14608 4060 14614 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14608 4032 14657 4060
rect 14608 4020 14614 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 11296 3964 13676 3992
rect 11296 3952 11302 3964
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14185 3995 14243 4001
rect 14185 3992 14197 3995
rect 13872 3964 14197 3992
rect 13872 3952 13878 3964
rect 14185 3961 14197 3964
rect 14231 3961 14243 3995
rect 14185 3955 14243 3961
rect 11330 3924 11336 3936
rect 11164 3896 11336 3924
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12158 3924 12164 3936
rect 11756 3896 12164 3924
rect 11756 3884 11762 3896
rect 12158 3884 12164 3896
rect 12216 3924 12222 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 12216 3896 12633 3924
rect 12216 3884 12222 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 12768 3896 13921 3924
rect 12768 3884 12774 3896
rect 13909 3893 13921 3896
rect 13955 3924 13967 3927
rect 14752 3924 14780 4023
rect 14826 3924 14832 3936
rect 13955 3896 14832 3924
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2556 3692 2697 3720
rect 2556 3680 2562 3692
rect 2685 3689 2697 3692
rect 2731 3720 2743 3723
rect 3418 3720 3424 3732
rect 2731 3692 3424 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 3970 3720 3976 3732
rect 3883 3692 3976 3720
rect 3970 3680 3976 3692
rect 4028 3720 4034 3732
rect 4798 3720 4804 3732
rect 4028 3692 4804 3720
rect 4028 3680 4034 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5074 3720 5080 3732
rect 4939 3692 5080 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5442 3720 5448 3732
rect 5307 3692 5448 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5442 3680 5448 3692
rect 5500 3720 5506 3732
rect 7006 3720 7012 3732
rect 5500 3692 7012 3720
rect 5500 3680 5506 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8812 3692 8953 3720
rect 8812 3680 8818 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9582 3720 9588 3732
rect 9364 3692 9588 3720
rect 9364 3680 9370 3692
rect 9582 3680 9588 3692
rect 9640 3720 9646 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9640 3692 9781 3720
rect 9640 3680 9646 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 9769 3683 9827 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11698 3720 11704 3732
rect 11020 3692 11704 3720
rect 11020 3680 11026 3692
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 12124 3692 12357 3720
rect 12124 3680 12130 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12710 3720 12716 3732
rect 12492 3692 12537 3720
rect 12671 3692 12716 3720
rect 12492 3680 12498 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 13262 3720 13268 3732
rect 12943 3692 13268 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 6181 3655 6239 3661
rect 6181 3652 6193 3655
rect 4580 3624 6193 3652
rect 4580 3612 4586 3624
rect 6181 3621 6193 3624
rect 6227 3621 6239 3655
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 6181 3615 6239 3621
rect 7392 3624 7849 3652
rect 4062 3584 4068 3596
rect 2148 3556 4068 3584
rect 2148 3525 2176 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 4396 3556 5917 3584
rect 4396 3544 4402 3556
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6512 3556 6745 3584
rect 6512 3544 6518 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2498 3516 2504 3528
rect 2459 3488 2504 3516
rect 2133 3479 2191 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 4356 3488 4752 3516
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 3237 3451 3295 3457
rect 3237 3448 3249 3451
rect 3108 3420 3249 3448
rect 3108 3408 3114 3420
rect 3237 3417 3249 3420
rect 3283 3448 3295 3451
rect 3283 3420 3648 3448
rect 3283 3417 3295 3420
rect 3237 3411 3295 3417
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2317 3383 2375 3389
rect 2317 3380 2329 3383
rect 2096 3352 2329 3380
rect 2096 3340 2102 3352
rect 2317 3349 2329 3352
rect 2363 3349 2375 3383
rect 2317 3343 2375 3349
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2556 3352 2881 3380
rect 2556 3340 2562 3352
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 3510 3380 3516 3392
rect 3471 3352 3516 3380
rect 2869 3343 2927 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 3620 3380 3648 3420
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 4356 3448 4384 3488
rect 3752 3420 4384 3448
rect 4433 3451 4491 3457
rect 3752 3408 3758 3420
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4724 3448 4752 3488
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 6362 3516 6368 3528
rect 5776 3488 6368 3516
rect 5776 3476 5782 3488
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 7392 3525 7420 3624
rect 7837 3621 7849 3624
rect 7883 3652 7895 3655
rect 9674 3652 9680 3664
rect 7883 3624 9680 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9950 3652 9956 3664
rect 9863 3624 9956 3652
rect 9950 3612 9956 3624
rect 10008 3652 10014 3664
rect 10870 3652 10876 3664
rect 10008 3624 10876 3652
rect 10008 3612 10014 3624
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 11054 3612 11060 3664
rect 11112 3652 11118 3664
rect 12912 3652 12940 3683
rect 13262 3680 13268 3692
rect 13320 3720 13326 3732
rect 13630 3720 13636 3732
rect 13320 3692 13636 3720
rect 13320 3680 13326 3692
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 13722 3680 13728 3732
rect 13780 3720 13786 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13780 3692 14105 3720
rect 13780 3680 13786 3692
rect 14093 3689 14105 3692
rect 14139 3720 14151 3723
rect 14458 3720 14464 3732
rect 14139 3692 14464 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 15470 3720 15476 3732
rect 14568 3692 15476 3720
rect 11112 3624 12940 3652
rect 13081 3655 13139 3661
rect 11112 3612 11118 3624
rect 13081 3621 13093 3655
rect 13127 3652 13139 3655
rect 14568 3652 14596 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 15746 3720 15752 3732
rect 15703 3692 15752 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 13127 3624 14596 3652
rect 14844 3624 15332 3652
rect 13127 3621 13139 3624
rect 13081 3615 13139 3621
rect 14844 3596 14872 3624
rect 7558 3584 7564 3596
rect 7519 3556 7564 3584
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8018 3584 8024 3596
rect 7668 3556 8024 3584
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 7668 3516 7696 3556
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 8260 3556 9505 3584
rect 8260 3544 8266 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10100 3556 10701 3584
rect 10100 3544 10106 3556
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 10689 3547 10747 3553
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11296 3556 11713 3584
rect 11296 3544 11302 3556
rect 11701 3553 11713 3556
rect 11747 3553 11759 3587
rect 11701 3547 11759 3553
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 13998 3584 14004 3596
rect 13771 3556 14004 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 13998 3544 14004 3556
rect 14056 3584 14062 3596
rect 14553 3587 14611 3593
rect 14056 3556 14320 3584
rect 14056 3544 14062 3556
rect 7515 3488 7696 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 7800 3488 10088 3516
rect 7800 3476 7806 3488
rect 10060 3460 10088 3488
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 11054 3516 11060 3528
rect 10284 3488 11060 3516
rect 10284 3476 10290 3488
rect 11054 3476 11060 3488
rect 11112 3476 11118 3528
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 12434 3516 12440 3528
rect 11563 3488 12440 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14292 3516 14320 3556
rect 14553 3553 14565 3587
rect 14599 3584 14611 3587
rect 14826 3584 14832 3596
rect 14599 3556 14832 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15194 3584 15200 3596
rect 15155 3556 15200 3584
rect 15194 3544 15200 3556
rect 15252 3544 15258 3596
rect 15304 3593 15332 3624
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15102 3516 15108 3528
rect 14292 3488 15108 3516
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 6822 3448 6828 3460
rect 4479 3420 4660 3448
rect 4724 3420 6828 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4062 3380 4068 3392
rect 3620 3352 4068 3380
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4212 3352 4537 3380
rect 4212 3340 4218 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 4632 3380 4660 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 8803 3420 9321 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 9401 3451 9459 3457
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 9582 3448 9588 3460
rect 9447 3420 9588 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 10042 3408 10048 3460
rect 10100 3408 10106 3460
rect 10505 3451 10563 3457
rect 10505 3417 10517 3451
rect 10551 3448 10563 3451
rect 10965 3451 11023 3457
rect 10965 3448 10977 3451
rect 10551 3420 10977 3448
rect 10551 3417 10563 3420
rect 10505 3411 10563 3417
rect 10965 3417 10977 3420
rect 11011 3417 11023 3451
rect 10965 3411 11023 3417
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 13633 3451 13691 3457
rect 11931 3420 13216 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 4890 3380 4896 3392
rect 4632 3352 4896 3380
rect 4525 3343 4583 3349
rect 4890 3340 4896 3352
rect 4948 3380 4954 3392
rect 4985 3383 5043 3389
rect 4985 3380 4997 3383
rect 4948 3352 4997 3380
rect 4948 3340 4954 3352
rect 4985 3349 4997 3352
rect 5031 3349 5043 3383
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 4985 3343 5043 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 6270 3380 6276 3392
rect 5859 3352 6276 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6546 3380 6552 3392
rect 6507 3352 6552 3380
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6641 3383 6699 3389
rect 6641 3349 6653 3383
rect 6687 3380 6699 3383
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6687 3352 7021 3380
rect 6687 3349 6699 3352
rect 6641 3343 6699 3349
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 9950 3380 9956 3392
rect 7984 3352 9956 3380
rect 7984 3340 7990 3352
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10597 3383 10655 3389
rect 10597 3349 10609 3383
rect 10643 3380 10655 3383
rect 10686 3380 10692 3392
rect 10643 3352 10692 3380
rect 10643 3349 10655 3352
rect 10597 3343 10655 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11330 3380 11336 3392
rect 11291 3352 11336 3380
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 13188 3389 13216 3420
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13679 3420 14780 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13173 3383 13231 3389
rect 12032 3352 12077 3380
rect 12032 3340 12038 3352
rect 13173 3349 13185 3383
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 14550 3380 14556 3392
rect 14415 3352 14556 3380
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14752 3389 14780 3420
rect 14737 3383 14795 3389
rect 14737 3349 14749 3383
rect 14783 3349 14795 3383
rect 14737 3343 14795 3349
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15746 3380 15752 3392
rect 15151 3352 15752 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 3418 3176 3424 3188
rect 2915 3148 3424 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5994 3176 6000 3188
rect 5399 3148 6000 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6178 3176 6184 3188
rect 6139 3148 6184 3176
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 6733 3179 6791 3185
rect 6733 3176 6745 3179
rect 6604 3148 6745 3176
rect 6604 3136 6610 3148
rect 6733 3145 6745 3148
rect 6779 3145 6791 3179
rect 6733 3139 6791 3145
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 6880 3148 8033 3176
rect 6880 3136 6886 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 9125 3179 9183 3185
rect 9125 3176 9137 3179
rect 8711 3148 9137 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 9125 3145 9137 3148
rect 9171 3145 9183 3179
rect 9125 3139 9183 3145
rect 9585 3179 9643 3185
rect 9585 3145 9597 3179
rect 9631 3176 9643 3179
rect 9950 3176 9956 3188
rect 9631 3148 9956 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 2317 3111 2375 3117
rect 2317 3077 2329 3111
rect 2363 3108 2375 3111
rect 2406 3108 2412 3120
rect 2363 3080 2412 3108
rect 2363 3077 2375 3080
rect 2317 3071 2375 3077
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 4522 3108 4528 3120
rect 3528 3080 4528 3108
rect 3528 3052 3556 3080
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4617 3111 4675 3117
rect 4617 3077 4629 3111
rect 4663 3108 4675 3111
rect 8312 3108 8340 3139
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10870 3176 10876 3188
rect 10831 3148 10876 3176
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11238 3176 11244 3188
rect 11199 3148 11244 3176
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11609 3179 11667 3185
rect 11609 3145 11621 3179
rect 11655 3145 11667 3179
rect 11974 3176 11980 3188
rect 11935 3148 11980 3176
rect 11609 3139 11667 3145
rect 11624 3108 11652 3139
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12805 3179 12863 3185
rect 12805 3176 12817 3179
rect 12483 3148 12817 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12805 3145 12817 3148
rect 12851 3145 12863 3179
rect 13262 3176 13268 3188
rect 13223 3148 13268 3176
rect 12805 3139 12863 3145
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14734 3176 14740 3188
rect 14292 3148 14740 3176
rect 12342 3108 12348 3120
rect 4663 3080 8340 3108
rect 8404 3080 11652 3108
rect 12303 3080 12348 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2222 3040 2228 3052
rect 2087 3012 2228 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2556 3012 2605 3040
rect 2556 3000 2562 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 3050 3040 3056 3052
rect 3011 3012 3056 3040
rect 2593 3003 2651 3009
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3040 3479 3043
rect 3510 3040 3516 3052
rect 3467 3012 3516 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3660 3012 3801 3040
rect 3660 3000 3666 3012
rect 3789 3009 3801 3012
rect 3835 3040 3847 3043
rect 3878 3040 3884 3052
rect 3835 3012 3884 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2608 2944 2774 2972
rect 2608 2916 2636 2944
rect 2590 2864 2596 2916
rect 2648 2864 2654 2916
rect 2746 2904 2774 2944
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3200 2944 4016 2972
rect 3200 2932 3206 2944
rect 3988 2913 4016 2944
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 2746 2876 3617 2904
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 3605 2867 3663 2873
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2873 4031 2907
rect 4172 2904 4200 3003
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 5445 3043 5503 3049
rect 4396 3012 5212 3040
rect 4396 3000 4402 3012
rect 4706 2972 4712 2984
rect 4667 2944 4712 2972
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 5074 2972 5080 2984
rect 4939 2944 5080 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5184 2981 5212 3012
rect 5445 3009 5457 3043
rect 5491 3040 5503 3043
rect 6178 3040 6184 3052
rect 5491 3012 6184 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 7098 3040 7104 3052
rect 7059 3012 7104 3040
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7239 3012 7849 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7837 3009 7849 3012
rect 7883 3040 7895 3043
rect 7926 3040 7932 3052
rect 7883 3012 7932 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8202 3040 8208 3052
rect 8163 3012 8208 3040
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2941 5227 2975
rect 6086 2972 6092 2984
rect 5169 2935 5227 2941
rect 5276 2944 6092 2972
rect 4246 2904 4252 2916
rect 4159 2876 4252 2904
rect 3973 2867 4031 2873
rect 4246 2864 4252 2876
rect 4304 2904 4310 2916
rect 5276 2904 5304 2944
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 7282 2972 7288 2984
rect 6972 2944 7288 2972
rect 6972 2932 6978 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7374 2932 7380 2984
rect 7432 2972 7438 2984
rect 7432 2944 7477 2972
rect 7432 2932 7438 2944
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 8404 2972 8432 3080
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 13078 3068 13084 3120
rect 13136 3108 13142 3120
rect 13173 3111 13231 3117
rect 13173 3108 13185 3111
rect 13136 3080 13185 3108
rect 13136 3068 13142 3080
rect 13173 3077 13185 3080
rect 13219 3108 13231 3111
rect 14292 3108 14320 3148
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 13219 3080 14320 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 14458 3068 14464 3120
rect 14516 3108 14522 3120
rect 15013 3111 15071 3117
rect 15013 3108 15025 3111
rect 14516 3080 15025 3108
rect 14516 3068 14522 3080
rect 15013 3077 15025 3080
rect 15059 3077 15071 3111
rect 15013 3071 15071 3077
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 9490 3040 9496 3052
rect 8536 3012 8892 3040
rect 9451 3012 9496 3040
rect 8536 3000 8542 3012
rect 8864 2981 8892 3012
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 10226 3040 10232 3052
rect 10139 3012 10232 3040
rect 10226 3000 10232 3012
rect 10284 3040 10290 3052
rect 10686 3040 10692 3052
rect 10284 3012 10692 3040
rect 10284 3000 10290 3012
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11238 3040 11244 3052
rect 10827 3012 11244 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 12434 3040 12440 3052
rect 11793 3003 11851 3009
rect 7616 2944 8432 2972
rect 8757 2975 8815 2981
rect 7616 2932 7622 2944
rect 8757 2941 8769 2975
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 4304 2876 5304 2904
rect 4304 2864 4310 2876
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 7653 2907 7711 2913
rect 7653 2904 7665 2907
rect 5684 2876 7665 2904
rect 5684 2864 5690 2876
rect 7653 2873 7665 2876
rect 7699 2873 7711 2907
rect 8772 2904 8800 2935
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 9732 2944 9781 2972
rect 9732 2932 9738 2944
rect 9769 2941 9781 2944
rect 9815 2972 9827 2975
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 9815 2944 10977 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 10965 2941 10977 2944
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11808 2972 11836 3003
rect 12406 3000 12440 3040
rect 12492 3000 12498 3052
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 13633 3043 13691 3049
rect 13633 3040 13645 3043
rect 13504 3012 13645 3040
rect 13504 3000 13510 3012
rect 13633 3009 13645 3012
rect 13679 3009 13691 3043
rect 14182 3040 14188 3052
rect 14143 3012 14188 3040
rect 13633 3003 13691 3009
rect 14182 3000 14188 3012
rect 14240 3040 14246 3052
rect 14550 3040 14556 3052
rect 14240 3012 14556 3040
rect 14240 3000 14246 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 15470 3040 15476 3052
rect 14783 3012 15476 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 12406 2972 12434 3000
rect 11112 2944 11744 2972
rect 11808 2944 12434 2972
rect 12621 2975 12679 2981
rect 11112 2932 11118 2944
rect 10413 2907 10471 2913
rect 10413 2904 10425 2907
rect 7653 2867 7711 2873
rect 7760 2876 8156 2904
rect 8772 2876 10425 2904
rect 3234 2836 3240 2848
rect 3195 2808 3240 2836
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 5442 2836 5448 2848
rect 4120 2808 5448 2836
rect 4120 2796 4126 2808
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 7760 2836 7788 2876
rect 6512 2808 7788 2836
rect 8128 2836 8156 2876
rect 10413 2873 10425 2876
rect 10459 2873 10471 2907
rect 11514 2904 11520 2916
rect 10413 2867 10471 2873
rect 11072 2876 11520 2904
rect 10045 2839 10103 2845
rect 10045 2836 10057 2839
rect 8128 2808 10057 2836
rect 6512 2796 6518 2808
rect 10045 2805 10057 2808
rect 10091 2805 10103 2839
rect 10045 2799 10103 2805
rect 10686 2796 10692 2848
rect 10744 2836 10750 2848
rect 11072 2836 11100 2876
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 11716 2904 11744 2944
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 12342 2904 12348 2916
rect 11716 2876 12348 2904
rect 12342 2864 12348 2876
rect 12400 2864 12406 2916
rect 12636 2904 12664 2935
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12768 2944 13369 2972
rect 12768 2932 12774 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13906 2972 13912 2984
rect 13867 2944 13912 2972
rect 13357 2935 13415 2941
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 14507 2944 14780 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 14752 2916 14780 2944
rect 13998 2904 14004 2916
rect 12636 2876 14004 2904
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 14734 2864 14740 2916
rect 14792 2864 14798 2916
rect 10744 2808 11100 2836
rect 10744 2796 10750 2808
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14844 2836 14872 3012
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 15654 3040 15660 3052
rect 15611 3012 15660 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15378 2904 15384 2916
rect 15339 2876 15384 2904
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 13780 2808 14872 2836
rect 13780 2796 13786 2808
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 3878 2632 3884 2644
rect 3384 2604 3884 2632
rect 3384 2592 3390 2604
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 4246 2632 4252 2644
rect 4019 2604 4252 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4764 2604 4813 2632
rect 4764 2592 4770 2604
rect 4801 2601 4813 2604
rect 4847 2601 4859 2635
rect 4801 2595 4859 2601
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 10689 2635 10747 2641
rect 5040 2604 5856 2632
rect 5040 2592 5046 2604
rect 1854 2524 1860 2576
rect 1912 2564 1918 2576
rect 2685 2567 2743 2573
rect 2685 2564 2697 2567
rect 1912 2536 2697 2564
rect 1912 2524 1918 2536
rect 2685 2533 2697 2536
rect 2731 2533 2743 2567
rect 2685 2527 2743 2533
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 3237 2567 3295 2573
rect 3237 2564 3249 2567
rect 2924 2536 3249 2564
rect 2924 2524 2930 2536
rect 3237 2533 3249 2536
rect 3283 2533 3295 2567
rect 5718 2564 5724 2576
rect 3237 2527 3295 2533
rect 4172 2536 5724 2564
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 4172 2496 4200 2536
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 2179 2468 4200 2496
rect 4249 2499 4307 2505
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 1995 2400 2513 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2516 2360 2544 2391
rect 2682 2388 2688 2440
rect 2740 2428 2746 2440
rect 2884 2437 2912 2468
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 5258 2496 5264 2508
rect 4295 2468 5264 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5408 2468 5549 2496
rect 5408 2456 5414 2468
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 5828 2496 5856 2604
rect 6886 2604 10364 2632
rect 5902 2524 5908 2576
rect 5960 2564 5966 2576
rect 6886 2564 6914 2604
rect 7653 2567 7711 2573
rect 5960 2536 6914 2564
rect 7015 2536 7328 2564
rect 5960 2524 5966 2536
rect 5675 2468 5948 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2740 2400 2881 2428
rect 2740 2388 2746 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 3099 2400 3433 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3421 2397 3433 2400
rect 3467 2428 3479 2431
rect 4062 2428 4068 2440
rect 3467 2400 4068 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4430 2428 4436 2440
rect 4391 2400 4436 2428
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 3326 2360 3332 2372
rect 2516 2332 3332 2360
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 4341 2363 4399 2369
rect 4341 2329 4353 2363
rect 4387 2360 4399 2363
rect 4387 2332 5120 2360
rect 4387 2329 4399 2332
rect 4341 2323 4399 2329
rect 2314 2292 2320 2304
rect 2275 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 3602 2292 3608 2304
rect 3563 2264 3608 2292
rect 3602 2252 3608 2264
rect 3660 2252 3666 2304
rect 5092 2301 5120 2332
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2261 5135 2295
rect 5276 2292 5304 2456
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5810 2428 5816 2440
rect 5491 2400 5816 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 5920 2428 5948 2468
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 7015 2496 7043 2536
rect 6052 2468 7043 2496
rect 6052 2456 6058 2468
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 7156 2468 7205 2496
rect 7156 2456 7162 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7300 2496 7328 2536
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 8018 2564 8024 2576
rect 7699 2536 8024 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9732 2536 10241 2564
rect 9732 2524 9738 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10336 2564 10364 2604
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 10778 2632 10784 2644
rect 10735 2604 10784 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11514 2632 11520 2644
rect 11475 2604 11520 2632
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 12342 2592 12348 2644
rect 12400 2632 12406 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 12400 2604 12449 2632
rect 12400 2592 12406 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 12437 2595 12495 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13081 2635 13139 2641
rect 13081 2601 13093 2635
rect 13127 2632 13139 2635
rect 13262 2632 13268 2644
rect 13127 2604 13268 2632
rect 13127 2601 13139 2604
rect 13081 2595 13139 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13722 2632 13728 2644
rect 13412 2604 13728 2632
rect 13412 2592 13418 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 15286 2564 15292 2576
rect 10336 2536 15292 2564
rect 10229 2527 10287 2533
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 8478 2496 8484 2508
rect 7300 2468 8484 2496
rect 7193 2459 7251 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8757 2499 8815 2505
rect 8757 2465 8769 2499
rect 8803 2496 8815 2499
rect 8803 2468 9260 2496
rect 8803 2465 8815 2468
rect 8757 2459 8815 2465
rect 9030 2428 9036 2440
rect 5920 2400 9036 2428
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9232 2437 9260 2468
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9548 2468 9597 2496
rect 9548 2456 9554 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 10778 2496 10784 2508
rect 9585 2459 9643 2465
rect 10152 2468 10784 2496
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9306 2428 9312 2440
rect 9263 2400 9312 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 10152 2437 10180 2468
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 12618 2496 12624 2508
rect 11379 2468 12624 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 10137 2431 10195 2437
rect 10137 2397 10149 2431
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11992 2437 12020 2468
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13357 2499 13415 2505
rect 13357 2465 13369 2499
rect 13403 2496 13415 2499
rect 13630 2496 13636 2508
rect 13403 2468 13636 2496
rect 13403 2465 13415 2468
rect 13357 2459 13415 2465
rect 13630 2456 13636 2468
rect 13688 2496 13694 2508
rect 16022 2496 16028 2508
rect 13688 2468 16028 2496
rect 13688 2456 13694 2468
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10284 2400 10425 2428
rect 10284 2388 10290 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 13262 2428 13268 2440
rect 12391 2400 13268 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14660 2437 14688 2468
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 13872 2400 13921 2428
rect 13872 2388 13878 2400
rect 13909 2397 13921 2400
rect 13955 2428 13967 2431
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 13955 2400 14381 2428
rect 13955 2397 13967 2400
rect 13909 2391 13967 2397
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 15194 2428 15200 2440
rect 15107 2400 15200 2428
rect 14645 2391 14703 2397
rect 15194 2388 15200 2400
rect 15252 2428 15258 2440
rect 15838 2428 15844 2440
rect 15252 2400 15844 2428
rect 15252 2388 15258 2400
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 5350 2320 5356 2372
rect 5408 2360 5414 2372
rect 5408 2332 6914 2360
rect 5408 2320 5414 2332
rect 5994 2292 6000 2304
rect 5276 2264 6000 2292
rect 5077 2255 5135 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 6886 2292 6914 2332
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 8297 2363 8355 2369
rect 8297 2360 8309 2363
rect 8260 2332 8309 2360
rect 8260 2320 8266 2332
rect 8297 2329 8309 2332
rect 8343 2360 8355 2363
rect 8343 2332 12388 2360
rect 8343 2329 8355 2332
rect 8297 2323 8355 2329
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 6886 2264 9045 2292
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9180 2264 9321 2292
rect 9180 2252 9186 2264
rect 9309 2261 9321 2264
rect 9355 2292 9367 2295
rect 9674 2292 9680 2304
rect 9355 2264 9680 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11238 2292 11244 2304
rect 11195 2264 11244 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11790 2292 11796 2304
rect 11751 2264 11796 2292
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 11940 2264 12173 2292
rect 11940 2252 11946 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12360 2292 12388 2332
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12713 2363 12771 2369
rect 12713 2360 12725 2363
rect 12492 2332 12725 2360
rect 12492 2320 12498 2332
rect 12713 2329 12725 2332
rect 12759 2360 12771 2363
rect 14550 2360 14556 2372
rect 12759 2332 14556 2360
rect 12759 2329 12771 2332
rect 12713 2323 12771 2329
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 14921 2363 14979 2369
rect 14921 2329 14933 2363
rect 14967 2360 14979 2363
rect 15010 2360 15016 2372
rect 14967 2332 15016 2360
rect 14967 2329 14979 2332
rect 14921 2323 14979 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 15286 2320 15292 2372
rect 15344 2360 15350 2372
rect 15473 2363 15531 2369
rect 15473 2360 15485 2363
rect 15344 2332 15485 2360
rect 15344 2320 15350 2332
rect 15473 2329 15485 2332
rect 15519 2329 15531 2363
rect 15473 2323 15531 2329
rect 12894 2292 12900 2304
rect 12360 2264 12900 2292
rect 12161 2255 12219 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 13446 2292 13452 2304
rect 13407 2264 13452 2292
rect 13446 2252 13452 2264
rect 13504 2252 13510 2304
rect 14182 2292 14188 2304
rect 14143 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 5074 2048 5080 2100
rect 5132 2088 5138 2100
rect 11790 2088 11796 2100
rect 5132 2060 11796 2088
rect 5132 2048 5138 2060
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
rect 4522 1980 4528 2032
rect 4580 2020 4586 2032
rect 9950 2020 9956 2032
rect 4580 1992 9956 2020
rect 4580 1980 4586 1992
rect 9950 1980 9956 1992
rect 10008 1980 10014 2032
rect 6454 1912 6460 1964
rect 6512 1952 6518 1964
rect 11882 1952 11888 1964
rect 6512 1924 11888 1952
rect 6512 1912 6518 1924
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 3602 1844 3608 1896
rect 3660 1884 3666 1896
rect 9858 1884 9864 1896
rect 3660 1856 9864 1884
rect 3660 1844 3666 1856
rect 9858 1844 9864 1856
rect 9916 1844 9922 1896
rect 2498 1776 2504 1828
rect 2556 1816 2562 1828
rect 13078 1816 13084 1828
rect 2556 1788 13084 1816
rect 2556 1776 2562 1788
rect 13078 1776 13084 1788
rect 13136 1816 13142 1828
rect 13446 1816 13452 1828
rect 13136 1788 13452 1816
rect 13136 1776 13142 1788
rect 13446 1776 13452 1788
rect 13504 1776 13510 1828
rect 2130 1640 2136 1692
rect 2188 1680 2194 1692
rect 11606 1680 11612 1692
rect 2188 1652 11612 1680
rect 2188 1640 2194 1652
rect 11606 1640 11612 1652
rect 11664 1640 11670 1692
rect 11238 1436 11244 1488
rect 11296 1476 11302 1488
rect 13906 1476 13912 1488
rect 11296 1448 13912 1476
rect 11296 1436 11302 1448
rect 13906 1436 13912 1448
rect 13964 1476 13970 1488
rect 15194 1476 15200 1488
rect 13964 1448 15200 1476
rect 13964 1436 13970 1448
rect 15194 1436 15200 1448
rect 15252 1436 15258 1488
rect 6086 1368 6092 1420
rect 6144 1408 6150 1420
rect 7834 1408 7840 1420
rect 6144 1380 7840 1408
rect 6144 1368 6150 1380
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
<< via1 >>
rect 664 17484 716 17536
rect 12072 17484 12124 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 2504 17280 2556 17332
rect 3608 17280 3660 17332
rect 4344 17323 4396 17332
rect 4344 17289 4353 17323
rect 4353 17289 4387 17323
rect 4387 17289 4396 17323
rect 4344 17280 4396 17289
rect 7656 17280 7708 17332
rect 8852 17280 8904 17332
rect 11980 17280 12032 17332
rect 16488 17280 16540 17332
rect 1400 17212 1452 17264
rect 2596 17212 2648 17264
rect 2780 17144 2832 17196
rect 3148 17144 3200 17196
rect 3332 17144 3384 17196
rect 12072 17212 12124 17264
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4252 17076 4304 17128
rect 6368 17076 6420 17128
rect 10048 17076 10100 17128
rect 15568 17144 15620 17196
rect 12624 17076 12676 17128
rect 13360 17076 13412 17128
rect 16120 17076 16172 17128
rect 2872 17008 2924 17060
rect 7012 17008 7064 17060
rect 7932 17008 7984 17060
rect 10968 17008 11020 17060
rect 13636 17008 13688 17060
rect 14556 17008 14608 17060
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 3148 16983 3200 16992
rect 3148 16949 3157 16983
rect 3157 16949 3191 16983
rect 3191 16949 3200 16983
rect 3148 16940 3200 16949
rect 3792 16940 3844 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 9864 16940 9916 16992
rect 10600 16940 10652 16992
rect 12624 16983 12676 16992
rect 12624 16949 12633 16983
rect 12633 16949 12667 16983
rect 12667 16949 12676 16983
rect 12624 16940 12676 16949
rect 14740 16940 14792 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 8392 16736 8444 16788
rect 9404 16736 9456 16788
rect 9588 16736 9640 16788
rect 6736 16711 6788 16720
rect 6736 16677 6745 16711
rect 6745 16677 6779 16711
rect 6779 16677 6788 16711
rect 6736 16668 6788 16677
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 2044 16532 2096 16584
rect 2596 16532 2648 16584
rect 5724 16643 5776 16652
rect 5724 16609 5733 16643
rect 5733 16609 5767 16643
rect 5767 16609 5776 16643
rect 5724 16600 5776 16609
rect 3608 16575 3660 16584
rect 2136 16507 2188 16516
rect 2136 16473 2145 16507
rect 2145 16473 2179 16507
rect 2179 16473 2188 16507
rect 2136 16464 2188 16473
rect 2228 16464 2280 16516
rect 2780 16464 2832 16516
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 3240 16396 3292 16448
rect 3700 16396 3752 16448
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 5264 16532 5316 16584
rect 5540 16532 5592 16584
rect 6368 16532 6420 16584
rect 7012 16600 7064 16652
rect 8392 16600 8444 16652
rect 9036 16600 9088 16652
rect 9404 16600 9456 16652
rect 4068 16464 4120 16516
rect 9588 16532 9640 16584
rect 13176 16736 13228 16788
rect 12716 16668 12768 16720
rect 10784 16532 10836 16584
rect 12072 16600 12124 16652
rect 12992 16600 13044 16652
rect 13360 16668 13412 16720
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 12900 16532 12952 16584
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 4344 16396 4396 16448
rect 5080 16396 5132 16448
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 6460 16396 6512 16448
rect 7288 16439 7340 16448
rect 7288 16405 7297 16439
rect 7297 16405 7331 16439
rect 7331 16405 7340 16439
rect 7288 16396 7340 16405
rect 7380 16439 7432 16448
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 9128 16464 9180 16516
rect 7380 16396 7432 16405
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 9864 16396 9916 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 10600 16439 10652 16448
rect 10600 16405 10609 16439
rect 10609 16405 10643 16439
rect 10643 16405 10652 16439
rect 10600 16396 10652 16405
rect 13360 16396 13412 16448
rect 14740 16396 14792 16448
rect 15844 16396 15896 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 4528 16192 4580 16244
rect 5448 16192 5500 16244
rect 6184 16192 6236 16244
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 7288 16192 7340 16244
rect 8024 16192 8076 16244
rect 9680 16192 9732 16244
rect 9956 16192 10008 16244
rect 3148 16167 3200 16176
rect 3148 16133 3182 16167
rect 3182 16133 3200 16167
rect 3148 16124 3200 16133
rect 3608 16124 3660 16176
rect 7380 16124 7432 16176
rect 7748 16124 7800 16176
rect 8392 16124 8444 16176
rect 10140 16192 10192 16244
rect 11980 16235 12032 16244
rect 11980 16201 11989 16235
rect 11989 16201 12023 16235
rect 12023 16201 12032 16235
rect 11980 16192 12032 16201
rect 12440 16192 12492 16244
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 15752 16192 15804 16244
rect 12256 16124 12308 16176
rect 14464 16124 14516 16176
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2688 16056 2740 16108
rect 2504 15988 2556 16040
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 4988 16056 5040 16108
rect 6460 16056 6512 16108
rect 7196 16056 7248 16108
rect 8116 16056 8168 16108
rect 6092 15988 6144 16040
rect 7840 15988 7892 16040
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 9680 16056 9732 16108
rect 4436 15920 4488 15972
rect 4620 15920 4672 15972
rect 5080 15920 5132 15972
rect 5816 15920 5868 15972
rect 4344 15895 4396 15904
rect 4344 15861 4353 15895
rect 4353 15861 4387 15895
rect 4387 15861 4396 15895
rect 4344 15852 4396 15861
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 6184 15852 6236 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 8116 15920 8168 15972
rect 9312 15988 9364 16040
rect 10324 16056 10376 16108
rect 11704 16056 11756 16108
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12164 16056 12216 16108
rect 13636 16099 13688 16108
rect 9496 15920 9548 15972
rect 8300 15852 8352 15904
rect 8392 15852 8444 15904
rect 9680 15852 9732 15904
rect 9772 15852 9824 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11520 15988 11572 16040
rect 12348 15988 12400 16040
rect 13636 16065 13645 16099
rect 13645 16065 13679 16099
rect 13679 16065 13688 16099
rect 13636 16056 13688 16065
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 11980 15920 12032 15972
rect 16028 15920 16080 15972
rect 11520 15852 11572 15904
rect 11796 15852 11848 15904
rect 12532 15852 12584 15904
rect 15936 15852 15988 15904
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 2320 15648 2372 15700
rect 2780 15648 2832 15700
rect 2044 15512 2096 15564
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 2504 15444 2556 15496
rect 6184 15648 6236 15700
rect 6920 15648 6972 15700
rect 10692 15648 10744 15700
rect 12256 15691 12308 15700
rect 12256 15657 12265 15691
rect 12265 15657 12299 15691
rect 12299 15657 12308 15691
rect 12256 15648 12308 15657
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12716 15691 12768 15700
rect 12440 15648 12492 15657
rect 12716 15657 12725 15691
rect 12725 15657 12759 15691
rect 12759 15657 12768 15691
rect 12716 15648 12768 15657
rect 13820 15648 13872 15700
rect 14464 15648 14516 15700
rect 11704 15580 11756 15632
rect 14832 15580 14884 15632
rect 1400 15376 1452 15428
rect 2780 15376 2832 15428
rect 4160 15512 4212 15564
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 12992 15512 13044 15564
rect 13636 15512 13688 15564
rect 4344 15444 4396 15496
rect 5540 15444 5592 15496
rect 6184 15444 6236 15496
rect 7196 15444 7248 15496
rect 8208 15444 8260 15496
rect 11336 15444 11388 15496
rect 12164 15444 12216 15496
rect 13360 15444 13412 15496
rect 4160 15376 4212 15428
rect 8300 15376 8352 15428
rect 9496 15376 9548 15428
rect 13912 15376 13964 15428
rect 296 15308 348 15360
rect 2320 15308 2372 15360
rect 2504 15351 2556 15360
rect 2504 15317 2513 15351
rect 2513 15317 2547 15351
rect 2547 15317 2556 15351
rect 2504 15308 2556 15317
rect 2688 15308 2740 15360
rect 4068 15308 4120 15360
rect 5172 15308 5224 15360
rect 5816 15308 5868 15360
rect 6000 15308 6052 15360
rect 7472 15308 7524 15360
rect 10968 15308 11020 15360
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 1952 15104 2004 15156
rect 2596 15104 2648 15156
rect 4344 15147 4396 15156
rect 2412 15079 2464 15088
rect 2412 15045 2421 15079
rect 2421 15045 2455 15079
rect 2455 15045 2464 15079
rect 2412 15036 2464 15045
rect 2504 14968 2556 15020
rect 4068 15036 4120 15088
rect 3608 14968 3660 15020
rect 1584 14943 1636 14952
rect 1584 14909 1593 14943
rect 1593 14909 1627 14943
rect 1627 14909 1636 14943
rect 1584 14900 1636 14909
rect 4344 15113 4353 15147
rect 4353 15113 4387 15147
rect 4387 15113 4396 15147
rect 4344 15104 4396 15113
rect 13544 15104 13596 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 16856 15104 16908 15156
rect 6000 15036 6052 15088
rect 5356 14968 5408 15020
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 7196 14968 7248 15020
rect 7472 15036 7524 15088
rect 10324 15036 10376 15088
rect 11796 15079 11848 15088
rect 2688 14832 2740 14884
rect 2136 14807 2188 14816
rect 2136 14773 2145 14807
rect 2145 14773 2179 14807
rect 2179 14773 2188 14807
rect 2136 14764 2188 14773
rect 3148 14764 3200 14816
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 8208 14968 8260 15020
rect 10692 15011 10744 15020
rect 10692 14977 10710 15011
rect 10710 14977 10744 15011
rect 10692 14968 10744 14977
rect 10876 14968 10928 15020
rect 11796 15045 11805 15079
rect 11805 15045 11839 15079
rect 11839 15045 11848 15079
rect 11796 15036 11848 15045
rect 11980 15036 12032 15088
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 13452 15036 13504 15088
rect 13636 15036 13688 15088
rect 14648 14968 14700 15020
rect 9312 14764 9364 14816
rect 11888 14900 11940 14952
rect 13084 14900 13136 14952
rect 10968 14832 11020 14884
rect 16304 14900 16356 14952
rect 12624 14764 12676 14816
rect 12716 14764 12768 14816
rect 13820 14764 13872 14816
rect 15016 14764 15068 14816
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 2872 14560 2924 14612
rect 4068 14560 4120 14612
rect 4344 14560 4396 14612
rect 5448 14560 5500 14612
rect 9312 14560 9364 14612
rect 9496 14560 9548 14612
rect 13084 14603 13136 14612
rect 1952 14356 2004 14408
rect 2872 14356 2924 14408
rect 8944 14424 8996 14476
rect 11888 14467 11940 14476
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 1768 14288 1820 14340
rect 2688 14288 2740 14340
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 4160 14220 4212 14272
rect 5356 14220 5408 14272
rect 5816 14220 5868 14272
rect 7104 14356 7156 14408
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 13268 14560 13320 14612
rect 12900 14492 12952 14544
rect 13452 14492 13504 14544
rect 15200 14424 15252 14476
rect 7932 14288 7984 14340
rect 8208 14288 8260 14340
rect 15660 14356 15712 14408
rect 9588 14288 9640 14340
rect 11888 14288 11940 14340
rect 13820 14288 13872 14340
rect 9864 14220 9916 14272
rect 10692 14220 10744 14272
rect 12072 14263 12124 14272
rect 12072 14229 12081 14263
rect 12081 14229 12115 14263
rect 12115 14229 12124 14263
rect 12072 14220 12124 14229
rect 12808 14220 12860 14272
rect 13268 14220 13320 14272
rect 14556 14263 14608 14272
rect 14556 14229 14565 14263
rect 14565 14229 14599 14263
rect 14599 14229 14608 14263
rect 14556 14220 14608 14229
rect 15476 14288 15528 14340
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 4252 14016 4304 14068
rect 5080 14016 5132 14068
rect 9128 14016 9180 14068
rect 9404 14016 9456 14068
rect 9496 14016 9548 14068
rect 11612 14016 11664 14068
rect 12256 14016 12308 14068
rect 12808 14059 12860 14068
rect 2872 13948 2924 14000
rect 3516 13948 3568 14000
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 13268 14016 13320 14068
rect 13636 14059 13688 14068
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 13912 14016 13964 14068
rect 15016 14016 15068 14068
rect 15752 14016 15804 14068
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 4068 13880 4120 13932
rect 5908 13880 5960 13932
rect 6828 13880 6880 13932
rect 7380 13880 7432 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 12624 13948 12676 14000
rect 13084 13948 13136 14000
rect 14648 13948 14700 14000
rect 8852 13880 8904 13932
rect 9312 13880 9364 13932
rect 11152 13880 11204 13932
rect 12532 13880 12584 13932
rect 11060 13812 11112 13864
rect 13452 13880 13504 13932
rect 13912 13880 13964 13932
rect 14464 13880 14516 13932
rect 3516 13676 3568 13728
rect 6184 13744 6236 13796
rect 9772 13744 9824 13796
rect 4436 13676 4488 13728
rect 6276 13676 6328 13728
rect 11520 13719 11572 13728
rect 11520 13685 11529 13719
rect 11529 13685 11563 13719
rect 11563 13685 11572 13719
rect 11520 13676 11572 13685
rect 11796 13744 11848 13796
rect 13728 13676 13780 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 4160 13472 4212 13524
rect 5264 13472 5316 13524
rect 7196 13515 7248 13524
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7564 13472 7616 13524
rect 11888 13515 11940 13524
rect 8944 13404 8996 13456
rect 11060 13447 11112 13456
rect 11060 13413 11069 13447
rect 11069 13413 11103 13447
rect 11103 13413 11112 13447
rect 11060 13404 11112 13413
rect 1584 13336 1636 13388
rect 2596 13336 2648 13388
rect 4068 13336 4120 13388
rect 4252 13336 4304 13388
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 11980 13472 12032 13524
rect 13360 13472 13412 13524
rect 13636 13472 13688 13524
rect 14556 13472 14608 13524
rect 11336 13336 11388 13388
rect 11520 13336 11572 13388
rect 13360 13336 13412 13388
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 14740 13336 14792 13388
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 15292 13336 15344 13388
rect 2688 13268 2740 13320
rect 3700 13268 3752 13320
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 4528 13200 4580 13252
rect 5908 13268 5960 13320
rect 7288 13268 7340 13320
rect 7932 13268 7984 13320
rect 7104 13200 7156 13252
rect 4436 13132 4488 13184
rect 8852 13200 8904 13252
rect 9864 13268 9916 13320
rect 10876 13268 10928 13320
rect 12900 13268 12952 13320
rect 14004 13268 14056 13320
rect 15384 13268 15436 13320
rect 10048 13200 10100 13252
rect 11428 13200 11480 13252
rect 11704 13200 11756 13252
rect 11060 13132 11112 13184
rect 11612 13132 11664 13184
rect 11796 13132 11848 13184
rect 11980 13132 12032 13184
rect 12256 13132 12308 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 13912 13132 13964 13184
rect 14832 13132 14884 13184
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 4068 12928 4120 12980
rect 4252 12928 4304 12980
rect 4804 12928 4856 12980
rect 5908 12928 5960 12980
rect 10140 12928 10192 12980
rect 11428 12928 11480 12980
rect 11704 12928 11756 12980
rect 13544 12928 13596 12980
rect 13820 12928 13872 12980
rect 15200 12928 15252 12980
rect 15384 12928 15436 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 4160 12792 4212 12844
rect 4712 12792 4764 12844
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 5080 12835 5132 12844
rect 4804 12792 4856 12801
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 6092 12792 6144 12844
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 5172 12724 5224 12776
rect 6276 12724 6328 12776
rect 8852 12860 8904 12912
rect 6828 12835 6880 12844
rect 6828 12801 6862 12835
rect 6862 12801 6880 12835
rect 6828 12792 6880 12801
rect 10140 12792 10192 12844
rect 11244 12792 11296 12844
rect 5908 12656 5960 12708
rect 6460 12656 6512 12708
rect 4160 12588 4212 12640
rect 4896 12588 4948 12640
rect 7932 12724 7984 12776
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 11152 12724 11204 12776
rect 7656 12656 7708 12708
rect 13360 12792 13412 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 13544 12724 13596 12776
rect 14740 12860 14792 12912
rect 15016 12792 15068 12844
rect 14740 12767 14792 12776
rect 8760 12588 8812 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 14740 12733 14749 12767
rect 14749 12733 14783 12767
rect 14783 12733 14792 12767
rect 14740 12724 14792 12733
rect 15292 12724 15344 12776
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 12256 12588 12308 12597
rect 14004 12588 14056 12640
rect 15016 12588 15068 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 1400 12384 1452 12436
rect 3332 12316 3384 12368
rect 4252 12384 4304 12436
rect 5632 12384 5684 12436
rect 10784 12384 10836 12436
rect 12072 12384 12124 12436
rect 13912 12384 13964 12436
rect 14096 12384 14148 12436
rect 14832 12384 14884 12436
rect 14924 12384 14976 12436
rect 11152 12316 11204 12368
rect 14188 12316 14240 12368
rect 2228 12248 2280 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 3700 12180 3752 12232
rect 4896 12223 4948 12232
rect 4896 12189 4914 12223
rect 4914 12189 4948 12223
rect 4896 12180 4948 12189
rect 6000 12180 6052 12232
rect 6552 12180 6604 12232
rect 9312 12248 9364 12300
rect 10876 12248 10928 12300
rect 11336 12248 11388 12300
rect 12256 12248 12308 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 8944 12180 8996 12232
rect 9404 12180 9456 12232
rect 4068 12112 4120 12164
rect 5080 12112 5132 12164
rect 6920 12112 6972 12164
rect 8116 12112 8168 12164
rect 9036 12112 9088 12164
rect 9956 12112 10008 12164
rect 12992 12180 13044 12232
rect 13912 12180 13964 12232
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 11796 12112 11848 12164
rect 12256 12112 12308 12164
rect 14096 12112 14148 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 3608 12044 3660 12096
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 6460 12044 6512 12096
rect 9680 12044 9732 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 12992 12044 13044 12096
rect 13636 12044 13688 12096
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 1952 11840 2004 11892
rect 2136 11840 2188 11892
rect 2228 11840 2280 11892
rect 7472 11840 7524 11892
rect 7564 11840 7616 11892
rect 4252 11772 4304 11824
rect 4436 11772 4488 11824
rect 5448 11772 5500 11824
rect 6552 11815 6604 11824
rect 6552 11781 6561 11815
rect 6561 11781 6595 11815
rect 6595 11781 6604 11815
rect 6552 11772 6604 11781
rect 2320 11704 2372 11756
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 2596 11636 2648 11688
rect 4896 11704 4948 11756
rect 7564 11704 7616 11756
rect 10232 11772 10284 11824
rect 10968 11772 11020 11824
rect 8484 11704 8536 11756
rect 11152 11704 11204 11756
rect 11520 11704 11572 11756
rect 9496 11636 9548 11688
rect 9680 11636 9732 11688
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 12072 11840 12124 11892
rect 13176 11840 13228 11892
rect 13636 11840 13688 11892
rect 13820 11772 13872 11824
rect 13636 11704 13688 11756
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14556 11704 14608 11756
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5448 11500 5500 11552
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 6460 11500 6512 11552
rect 8116 11568 8168 11620
rect 11520 11568 11572 11620
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 14464 11636 14516 11688
rect 15200 11568 15252 11620
rect 11428 11500 11480 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 2320 11296 2372 11348
rect 2504 11296 2556 11348
rect 4528 11296 4580 11348
rect 4896 11296 4948 11348
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 8208 11296 8260 11348
rect 10140 11296 10192 11348
rect 11060 11296 11112 11348
rect 3700 11160 3752 11212
rect 7748 11228 7800 11280
rect 8484 11228 8536 11280
rect 6276 11160 6328 11212
rect 6460 11160 6512 11212
rect 8208 11160 8260 11212
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 1952 11024 2004 11076
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 5540 11135 5592 11144
rect 5540 11101 5558 11135
rect 5558 11101 5592 11135
rect 5540 11092 5592 11101
rect 5448 11024 5500 11076
rect 1492 10956 1544 11008
rect 9680 11024 9732 11076
rect 10784 11092 10836 11144
rect 11520 11296 11572 11348
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 13084 11296 13136 11348
rect 13728 11296 13780 11348
rect 11612 11160 11664 11212
rect 14096 11228 14148 11280
rect 14372 11271 14424 11280
rect 14372 11237 14381 11271
rect 14381 11237 14415 11271
rect 14415 11237 14424 11271
rect 14372 11228 14424 11237
rect 15200 11203 15252 11212
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 15292 11092 15344 11144
rect 11428 11024 11480 11076
rect 12072 11024 12124 11076
rect 14188 11024 14240 11076
rect 5816 10956 5868 11008
rect 6460 10956 6512 11008
rect 6644 10956 6696 11008
rect 11244 10956 11296 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 14372 10956 14424 11008
rect 14556 10999 14608 11008
rect 14556 10965 14565 10999
rect 14565 10965 14599 10999
rect 14599 10965 14608 10999
rect 14556 10956 14608 10965
rect 15660 10956 15712 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 2228 10752 2280 10804
rect 2688 10752 2740 10804
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 3608 10659 3660 10668
rect 3608 10625 3626 10659
rect 3626 10625 3660 10659
rect 3884 10659 3936 10668
rect 3608 10616 3660 10625
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 4252 10752 4304 10804
rect 6000 10752 6052 10804
rect 5540 10684 5592 10736
rect 6184 10684 6236 10736
rect 6460 10752 6512 10804
rect 8852 10684 8904 10736
rect 10232 10752 10284 10804
rect 10968 10752 11020 10804
rect 11980 10752 12032 10804
rect 12348 10752 12400 10804
rect 13084 10795 13136 10804
rect 13084 10761 13093 10795
rect 13093 10761 13127 10795
rect 13127 10761 13136 10795
rect 13084 10752 13136 10761
rect 3884 10616 3936 10625
rect 1400 10548 1452 10600
rect 8760 10616 8812 10668
rect 9404 10616 9456 10668
rect 10232 10616 10284 10668
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 13636 10684 13688 10736
rect 13820 10684 13872 10736
rect 14096 10752 14148 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15752 10752 15804 10804
rect 14556 10684 14608 10736
rect 14648 10616 14700 10668
rect 2504 10455 2556 10464
rect 2504 10421 2513 10455
rect 2513 10421 2547 10455
rect 2547 10421 2556 10455
rect 2504 10412 2556 10421
rect 7656 10412 7708 10464
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 8300 10412 8352 10464
rect 9772 10480 9824 10532
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 13360 10548 13412 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 4252 10208 4304 10260
rect 4068 10140 4120 10192
rect 5264 9936 5316 9988
rect 8116 10208 8168 10260
rect 9220 10208 9272 10260
rect 11428 10251 11480 10260
rect 7656 10140 7708 10192
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 11612 10208 11664 10260
rect 12348 10208 12400 10260
rect 7104 10072 7156 10124
rect 7380 10072 7432 10124
rect 10876 10115 10928 10124
rect 10876 10081 10885 10115
rect 10885 10081 10919 10115
rect 10919 10081 10928 10115
rect 10876 10072 10928 10081
rect 10968 10072 11020 10124
rect 12900 10072 12952 10124
rect 14556 10208 14608 10260
rect 13820 10072 13872 10124
rect 14464 10115 14516 10124
rect 14464 10081 14473 10115
rect 14473 10081 14507 10115
rect 14507 10081 14516 10115
rect 15108 10115 15160 10124
rect 14464 10072 14516 10081
rect 14740 10004 14792 10056
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 6000 9936 6052 9988
rect 6460 9936 6512 9988
rect 9220 9936 9272 9988
rect 2596 9868 2648 9920
rect 7196 9868 7248 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 9680 9868 9732 9920
rect 10140 9936 10192 9988
rect 13176 9936 13228 9988
rect 13544 9936 13596 9988
rect 10508 9868 10560 9920
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 12992 9868 13044 9920
rect 15752 9936 15804 9988
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 2780 9596 2832 9648
rect 5172 9664 5224 9716
rect 3332 9596 3384 9648
rect 6644 9664 6696 9716
rect 7196 9664 7248 9716
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 2596 9528 2648 9580
rect 4620 9528 4672 9580
rect 7472 9596 7524 9648
rect 9680 9664 9732 9716
rect 12716 9707 12768 9716
rect 10508 9596 10560 9648
rect 12716 9673 12725 9707
rect 12725 9673 12759 9707
rect 12759 9673 12768 9707
rect 12716 9664 12768 9673
rect 12992 9707 13044 9716
rect 12992 9673 13001 9707
rect 13001 9673 13035 9707
rect 13035 9673 13044 9707
rect 12992 9664 13044 9673
rect 13176 9707 13228 9716
rect 13176 9673 13185 9707
rect 13185 9673 13219 9707
rect 13219 9673 13228 9707
rect 13176 9664 13228 9673
rect 12900 9596 12952 9648
rect 13360 9596 13412 9648
rect 6644 9571 6696 9580
rect 6644 9537 6678 9571
rect 6678 9537 6696 9571
rect 6644 9528 6696 9537
rect 7840 9528 7892 9580
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 13452 9528 13504 9580
rect 15200 9596 15252 9648
rect 11060 9503 11112 9512
rect 5080 9324 5132 9376
rect 5448 9324 5500 9376
rect 7840 9324 7892 9376
rect 9312 9324 9364 9376
rect 9588 9324 9640 9376
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 11704 9392 11756 9444
rect 12532 9460 12584 9512
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 12716 9392 12768 9444
rect 13820 9392 13872 9444
rect 15016 9392 15068 9444
rect 12072 9324 12124 9376
rect 13636 9324 13688 9376
rect 14464 9324 14516 9376
rect 14556 9324 14608 9376
rect 15384 9324 15436 9376
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 6000 9120 6052 9172
rect 5632 9052 5684 9104
rect 7104 9095 7156 9104
rect 7104 9061 7113 9095
rect 7113 9061 7147 9095
rect 7147 9061 7156 9095
rect 7104 9052 7156 9061
rect 8852 9120 8904 9172
rect 10968 9052 11020 9104
rect 14648 9120 14700 9172
rect 3884 8984 3936 9036
rect 5448 8984 5500 9036
rect 9036 8984 9088 9036
rect 9588 8984 9640 9036
rect 2136 8916 2188 8968
rect 2688 8848 2740 8900
rect 5448 8848 5500 8900
rect 6736 8916 6788 8968
rect 8852 8916 8904 8968
rect 11060 8916 11112 8968
rect 5816 8848 5868 8900
rect 6184 8848 6236 8900
rect 9772 8848 9824 8900
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4620 8780 4672 8832
rect 11980 8984 12032 9036
rect 11244 8916 11296 8968
rect 12900 8984 12952 9036
rect 13452 9052 13504 9104
rect 13728 9095 13780 9104
rect 13728 9061 13737 9095
rect 13737 9061 13771 9095
rect 13771 9061 13780 9095
rect 13728 9052 13780 9061
rect 15292 9120 15344 9172
rect 15108 9052 15160 9104
rect 15476 9052 15528 9104
rect 16396 9052 16448 9104
rect 12532 8916 12584 8968
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 13728 8848 13780 8900
rect 15476 8916 15528 8968
rect 15292 8848 15344 8900
rect 11428 8780 11480 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 13084 8780 13136 8832
rect 13636 8780 13688 8832
rect 13820 8780 13872 8832
rect 14924 8780 14976 8832
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 2688 8576 2740 8628
rect 3148 8576 3200 8628
rect 8852 8619 8904 8628
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 7104 8508 7156 8560
rect 9956 8576 10008 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 12808 8619 12860 8628
rect 12808 8585 12817 8619
rect 12817 8585 12851 8619
rect 12851 8585 12860 8619
rect 12808 8576 12860 8585
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 4160 8440 4212 8492
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 11704 8508 11756 8560
rect 13176 8508 13228 8560
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 14832 8508 14884 8560
rect 2136 8372 2188 8424
rect 5816 8372 5868 8424
rect 8852 8440 8904 8492
rect 7932 8372 7984 8424
rect 12900 8440 12952 8492
rect 10048 8372 10100 8424
rect 13360 8372 13412 8424
rect 14740 8372 14792 8424
rect 3884 8304 3936 8356
rect 4252 8304 4304 8356
rect 5448 8304 5500 8356
rect 6644 8304 6696 8356
rect 5080 8236 5132 8288
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 11336 8236 11388 8288
rect 14004 8236 14056 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 1676 8032 1728 8084
rect 6184 8032 6236 8084
rect 7380 8032 7432 8084
rect 8852 8032 8904 8084
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 3332 7964 3384 8016
rect 9404 7964 9456 8016
rect 11612 8032 11664 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 2136 7896 2188 7948
rect 2504 7896 2556 7948
rect 5448 7896 5500 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 4252 7828 4304 7880
rect 5632 7828 5684 7880
rect 9036 7828 9088 7880
rect 9128 7828 9180 7880
rect 11244 7896 11296 7948
rect 12900 7896 12952 7948
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 14832 7896 14884 7948
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 3884 7760 3936 7812
rect 4620 7803 4672 7812
rect 4620 7769 4654 7803
rect 4654 7769 4672 7803
rect 4620 7760 4672 7769
rect 3700 7692 3752 7744
rect 4160 7692 4212 7744
rect 9772 7760 9824 7812
rect 11060 7760 11112 7812
rect 12440 7760 12492 7812
rect 12808 7760 12860 7812
rect 14280 7760 14332 7812
rect 8116 7692 8168 7744
rect 11244 7692 11296 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 13544 7692 13596 7744
rect 15200 7692 15252 7744
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 3240 7488 3292 7540
rect 12624 7488 12676 7540
rect 13176 7531 13228 7540
rect 13176 7497 13185 7531
rect 13185 7497 13219 7531
rect 13219 7497 13228 7531
rect 13176 7488 13228 7497
rect 13544 7531 13596 7540
rect 13544 7497 13553 7531
rect 13553 7497 13587 7531
rect 13587 7497 13596 7531
rect 13544 7488 13596 7497
rect 14280 7531 14332 7540
rect 14280 7497 14289 7531
rect 14289 7497 14323 7531
rect 14323 7497 14332 7531
rect 14280 7488 14332 7497
rect 15200 7488 15252 7540
rect 16120 7488 16172 7540
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 6276 7420 6328 7472
rect 8024 7463 8076 7472
rect 8024 7429 8058 7463
rect 8058 7429 8076 7463
rect 8024 7420 8076 7429
rect 9128 7420 9180 7472
rect 11244 7463 11296 7472
rect 11244 7429 11253 7463
rect 11253 7429 11287 7463
rect 11287 7429 11296 7463
rect 11244 7420 11296 7429
rect 11980 7420 12032 7472
rect 5080 7395 5132 7404
rect 5080 7361 5114 7395
rect 5114 7361 5132 7395
rect 5080 7352 5132 7361
rect 7840 7352 7892 7404
rect 6092 7284 6144 7336
rect 3240 7148 3292 7200
rect 5172 7148 5224 7200
rect 7104 7216 7156 7268
rect 11612 7284 11664 7336
rect 13820 7420 13872 7472
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 13636 7327 13688 7336
rect 13636 7293 13645 7327
rect 13645 7293 13679 7327
rect 13679 7293 13688 7327
rect 13636 7284 13688 7293
rect 14740 7327 14792 7336
rect 13452 7216 13504 7268
rect 14740 7293 14749 7327
rect 14749 7293 14783 7327
rect 14783 7293 14792 7327
rect 14740 7284 14792 7293
rect 14832 7327 14884 7336
rect 14832 7293 14841 7327
rect 14841 7293 14875 7327
rect 14875 7293 14884 7327
rect 14832 7284 14884 7293
rect 8668 7148 8720 7200
rect 9220 7148 9272 7200
rect 10140 7148 10192 7200
rect 11520 7191 11572 7200
rect 11520 7157 11529 7191
rect 11529 7157 11563 7191
rect 11563 7157 11572 7191
rect 11520 7148 11572 7157
rect 15292 7148 15344 7200
rect 15660 7148 15712 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 2504 6944 2556 6996
rect 4160 6944 4212 6996
rect 4804 6944 4856 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 3608 6808 3660 6860
rect 7472 6944 7524 6996
rect 7840 6944 7892 6996
rect 8668 6987 8720 6996
rect 8668 6953 8677 6987
rect 8677 6953 8711 6987
rect 8711 6953 8720 6987
rect 8668 6944 8720 6953
rect 10232 6944 10284 6996
rect 12072 6944 12124 6996
rect 3516 6740 3568 6792
rect 3424 6672 3476 6724
rect 4252 6672 4304 6724
rect 4712 6740 4764 6792
rect 6000 6740 6052 6792
rect 6460 6740 6512 6792
rect 13636 6944 13688 6996
rect 14648 6944 14700 6996
rect 15108 6944 15160 6996
rect 11520 6851 11572 6860
rect 11520 6817 11529 6851
rect 11529 6817 11563 6851
rect 11563 6817 11572 6851
rect 11520 6808 11572 6817
rect 9220 6783 9272 6792
rect 7012 6715 7064 6724
rect 1952 6604 2004 6656
rect 2320 6604 2372 6656
rect 5816 6604 5868 6656
rect 7012 6681 7046 6715
rect 7046 6681 7064 6715
rect 7012 6672 7064 6681
rect 7656 6672 7708 6724
rect 8024 6672 8076 6724
rect 9220 6749 9254 6783
rect 9254 6749 9272 6783
rect 9220 6740 9272 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 13084 6808 13136 6860
rect 13820 6808 13872 6860
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 14096 6808 14148 6860
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 14832 6808 14884 6860
rect 15476 6851 15528 6860
rect 12716 6740 12768 6792
rect 13360 6740 13412 6792
rect 7472 6604 7524 6656
rect 8208 6604 8260 6656
rect 8852 6604 8904 6656
rect 11520 6604 11572 6656
rect 14004 6672 14056 6724
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 15016 6740 15068 6792
rect 15292 6740 15344 6792
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 12072 6604 12124 6656
rect 12624 6604 12676 6656
rect 12900 6604 12952 6656
rect 13084 6604 13136 6656
rect 14556 6604 14608 6656
rect 14832 6604 14884 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 1584 6332 1636 6384
rect 3976 6400 4028 6452
rect 4068 6400 4120 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 5816 6400 5868 6452
rect 6000 6400 6052 6452
rect 7748 6400 7800 6452
rect 8852 6400 8904 6452
rect 9312 6400 9364 6452
rect 9588 6400 9640 6452
rect 11060 6400 11112 6452
rect 12440 6400 12492 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 13360 6400 13412 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14556 6400 14608 6452
rect 15292 6400 15344 6452
rect 2320 6332 2372 6384
rect 4252 6332 4304 6384
rect 3240 6307 3292 6316
rect 3240 6273 3274 6307
rect 3274 6273 3292 6307
rect 6092 6332 6144 6384
rect 7012 6332 7064 6384
rect 14648 6332 14700 6384
rect 3240 6264 3292 6273
rect 8300 6264 8352 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 12440 6264 12492 6316
rect 12624 6264 12676 6316
rect 12808 6264 12860 6316
rect 1492 6196 1544 6248
rect 2596 6196 2648 6248
rect 4068 6196 4120 6248
rect 5632 6196 5684 6248
rect 7104 6239 7156 6248
rect 2504 6128 2556 6180
rect 4620 6128 4672 6180
rect 5540 6128 5592 6180
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7380 6128 7432 6180
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 9312 6196 9364 6248
rect 10048 6128 10100 6180
rect 11428 6196 11480 6248
rect 13452 6239 13504 6248
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 14004 6196 14056 6248
rect 14096 6196 14148 6248
rect 15108 6196 15160 6248
rect 3240 6060 3292 6112
rect 4712 6060 4764 6112
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 11704 6060 11756 6112
rect 13728 6128 13780 6180
rect 11888 6060 11940 6112
rect 12716 6060 12768 6112
rect 12808 6060 12860 6112
rect 13544 6060 13596 6112
rect 14832 6060 14884 6112
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 1676 5856 1728 5908
rect 2596 5899 2648 5908
rect 2596 5865 2605 5899
rect 2605 5865 2639 5899
rect 2639 5865 2648 5899
rect 2596 5856 2648 5865
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 4804 5856 4856 5908
rect 5080 5856 5132 5908
rect 7748 5856 7800 5908
rect 9312 5856 9364 5908
rect 9772 5856 9824 5908
rect 12072 5856 12124 5908
rect 13268 5856 13320 5908
rect 14740 5856 14792 5908
rect 2136 5763 2188 5772
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 5908 5788 5960 5840
rect 2136 5720 2188 5729
rect 3608 5720 3660 5772
rect 4436 5720 4488 5772
rect 4712 5763 4764 5772
rect 4712 5729 4721 5763
rect 4721 5729 4755 5763
rect 4755 5729 4764 5763
rect 4712 5720 4764 5729
rect 5356 5720 5408 5772
rect 5816 5720 5868 5772
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 6276 5720 6328 5772
rect 7288 5720 7340 5772
rect 2780 5584 2832 5636
rect 7656 5720 7708 5772
rect 7932 5720 7984 5772
rect 6000 5584 6052 5636
rect 9128 5652 9180 5704
rect 9496 5720 9548 5772
rect 10324 5720 10376 5772
rect 11336 5720 11388 5772
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11796 5788 11848 5840
rect 13820 5788 13872 5840
rect 12348 5720 12400 5772
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 9588 5652 9640 5704
rect 13544 5695 13596 5704
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4620 5559 4672 5568
rect 4620 5525 4629 5559
rect 4629 5525 4663 5559
rect 4663 5525 4672 5559
rect 4620 5516 4672 5525
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 6368 5516 6420 5568
rect 7472 5584 7524 5636
rect 7564 5584 7616 5636
rect 8852 5584 8904 5636
rect 10784 5584 10836 5636
rect 11612 5584 11664 5636
rect 12072 5584 12124 5636
rect 7840 5516 7892 5568
rect 9220 5516 9272 5568
rect 9772 5516 9824 5568
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 10968 5559 11020 5568
rect 10968 5525 10977 5559
rect 10977 5525 11011 5559
rect 11011 5525 11020 5559
rect 10968 5516 11020 5525
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 14372 5652 14424 5704
rect 15752 5652 15804 5704
rect 13360 5584 13412 5636
rect 12624 5516 12676 5525
rect 13912 5516 13964 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 15292 5516 15344 5568
rect 16120 5516 16172 5568
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 4068 5312 4120 5364
rect 4252 5312 4304 5364
rect 5448 5312 5500 5364
rect 7104 5312 7156 5364
rect 7932 5355 7984 5364
rect 7932 5321 7941 5355
rect 7941 5321 7975 5355
rect 7975 5321 7984 5355
rect 7932 5312 7984 5321
rect 8300 5312 8352 5364
rect 2688 5287 2740 5296
rect 2688 5253 2697 5287
rect 2697 5253 2731 5287
rect 2731 5253 2740 5287
rect 2688 5244 2740 5253
rect 3148 5176 3200 5228
rect 3608 5244 3660 5296
rect 6736 5287 6788 5296
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 4712 5176 4764 5228
rect 5448 5176 5500 5228
rect 6736 5253 6745 5287
rect 6745 5253 6779 5287
rect 6779 5253 6788 5287
rect 6736 5244 6788 5253
rect 9312 5244 9364 5296
rect 9588 5287 9640 5296
rect 9588 5253 9597 5287
rect 9597 5253 9631 5287
rect 9631 5253 9640 5287
rect 9588 5244 9640 5253
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 10968 5312 11020 5364
rect 11612 5355 11664 5364
rect 11612 5321 11621 5355
rect 11621 5321 11655 5355
rect 11655 5321 11664 5355
rect 11612 5312 11664 5321
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 13452 5312 13504 5364
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 14372 5312 14424 5364
rect 14556 5312 14608 5364
rect 15016 5355 15068 5364
rect 15016 5321 15025 5355
rect 15025 5321 15059 5355
rect 15059 5321 15068 5355
rect 15016 5312 15068 5321
rect 15936 5312 15988 5364
rect 10140 5244 10192 5296
rect 13544 5244 13596 5296
rect 15200 5244 15252 5296
rect 15476 5244 15528 5296
rect 7012 5176 7064 5228
rect 8208 5176 8260 5228
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 10508 5176 10560 5228
rect 11612 5176 11664 5228
rect 12072 5176 12124 5228
rect 14280 5176 14332 5228
rect 14740 5176 14792 5228
rect 15016 5176 15068 5228
rect 3976 5108 4028 5160
rect 3516 4972 3568 5024
rect 3976 4972 4028 5024
rect 4068 4972 4120 5024
rect 5540 5108 5592 5160
rect 5908 5108 5960 5160
rect 6184 5108 6236 5160
rect 7472 5108 7524 5160
rect 5724 5040 5776 5092
rect 6000 5040 6052 5092
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9404 5151 9456 5160
rect 9036 5108 9088 5117
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 9772 5108 9824 5160
rect 11796 5108 11848 5160
rect 13452 5151 13504 5160
rect 10140 5040 10192 5092
rect 12072 5040 12124 5092
rect 8392 4972 8444 5024
rect 9312 4972 9364 5024
rect 11980 4972 12032 5024
rect 12624 4972 12676 5024
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 12808 5040 12860 5092
rect 13636 5108 13688 5160
rect 15292 5108 15344 5160
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 4160 4811 4212 4820
rect 4160 4777 4169 4811
rect 4169 4777 4203 4811
rect 4203 4777 4212 4811
rect 4160 4768 4212 4777
rect 5080 4768 5132 4820
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 3976 4743 4028 4752
rect 3976 4709 3985 4743
rect 3985 4709 4019 4743
rect 4019 4709 4028 4743
rect 3976 4700 4028 4709
rect 7748 4768 7800 4820
rect 7932 4768 7984 4820
rect 8208 4768 8260 4820
rect 8852 4768 8904 4820
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10876 4768 10928 4820
rect 13636 4811 13688 4820
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4160 4632 4212 4684
rect 6920 4700 6972 4752
rect 6092 4675 6144 4684
rect 2136 4607 2188 4616
rect 2136 4573 2145 4607
rect 2145 4573 2179 4607
rect 2179 4573 2188 4607
rect 2136 4564 2188 4573
rect 3148 4564 3200 4616
rect 4252 4564 4304 4616
rect 5080 4564 5132 4616
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 8116 4700 8168 4752
rect 10324 4700 10376 4752
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 11980 4700 12032 4752
rect 12532 4700 12584 4752
rect 13084 4700 13136 4752
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 8392 4675 8444 4684
rect 8392 4641 8401 4675
rect 8401 4641 8435 4675
rect 8435 4641 8444 4675
rect 8392 4632 8444 4641
rect 9220 4632 9272 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 5908 4564 5960 4616
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 2228 4496 2280 4548
rect 8300 4564 8352 4616
rect 9036 4564 9088 4616
rect 9588 4564 9640 4616
rect 9864 4564 9916 4616
rect 11244 4564 11296 4616
rect 13820 4632 13872 4684
rect 15108 4632 15160 4684
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 15660 4564 15712 4616
rect 16396 4564 16448 4616
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 3148 4471 3200 4480
rect 2780 4428 2832 4437
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 4436 4428 4488 4480
rect 4528 4428 4580 4480
rect 4712 4428 4764 4480
rect 5080 4428 5132 4480
rect 6276 4428 6328 4480
rect 12716 4496 12768 4548
rect 7656 4428 7708 4480
rect 9036 4428 9088 4480
rect 9864 4428 9916 4480
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11612 4471 11664 4480
rect 11244 4428 11296 4437
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 2136 4224 2188 4276
rect 3148 4224 3200 4276
rect 3240 4267 3292 4276
rect 3240 4233 3249 4267
rect 3249 4233 3283 4267
rect 3283 4233 3292 4267
rect 3240 4224 3292 4233
rect 3700 4224 3752 4276
rect 3976 4224 4028 4276
rect 4528 4224 4580 4276
rect 6276 4224 6328 4276
rect 7196 4224 7248 4276
rect 7472 4224 7524 4276
rect 8116 4224 8168 4276
rect 8300 4224 8352 4276
rect 9956 4224 10008 4276
rect 10968 4224 11020 4276
rect 11244 4224 11296 4276
rect 2504 4156 2556 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 2136 4088 2188 4140
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2780 4088 2832 4140
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 3700 4020 3752 4072
rect 3884 4088 3936 4140
rect 4160 4156 4212 4208
rect 4988 4156 5040 4208
rect 8760 4156 8812 4208
rect 10140 4156 10192 4208
rect 4896 4020 4948 4072
rect 5356 4020 5408 4072
rect 5632 4020 5684 4072
rect 4620 3952 4672 4004
rect 4804 3952 4856 4004
rect 5816 4063 5868 4072
rect 5816 4029 5825 4063
rect 5825 4029 5859 4063
rect 5859 4029 5868 4063
rect 6092 4088 6144 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10784 4156 10836 4208
rect 12164 4199 12216 4208
rect 12164 4165 12173 4199
rect 12173 4165 12207 4199
rect 12207 4165 12216 4199
rect 12716 4224 12768 4276
rect 14924 4224 14976 4276
rect 15200 4224 15252 4276
rect 16120 4224 16172 4276
rect 12164 4156 12216 4165
rect 13176 4156 13228 4208
rect 14464 4156 14516 4208
rect 10692 4088 10744 4140
rect 11980 4088 12032 4140
rect 12440 4088 12492 4140
rect 13268 4088 13320 4140
rect 13728 4088 13780 4140
rect 14648 4156 14700 4208
rect 14832 4088 14884 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 8208 4063 8260 4072
rect 5816 4020 5868 4029
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 11796 4020 11848 4072
rect 3976 3884 4028 3936
rect 4160 3884 4212 3936
rect 4712 3884 4764 3936
rect 9864 3952 9916 4004
rect 6184 3884 6236 3936
rect 9404 3884 9456 3936
rect 11060 3884 11112 3936
rect 11244 3952 11296 4004
rect 14372 4020 14424 4072
rect 14556 4020 14608 4072
rect 13820 3952 13872 4004
rect 11336 3884 11388 3936
rect 11704 3884 11756 3936
rect 12164 3884 12216 3936
rect 12716 3884 12768 3936
rect 14832 3884 14884 3936
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 2504 3680 2556 3732
rect 3424 3680 3476 3732
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 4804 3680 4856 3732
rect 5080 3680 5132 3732
rect 5448 3680 5500 3732
rect 7012 3680 7064 3732
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 8760 3680 8812 3732
rect 9312 3680 9364 3732
rect 9588 3680 9640 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 10968 3680 11020 3732
rect 11704 3680 11756 3732
rect 12072 3680 12124 3732
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12716 3723 12768 3732
rect 12440 3680 12492 3689
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 4528 3612 4580 3664
rect 4068 3544 4120 3596
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 6460 3544 6512 3596
rect 2504 3519 2556 3528
rect 2504 3485 2513 3519
rect 2513 3485 2547 3519
rect 2547 3485 2556 3519
rect 2504 3476 2556 3485
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 3056 3408 3108 3460
rect 2044 3340 2096 3392
rect 2504 3340 2556 3392
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 3516 3340 3568 3349
rect 3700 3408 3752 3460
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6368 3476 6420 3528
rect 9680 3612 9732 3664
rect 9956 3655 10008 3664
rect 9956 3621 9965 3655
rect 9965 3621 9999 3655
rect 9999 3621 10008 3655
rect 9956 3612 10008 3621
rect 10876 3612 10928 3664
rect 11060 3612 11112 3664
rect 13268 3680 13320 3732
rect 13636 3680 13688 3732
rect 13728 3680 13780 3732
rect 14464 3680 14516 3732
rect 15476 3680 15528 3732
rect 15752 3680 15804 3732
rect 7564 3587 7616 3596
rect 7564 3553 7573 3587
rect 7573 3553 7607 3587
rect 7607 3553 7616 3587
rect 7564 3544 7616 3553
rect 8024 3544 8076 3596
rect 8208 3544 8260 3596
rect 10048 3544 10100 3596
rect 11244 3544 11296 3596
rect 14004 3544 14056 3596
rect 7748 3476 7800 3528
rect 10232 3476 10284 3528
rect 11060 3476 11112 3528
rect 12440 3476 12492 3528
rect 13820 3476 13872 3528
rect 14832 3544 14884 3596
rect 15200 3587 15252 3596
rect 15200 3553 15209 3587
rect 15209 3553 15243 3587
rect 15243 3553 15252 3587
rect 15200 3544 15252 3553
rect 15108 3476 15160 3528
rect 4068 3340 4120 3392
rect 4160 3340 4212 3392
rect 6828 3408 6880 3460
rect 9588 3408 9640 3460
rect 10048 3408 10100 3460
rect 4896 3340 4948 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6276 3340 6328 3392
rect 6552 3383 6604 3392
rect 6552 3349 6561 3383
rect 6561 3349 6595 3383
rect 6595 3349 6604 3383
rect 6552 3340 6604 3349
rect 7932 3340 7984 3392
rect 9956 3340 10008 3392
rect 10692 3340 10744 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 14556 3340 14608 3392
rect 15752 3340 15804 3392
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 3424 3136 3476 3188
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 6552 3136 6604 3188
rect 6828 3136 6880 3188
rect 2412 3068 2464 3120
rect 4528 3068 4580 3120
rect 9956 3136 10008 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 11980 3179 12032 3188
rect 11980 3145 11989 3179
rect 11989 3145 12023 3179
rect 12023 3145 12032 3179
rect 11980 3136 12032 3145
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 12348 3111 12400 3120
rect 2228 3000 2280 3052
rect 2504 3000 2556 3052
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3516 3000 3568 3052
rect 3608 3000 3660 3052
rect 3884 3000 3936 3052
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2596 2864 2648 2916
rect 3148 2932 3200 2984
rect 4344 3000 4396 3052
rect 4712 2975 4764 2984
rect 4712 2941 4721 2975
rect 4721 2941 4755 2975
rect 4755 2941 4764 2975
rect 4712 2932 4764 2941
rect 5080 2932 5132 2984
rect 6184 3000 6236 3052
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 7932 3000 7984 3052
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 4252 2864 4304 2916
rect 6092 2932 6144 2984
rect 6920 2932 6972 2984
rect 7288 2932 7340 2984
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 7564 2932 7616 2984
rect 12348 3077 12357 3111
rect 12357 3077 12391 3111
rect 12391 3077 12400 3111
rect 12348 3068 12400 3077
rect 13084 3068 13136 3120
rect 14740 3136 14792 3188
rect 14464 3068 14516 3120
rect 8484 3000 8536 3052
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 10692 3000 10744 3052
rect 11244 3000 11296 3052
rect 5632 2864 5684 2916
rect 9680 2932 9732 2984
rect 11060 2932 11112 2984
rect 12440 3000 12492 3052
rect 13452 3000 13504 3052
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 14556 3000 14608 3052
rect 3240 2839 3292 2848
rect 3240 2805 3249 2839
rect 3249 2805 3283 2839
rect 3283 2805 3292 2839
rect 3240 2796 3292 2805
rect 4068 2796 4120 2848
rect 5448 2796 5500 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 6460 2796 6512 2848
rect 10692 2796 10744 2848
rect 11520 2864 11572 2916
rect 12348 2864 12400 2916
rect 12716 2932 12768 2984
rect 13912 2975 13964 2984
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 14004 2864 14056 2916
rect 14740 2864 14792 2916
rect 13728 2796 13780 2848
rect 15476 3000 15528 3052
rect 15660 3000 15712 3052
rect 15384 2907 15436 2916
rect 15384 2873 15393 2907
rect 15393 2873 15427 2907
rect 15427 2873 15436 2907
rect 15384 2864 15436 2873
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 3332 2592 3384 2644
rect 3884 2592 3936 2644
rect 4252 2592 4304 2644
rect 4712 2592 4764 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 1860 2524 1912 2576
rect 2872 2524 2924 2576
rect 5724 2524 5776 2576
rect 2688 2388 2740 2440
rect 5264 2456 5316 2508
rect 5356 2456 5408 2508
rect 5908 2524 5960 2576
rect 4068 2388 4120 2440
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 3332 2320 3384 2372
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 3608 2295 3660 2304
rect 3608 2261 3617 2295
rect 3617 2261 3651 2295
rect 3651 2261 3660 2295
rect 3608 2252 3660 2261
rect 5816 2388 5868 2440
rect 6000 2456 6052 2508
rect 7104 2456 7156 2508
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 9680 2524 9732 2576
rect 10784 2592 10836 2644
rect 11520 2635 11572 2644
rect 11520 2601 11529 2635
rect 11529 2601 11563 2635
rect 11563 2601 11572 2635
rect 11520 2592 11572 2601
rect 12348 2592 12400 2644
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13268 2592 13320 2644
rect 13360 2592 13412 2644
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 15292 2524 15344 2576
rect 8484 2456 8536 2508
rect 9036 2388 9088 2440
rect 9496 2456 9548 2508
rect 9312 2388 9364 2440
rect 10784 2456 10836 2508
rect 10232 2388 10284 2440
rect 12624 2456 12676 2508
rect 13636 2456 13688 2508
rect 13268 2388 13320 2440
rect 13820 2388 13872 2440
rect 16028 2456 16080 2508
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 15844 2388 15896 2440
rect 5356 2320 5408 2372
rect 6000 2252 6052 2304
rect 8208 2320 8260 2372
rect 9128 2252 9180 2304
rect 9680 2252 9732 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 11244 2252 11296 2304
rect 11796 2295 11848 2304
rect 11796 2261 11805 2295
rect 11805 2261 11839 2295
rect 11839 2261 11848 2295
rect 11796 2252 11848 2261
rect 11888 2252 11940 2304
rect 12440 2320 12492 2372
rect 14556 2320 14608 2372
rect 15016 2320 15068 2372
rect 15292 2320 15344 2372
rect 12900 2252 12952 2304
rect 13452 2295 13504 2304
rect 13452 2261 13461 2295
rect 13461 2261 13495 2295
rect 13495 2261 13504 2295
rect 13452 2252 13504 2261
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 5080 2048 5132 2100
rect 11796 2048 11848 2100
rect 4528 1980 4580 2032
rect 9956 1980 10008 2032
rect 6460 1912 6512 1964
rect 11888 1912 11940 1964
rect 3608 1844 3660 1896
rect 9864 1844 9916 1896
rect 2504 1776 2556 1828
rect 13084 1776 13136 1828
rect 13452 1776 13504 1828
rect 2136 1640 2188 1692
rect 11612 1640 11664 1692
rect 11244 1436 11296 1488
rect 13912 1436 13964 1488
rect 15200 1436 15252 1488
rect 6092 1368 6144 1420
rect 7840 1368 7892 1420
<< metal2 >>
rect 294 19200 350 20000
rect 662 19200 718 20000
rect 1030 19200 1086 20000
rect 1136 19230 1348 19258
rect 308 15366 336 19200
rect 676 17542 704 19200
rect 1044 19122 1072 19200
rect 1136 19122 1164 19230
rect 1044 19094 1164 19122
rect 664 17536 716 17542
rect 664 17478 716 17484
rect 1320 17354 1348 19230
rect 1398 19200 1454 20000
rect 1504 19230 1716 19258
rect 1412 19122 1440 19200
rect 1504 19122 1532 19230
rect 1412 19094 1532 19122
rect 1582 18048 1638 18057
rect 1582 17983 1638 17992
rect 1320 17326 1440 17354
rect 1412 17270 1440 17326
rect 1400 17264 1452 17270
rect 1400 17206 1452 17212
rect 1596 16590 1624 17983
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1688 16017 1716 19230
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4448 19230 4660 19258
rect 1780 16289 1808 19200
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16590 2084 16934
rect 2148 16810 2176 19200
rect 2516 17338 2544 19200
rect 2778 19000 2834 19009
rect 2778 18935 2834 18944
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2608 16946 2636 17206
rect 2792 17202 2820 18935
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2884 17066 2912 19200
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 3160 16998 3188 17138
rect 3148 16992 3200 16998
rect 2608 16918 2728 16946
rect 3148 16934 3200 16940
rect 2148 16782 2268 16810
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1766 16280 1822 16289
rect 1766 16215 1822 16224
rect 1674 16008 1730 16017
rect 1674 15943 1730 15952
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 296 15360 348 15366
rect 296 15302 348 15308
rect 1412 14249 1440 15370
rect 1964 15162 1992 15846
rect 2056 15570 2084 16526
rect 2240 16522 2268 16782
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2148 16153 2176 16458
rect 2134 16144 2190 16153
rect 2134 16079 2190 16088
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2332 15706 2360 16050
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1398 14240 1454 14249
rect 1398 14175 1454 14184
rect 1596 13394 1624 14894
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1688 13297 1716 13806
rect 1674 13288 1730 13297
rect 1674 13223 1730 13232
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12442 1440 12786
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1596 11393 1624 12718
rect 1582 11384 1638 11393
rect 1582 11319 1638 11328
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10674 1532 10950
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1400 10600 1452 10606
rect 1780 10554 1808 14282
rect 1964 12850 1992 14350
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11898 1992 12038
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1400 10542 1452 10548
rect 1412 9489 1440 10542
rect 1504 10526 1808 10554
rect 1398 9480 1454 9489
rect 1398 9415 1454 9424
rect 1504 6254 1532 10526
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 8090 1716 9454
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1596 6390 1624 7511
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1688 5914 1716 7686
rect 1780 7449 1808 9522
rect 1964 8537 1992 11018
rect 2056 8945 2084 15506
rect 2516 15502 2544 15982
rect 2412 15496 2464 15502
rect 2410 15464 2412 15473
rect 2504 15496 2556 15502
rect 2464 15464 2466 15473
rect 2504 15438 2556 15444
rect 2410 15399 2466 15408
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2332 14906 2360 15302
rect 2410 15192 2466 15201
rect 2410 15127 2466 15136
rect 2424 15094 2452 15127
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2516 15026 2544 15302
rect 2608 15162 2636 16526
rect 2700 16114 2728 16918
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2792 15994 2820 16458
rect 3252 16454 3280 19200
rect 3620 17338 3648 19200
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 2700 15966 2820 15994
rect 2700 15366 2728 15966
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2792 15434 2820 15642
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2332 14878 2452 14906
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2148 11898 2176 14758
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11898 2268 12242
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2332 11762 2360 13126
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2136 8968 2188 8974
rect 2042 8936 2098 8945
rect 2136 8910 2188 8916
rect 2042 8871 2098 8880
rect 1950 8528 2006 8537
rect 1950 8463 2006 8472
rect 2148 8430 2176 8910
rect 2240 8537 2268 10746
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 1766 7440 1822 7449
rect 1766 7375 1822 7384
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1676 5908 1728 5914
rect 1676 5850 1728 5856
rect 1964 5778 1992 6598
rect 2148 5778 2176 7890
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 6633 2268 7278
rect 2332 6662 2360 11290
rect 2320 6656 2372 6662
rect 2226 6624 2282 6633
rect 2320 6598 2372 6604
rect 2226 6559 2282 6568
rect 2332 6390 2360 6598
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1596 4146 1624 4655
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1872 3777 1900 4490
rect 2148 4282 2176 4558
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1858 3768 1914 3777
rect 1858 3703 1914 3712
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1780 1873 1808 2926
rect 1872 2825 1900 3402
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1858 2816 1914 2825
rect 1858 2751 1914 2760
rect 1860 2576 1912 2582
rect 1860 2518 1912 2524
rect 1766 1864 1822 1873
rect 1766 1799 1822 1808
rect 1872 1170 1900 2518
rect 1780 1142 1900 1170
rect 1780 800 1808 1142
rect 2056 800 2084 3334
rect 2148 1698 2176 4082
rect 2240 3058 2268 4490
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2332 4049 2360 4082
rect 2318 4040 2374 4049
rect 2318 3975 2374 3984
rect 2424 3126 2452 14878
rect 2516 11354 2544 14962
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2700 14346 2728 14826
rect 3160 14822 3188 16118
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2884 14414 2912 14554
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2884 14006 2912 14350
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 11694 2636 13330
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9674 2544 10406
rect 2608 9926 2636 11630
rect 2700 10810 2728 13262
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 2964 11144 3016 11150
rect 2962 11112 2964 11121
rect 3016 11112 3018 11121
rect 2962 11047 3018 11056
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2686 10432 2742 10441
rect 2686 10367 2742 10376
rect 2700 10180 2728 10367
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 2700 10152 2820 10180
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2516 9646 2636 9674
rect 2792 9654 2820 10152
rect 2516 7954 2544 9646
rect 2608 9586 2636 9646
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 2686 9072 2742 9081
rect 2686 9007 2742 9016
rect 2700 8906 2728 9007
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 3160 8634 3188 14758
rect 3344 12434 3372 17138
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 16182 3648 16526
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3608 16176 3660 16182
rect 3608 16118 3660 16124
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3620 14278 3648 14962
rect 3608 14272 3660 14278
rect 3606 14240 3608 14249
rect 3660 14240 3662 14249
rect 3606 14175 3662 14184
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3528 13734 3556 13942
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3712 13326 3740 16390
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3804 12434 3832 16934
rect 3988 16538 4016 19200
rect 4356 17338 4384 19200
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4172 17105 4200 17138
rect 4252 17128 4304 17134
rect 4158 17096 4214 17105
rect 4252 17070 4304 17076
rect 4158 17031 4214 17040
rect 3988 16522 4108 16538
rect 3988 16516 4120 16522
rect 3988 16510 4068 16516
rect 4068 16458 4120 16464
rect 4158 15600 4214 15609
rect 4158 15535 4160 15544
rect 4212 15535 4214 15544
rect 4160 15506 4212 15512
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4080 15094 4108 15302
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4080 13938 4108 14554
rect 4172 14278 4200 15370
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14074 4200 14214
rect 4264 14074 4292 17070
rect 4448 16538 4476 19230
rect 4632 19122 4660 19230
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11440 19230 11652 19258
rect 4724 19122 4752 19200
rect 4632 19094 4752 19122
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 4356 16510 4476 16538
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4356 16454 4384 16510
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4356 15502 4384 15846
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4356 15162 4384 15438
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4356 14618 4384 15098
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4448 14498 4476 15914
rect 4356 14470 4476 14498
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13394 4108 13874
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4066 13288 4122 13297
rect 4066 13223 4122 13232
rect 4080 12986 4108 13223
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4172 12850 4200 13466
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4264 12986 4292 13330
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3344 12406 3556 12434
rect 3804 12406 4016 12434
rect 3332 12368 3384 12374
rect 3238 12336 3294 12345
rect 3332 12310 3384 12316
rect 3238 12271 3294 12280
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 7002 2544 7346
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2516 4214 2544 6122
rect 2608 5914 2636 6190
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2700 5794 2728 8570
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 3252 7546 3280 12271
rect 3344 11762 3372 12310
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3344 8022 3372 9590
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 3252 6322 3280 7142
rect 3528 6798 3556 12406
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 10674 3648 12038
rect 3712 11218 3740 12174
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3620 6866 3648 10610
rect 3896 10266 3924 10610
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3698 8664 3754 8673
rect 3698 8599 3754 8608
rect 3712 7750 3740 8599
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 2608 5766 2728 5794
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2608 4078 2636 5766
rect 2686 5672 2742 5681
rect 2686 5607 2742 5616
rect 2780 5636 2832 5642
rect 2700 5302 2728 5607
rect 2780 5578 2832 5584
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2792 5114 2820 5578
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2700 5086 2820 5114
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2516 3534 2544 3674
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2516 3058 2544 3334
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2136 1692 2188 1698
rect 2136 1634 2188 1640
rect 2332 800 2360 2246
rect 2516 1834 2544 2994
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2504 1828 2556 1834
rect 2504 1770 2556 1776
rect 2608 800 2636 2858
rect 2700 2446 2728 5086
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 3160 4622 3188 5170
rect 3252 4690 3280 6054
rect 3436 5234 3464 6666
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3330 4720 3386 4729
rect 3240 4684 3292 4690
rect 3330 4655 3332 4664
rect 3240 4626 3292 4632
rect 3384 4655 3386 4664
rect 3332 4626 3384 4632
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 2792 4146 2820 4422
rect 3160 4282 3188 4422
rect 3238 4312 3294 4321
rect 3148 4276 3200 4282
rect 3238 4247 3240 4256
rect 3148 4218 3200 4224
rect 3292 4247 3294 4256
rect 3240 4218 3292 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 3058 3096 3402
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2884 800 2912 2518
rect 3160 800 3188 2926
rect 3240 2848 3292 2854
rect 3238 2816 3240 2825
rect 3292 2816 3294 2825
rect 3238 2751 3294 2760
rect 3344 2650 3372 4014
rect 3436 3738 3464 5170
rect 3528 5030 3556 6734
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3620 5302 3648 5714
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3712 4282 3740 7686
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3712 3641 3740 4014
rect 3698 3632 3754 3641
rect 3698 3567 3754 3576
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3344 2378 3372 2586
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 3436 800 3464 3130
rect 3528 3058 3556 3334
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3620 2310 3648 2994
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3620 1902 3648 2246
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3712 800 3740 3402
rect 3804 921 3832 8774
rect 3896 8362 3924 8978
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 4146 3924 7754
rect 3988 6610 4016 12406
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 10198 4108 12106
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4172 8498 4200 12582
rect 4264 12442 4292 12922
rect 4252 12436 4304 12442
rect 4356 12434 4384 14470
rect 4540 14226 4568 16186
rect 4632 15978 4660 16526
rect 5092 16454 5120 19200
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16590 5304 16934
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 5000 15910 5028 16050
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 4988 15904 5040 15910
rect 4986 15872 4988 15881
rect 5040 15872 5042 15881
rect 4986 15807 5042 15816
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 5092 15178 5120 15914
rect 5184 15366 5212 16390
rect 5276 16153 5304 16526
rect 5460 16250 5488 19200
rect 5724 16652 5776 16658
rect 5644 16612 5724 16640
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5262 16144 5318 16153
rect 5262 16079 5318 16088
rect 5552 15910 5580 16526
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15502 5580 15846
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5092 15150 5212 15178
rect 4540 14198 4660 14226
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13190 4476 13670
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4356 12406 4476 12434
rect 4252 12378 4304 12384
rect 4264 11830 4292 12378
rect 4342 12336 4398 12345
rect 4342 12271 4398 12280
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4264 10810 4292 11766
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4264 9518 4292 10202
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4172 7834 4200 8434
rect 4264 8362 4292 9454
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7886 4292 8298
rect 4080 7806 4200 7834
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4080 6882 4108 7806
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7002 4200 7686
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4080 6854 4200 6882
rect 3988 6582 4108 6610
rect 4080 6458 4108 6582
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3988 5166 4016 6394
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4080 5370 4108 6190
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3988 4758 4016 4966
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 4593 4016 4694
rect 3974 4584 4030 4593
rect 3974 4519 4030 4528
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3896 3058 3924 4082
rect 3988 3942 4016 4218
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3988 2938 4016 3674
rect 4080 3602 4108 4966
rect 4172 4826 4200 6854
rect 4264 6730 4292 7822
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4264 6390 4292 6666
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5370 4292 5510
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4172 4690 4200 4762
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4214 4200 4626
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4160 3936 4212 3942
rect 4158 3904 4160 3913
rect 4212 3904 4214 3913
rect 4158 3839 4214 3848
rect 4158 3768 4214 3777
rect 4158 3703 4214 3712
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4172 3482 4200 3703
rect 4080 3454 4200 3482
rect 4080 3398 4108 3454
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3210 4200 3334
rect 3896 2910 4016 2938
rect 4080 3182 4200 3210
rect 4264 3194 4292 4558
rect 4356 3602 4384 12271
rect 4448 11937 4476 12406
rect 4434 11928 4490 11937
rect 4434 11863 4490 11872
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4448 5778 4476 11766
rect 4540 11354 4568 13194
rect 4632 12322 4660 14198
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4816 12850 4844 12922
rect 5092 12850 5120 14010
rect 5184 13161 5212 15150
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5368 14362 5396 14962
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5276 14334 5396 14362
rect 5276 13530 5304 14334
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5170 13152 5226 13161
rect 5170 13087 5226 13096
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4724 12481 4752 12786
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4710 12472 4766 12481
rect 4710 12407 4766 12416
rect 4632 12294 4752 12322
rect 4724 12209 4752 12294
rect 4908 12238 4936 12582
rect 5184 12306 5212 12718
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4896 12232 4948 12238
rect 4710 12200 4766 12209
rect 4896 12174 4948 12180
rect 4710 12135 4766 12144
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 4802 11792 4858 11801
rect 4802 11727 4858 11736
rect 4896 11756 4948 11762
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4724 11257 4752 11494
rect 4710 11248 4766 11257
rect 4710 11183 4766 11192
rect 4816 10996 4844 11727
rect 4896 11698 4948 11704
rect 4908 11354 4936 11698
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4540 10968 4844 10996
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4540 5001 4568 10968
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4632 8838 4660 9522
rect 5092 9382 5120 12106
rect 5276 12102 5304 12543
rect 5264 12096 5316 12102
rect 5170 12064 5226 12073
rect 5264 12038 5316 12044
rect 5170 11999 5226 12008
rect 5184 9722 5212 11999
rect 5276 9994 5304 12038
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4632 6186 4660 7754
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 5092 7410 5120 8230
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 5080 7404 5132 7410
rect 5132 7364 5212 7392
rect 5080 7346 5132 7352
rect 4724 6984 4752 7346
rect 5184 7324 5212 7364
rect 5184 7296 5304 7324
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 4804 6996 4856 7002
rect 4724 6956 4804 6984
rect 4724 6798 4752 6956
rect 4804 6938 4856 6944
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4724 5778 4752 6054
rect 4816 5914 4844 6394
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4620 5568 4672 5574
rect 5092 5545 5120 5850
rect 4620 5510 4672 5516
rect 5078 5536 5134 5545
rect 4526 4992 4582 5001
rect 4526 4927 4582 4936
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3188 4304 3194
rect 3896 2650 3924 2910
rect 4080 2854 4108 3182
rect 4252 3130 4304 3136
rect 4158 3088 4214 3097
rect 4356 3058 4384 3538
rect 4158 3023 4214 3032
rect 4344 3052 4396 3058
rect 4068 2848 4120 2854
rect 3974 2816 4030 2825
rect 4068 2790 4120 2796
rect 3974 2751 4030 2760
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3790 912 3846 921
rect 3790 847 3846 856
rect 3988 800 4016 2751
rect 4080 2446 4108 2790
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4172 1714 4200 3023
rect 4344 2994 4396 3000
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4264 2650 4292 2858
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4448 2446 4476 4422
rect 4540 4282 4568 4422
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4526 4040 4582 4049
rect 4632 4010 4660 5510
rect 4698 5468 5006 5477
rect 5078 5471 5134 5480
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 4486 4752 5170
rect 5078 4856 5134 4865
rect 5078 4791 5080 4800
rect 5132 4791 5134 4800
rect 5080 4762 5132 4768
rect 5092 4622 5120 4762
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4896 4072 4948 4078
rect 4710 4040 4766 4049
rect 4526 3975 4582 3984
rect 4620 4004 4672 4010
rect 4540 3670 4568 3975
rect 4896 4014 4948 4020
rect 4710 3975 4766 3984
rect 4804 4004 4856 4010
rect 4620 3946 4672 3952
rect 4724 3942 4752 3975
rect 4804 3946 4856 3952
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4526 3496 4582 3505
rect 4724 3482 4752 3878
rect 4816 3738 4844 3946
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4526 3431 4582 3440
rect 4632 3454 4752 3482
rect 4540 3126 4568 3431
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4632 2825 4660 3454
rect 4908 3398 4936 4014
rect 5000 3482 5028 4150
rect 5092 3738 5120 4422
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5000 3454 5120 3482
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 5092 3108 5120 3454
rect 5000 3080 5120 3108
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4724 2650 4752 2926
rect 5000 2650 5028 3080
rect 5080 2984 5132 2990
rect 5184 2972 5212 7142
rect 5132 2944 5212 2972
rect 5080 2926 5132 2932
rect 5078 2816 5134 2825
rect 5078 2751 5134 2760
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5092 2553 5120 2751
rect 5078 2544 5134 2553
rect 5276 2514 5304 7296
rect 5368 5778 5396 14214
rect 5460 13410 5488 14554
rect 5460 13382 5580 13410
rect 5552 12866 5580 13382
rect 5460 12838 5580 12866
rect 5460 11830 5488 12838
rect 5644 12442 5672 16612
rect 5724 16594 5776 16600
rect 5828 15978 5856 19200
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16046 6132 16934
rect 6196 16250 6224 19200
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6380 16590 6408 17070
rect 6564 16980 6592 19200
rect 6472 16952 6592 16980
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15706 6224 15846
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5828 14362 5856 15302
rect 6012 15094 6040 15302
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5736 14334 5856 14362
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11082 5488 11494
rect 5540 11144 5592 11150
rect 5644 11132 5672 12378
rect 5592 11104 5672 11132
rect 5540 11086 5592 11092
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9042 5488 9318
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5460 8906 5488 8978
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5460 8362 5488 8842
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 7954 5488 8298
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5552 7698 5580 10678
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5644 7886 5672 9046
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5552 7670 5672 7698
rect 5644 6254 5672 7670
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5354 5400 5410 5409
rect 5460 5370 5488 5510
rect 5354 5335 5410 5344
rect 5448 5364 5500 5370
rect 5368 5001 5396 5335
rect 5448 5306 5500 5312
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5368 4078 5396 4927
rect 5460 4826 5488 5170
rect 5552 5166 5580 6122
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5644 4078 5672 6190
rect 5736 5098 5764 14334
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 11014 5856 14214
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5920 13326 5948 13874
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 5920 12714 5948 12922
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 6012 12434 6040 15030
rect 6196 15026 6224 15438
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5920 12406 6040 12434
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5828 8430 5856 8842
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6458 5856 6598
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5920 5846 5948 12406
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6012 11354 6040 12174
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6012 10810 6040 11290
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6012 9994 6040 10746
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6012 6798 6040 9114
rect 6104 7857 6132 12786
rect 6196 11558 6224 13738
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6288 12782 6316 13670
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6288 11642 6316 12718
rect 6380 12209 6408 16526
rect 6472 16454 6500 16952
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 6736 16720 6788 16726
rect 6734 16688 6736 16697
rect 6788 16688 6790 16697
rect 6734 16623 6790 16632
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6932 16250 6960 19200
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 7024 16658 7052 17002
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7208 16114 7236 16934
rect 7300 16697 7328 19200
rect 7668 17338 7696 19200
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7286 16688 7342 16697
rect 7286 16623 7342 16632
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7300 16250 7328 16390
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7392 16182 7420 16390
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7944 16130 7972 17002
rect 8036 16250 8064 19200
rect 8404 17524 8432 19200
rect 8312 17496 8432 17524
rect 8772 17524 8800 19200
rect 8772 17496 8892 17524
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 8312 16130 8340 17496
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8864 17338 8892 17496
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8404 16658 8432 16730
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8392 16176 8444 16182
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 7196 16108 7248 16114
rect 7248 16068 7328 16096
rect 7196 16050 7248 16056
rect 6472 13410 6500 16050
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6932 15473 6960 15642
rect 7208 15502 7236 15846
rect 7196 15496 7248 15502
rect 6918 15464 6974 15473
rect 7196 15438 7248 15444
rect 6918 15399 6974 15408
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6840 13938 6868 14350
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 7116 13818 7144 14350
rect 7024 13790 7144 13818
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 6472 13382 6592 13410
rect 6564 12753 6592 13382
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6550 12744 6606 12753
rect 6460 12708 6512 12714
rect 6840 12730 6868 12786
rect 6840 12702 6960 12730
rect 6550 12679 6606 12688
rect 6460 12650 6512 12656
rect 6366 12200 6422 12209
rect 6366 12135 6422 12144
rect 6472 12102 6500 12650
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6564 11830 6592 12174
rect 6932 12170 6960 12702
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6288 11614 6408 11642
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 10742 6224 11494
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6184 10736 6236 10742
rect 6184 10678 6236 10684
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 8090 6224 8842
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6090 7848 6146 7857
rect 6090 7783 6146 7792
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 7002 6132 7278
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5828 4078 5856 5714
rect 6012 5642 6040 6394
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6104 5778 6132 6326
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 5636 6052 5642
rect 6000 5578 6052 5584
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4622 5948 5102
rect 6012 5098 6040 5578
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 2514 5396 3334
rect 5460 2854 5488 3674
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5078 2479 5134 2488
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4618 2408 4674 2417
rect 4618 2343 4674 2352
rect 5356 2372 5408 2378
rect 4528 2032 4580 2038
rect 4528 1974 4580 1980
rect 4172 1686 4292 1714
rect 4264 800 4292 1686
rect 4540 800 4568 1974
rect 4632 1170 4660 2343
rect 5356 2314 5408 2320
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 4632 1142 4844 1170
rect 4816 800 4844 1142
rect 5092 800 5120 2042
rect 5368 800 5396 2314
rect 5644 800 5672 2858
rect 5736 2582 5764 3470
rect 6012 3194 6040 5034
rect 6104 4690 6132 5714
rect 6196 5166 6224 8026
rect 6288 7478 6316 11154
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6288 5778 6316 7414
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6380 5658 6408 11614
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11218 6500 11494
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6472 10810 6500 10950
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6472 9994 6500 10746
rect 6656 10713 6684 10950
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 9586 6684 9658
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9489 6684 9522
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 6736 8968 6788 8974
rect 6656 8928 6736 8956
rect 6656 8498 6684 8928
rect 6736 8910 6788 8916
rect 7024 8514 7052 13790
rect 7208 13530 7236 14962
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 10130 7144 13194
rect 7208 12434 7236 13466
rect 7300 13433 7328 16068
rect 7760 15910 7788 16118
rect 7944 16102 8064 16130
rect 8312 16124 8392 16130
rect 8312 16118 8444 16124
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 15094 7512 15302
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7286 13424 7342 13433
rect 7392 13394 7420 13874
rect 7286 13359 7342 13368
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 13320 7340 13326
rect 7286 13288 7288 13297
rect 7340 13288 7342 13297
rect 7286 13223 7342 13232
rect 7208 12406 7328 12434
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7102 10024 7158 10033
rect 7102 9959 7158 9968
rect 7116 9110 7144 9959
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9722 7236 9862
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6932 8486 7052 8514
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 6656 8362 6684 8434
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 6458 7440 6514 7449
rect 6458 7375 6514 7384
rect 6472 6798 6500 7375
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6288 5630 6408 5658
rect 6184 5160 6236 5166
rect 6288 5137 6316 5630
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6184 5102 6236 5108
rect 6274 5128 6330 5137
rect 6274 5063 6330 5072
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6288 4486 6316 5063
rect 6276 4480 6328 4486
rect 6196 4440 6276 4468
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5828 2446 5856 2790
rect 6012 2632 6040 3130
rect 6104 2990 6132 4082
rect 6196 3942 6224 4440
rect 6276 4422 6328 4428
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3194 6224 3878
rect 6288 3398 6316 4218
rect 6380 3534 6408 5510
rect 6736 5296 6788 5302
rect 6734 5264 6736 5273
rect 6788 5264 6790 5273
rect 6734 5199 6790 5208
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 6932 4758 6960 8486
rect 7116 7274 7144 8502
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 6390 7052 6666
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 5370 7144 6190
rect 7300 5778 7328 12406
rect 7484 11898 7512 15030
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7576 13297 7604 13466
rect 7562 13288 7618 13297
rect 7562 13223 7618 13232
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7576 11762 7604 11834
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7668 10470 7696 12650
rect 7760 11286 7788 15846
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7392 8090 7420 10066
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 6186 7420 8026
rect 7484 7002 7512 9590
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7668 6730 7696 10134
rect 7852 10010 7880 15982
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7944 14346 7972 14758
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12782 7972 13262
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7760 9982 7880 10010
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7484 5642 7512 6598
rect 7760 6458 7788 9982
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9382 7880 9522
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7944 8430 7972 10406
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8036 8378 8064 16102
rect 8116 16108 8168 16114
rect 8312 16102 8432 16118
rect 8168 16068 8248 16096
rect 8116 16050 8168 16056
rect 8220 16028 8248 16068
rect 8220 16000 8432 16028
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8128 12434 8156 15914
rect 8220 15609 8248 16000
rect 8404 15910 8432 16000
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8206 15600 8262 15609
rect 8206 15535 8262 15544
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15026 8248 15438
rect 8312 15434 8340 15846
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14346 8248 14962
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8220 13938 8248 14282
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8128 12406 8248 12434
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8128 11626 8156 12106
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8128 10266 8156 11562
rect 8220 11354 8248 12406
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11257 8340 15370
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8864 13258 8892 13874
rect 8956 13462 8984 14418
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8864 12918 8892 13194
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8956 12730 8984 13398
rect 8864 12702 8984 12730
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12481 8800 12582
rect 8758 12472 8814 12481
rect 8758 12407 8814 12416
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11286 8524 11698
rect 8484 11280 8536 11286
rect 8298 11248 8354 11257
rect 8208 11212 8260 11218
rect 8484 11222 8536 11228
rect 8298 11183 8354 11192
rect 8208 11154 8260 11160
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8036 8350 8156 8378
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7478 8064 8230
rect 8128 7750 8156 8350
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 7002 7880 7346
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7576 5642 7604 6054
rect 7668 5778 7696 6054
rect 7760 5914 7788 6394
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6920 4752 6972 4758
rect 6458 4720 6514 4729
rect 6920 4694 6972 4700
rect 6458 4655 6514 4664
rect 6472 3602 6500 4655
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 7024 3738 7052 5170
rect 7484 5166 7512 5578
rect 7562 5536 7618 5545
rect 7562 5471 7618 5480
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4282 7512 5102
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6380 3194 6408 3470
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 3194 6592 3334
rect 6840 3194 6868 3402
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6196 3058 6224 3130
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7010 2952 7066 2961
rect 6460 2848 6512 2854
rect 6196 2796 6460 2802
rect 6196 2790 6512 2796
rect 6196 2774 6500 2790
rect 6012 2604 6132 2632
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5920 800 5948 2518
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6012 2310 6040 2450
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6104 1426 6132 2604
rect 6092 1420 6144 1426
rect 6092 1362 6144 1368
rect 6196 800 6224 2774
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 6932 2530 6960 2926
rect 7010 2887 7066 2896
rect 6748 2502 6960 2530
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 6472 800 6500 1906
rect 6748 800 6776 2502
rect 7024 800 7052 2887
rect 7116 2514 7144 2994
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7208 2394 7236 4218
rect 7576 4185 7604 5471
rect 7760 4826 7788 5850
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7944 5681 7972 5714
rect 7930 5672 7986 5681
rect 7930 5607 7986 5616
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7654 4584 7710 4593
rect 7654 4519 7710 4528
rect 7668 4486 7696 4519
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7562 4176 7618 4185
rect 7562 4111 7618 4120
rect 7562 3632 7618 3641
rect 7392 3576 7562 3584
rect 7392 3556 7564 3576
rect 7392 2990 7420 3556
rect 7616 3567 7618 3576
rect 7564 3538 7616 3544
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7380 2984 7432 2990
rect 7564 2984 7616 2990
rect 7380 2926 7432 2932
rect 7484 2932 7564 2938
rect 7484 2926 7616 2932
rect 7300 2802 7328 2926
rect 7484 2910 7604 2926
rect 7484 2802 7512 2910
rect 7668 2836 7696 4422
rect 7760 3534 7788 4762
rect 7852 4690 7880 5510
rect 7930 5400 7986 5409
rect 7930 5335 7932 5344
rect 7984 5335 7986 5344
rect 7932 5306 7984 5312
rect 7944 4826 7972 5306
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 8036 4049 8064 6666
rect 8128 4758 8156 7686
rect 8220 6662 8248 11154
rect 8312 10470 8340 11183
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 8864 10742 8892 12702
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8298 10296 8354 10305
rect 8298 10231 8354 10240
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8312 6440 8340 10231
rect 8772 9908 8800 10610
rect 8772 9880 8892 9908
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8864 9178 8892 9880
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8864 8634 8892 8910
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8864 8498 8892 8570
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8864 8090 8892 8434
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 7002 8708 7142
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8864 6458 8892 6598
rect 8220 6412 8340 6440
rect 8852 6452 8904 6458
rect 8220 5234 8248 6412
rect 8852 6394 8904 6400
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8312 5370 8340 6258
rect 8864 5642 8892 6258
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8850 5400 8906 5409
rect 8300 5364 8352 5370
rect 8850 5335 8906 5344
rect 8300 5306 8352 5312
rect 8864 5234 8892 5335
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8864 5137 8892 5170
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8128 4282 8156 4694
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8114 4176 8170 4185
rect 8220 4162 8248 4762
rect 8404 4690 8432 4966
rect 8864 4826 8892 5063
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8760 4208 8812 4214
rect 8220 4134 8340 4162
rect 8760 4150 8812 4156
rect 8114 4111 8170 4120
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8036 3738 8064 3975
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8036 3602 8064 3674
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 3058 7972 3334
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7300 2774 7512 2802
rect 7576 2808 7696 2836
rect 7208 2366 7328 2394
rect 7300 800 7328 2366
rect 7576 800 7604 2808
rect 7944 2774 7972 2994
rect 7944 2746 8064 2774
rect 8036 2582 8064 2746
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 7852 800 7880 1362
rect 8128 800 8156 4111
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3602 8248 4014
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8220 2378 8248 2994
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8312 1986 8340 4134
rect 8772 3738 8800 4150
rect 8956 3924 8984 12174
rect 9048 12170 9076 16594
rect 9140 16522 9168 19200
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9416 16658 9444 16730
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9218 16280 9274 16289
rect 9218 16215 9274 16224
rect 9126 16144 9182 16153
rect 9126 16079 9182 16088
rect 9140 14074 9168 16079
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9126 12472 9182 12481
rect 9126 12407 9182 12416
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 9042 9076 12106
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9140 7886 9168 12407
rect 9232 10266 9260 16215
rect 9324 16046 9352 16390
rect 9416 16289 9444 16594
rect 9402 16280 9458 16289
rect 9402 16215 9458 16224
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14618 9352 14758
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9324 13938 9352 14554
rect 9416 14521 9444 16050
rect 9508 15978 9536 19200
rect 9876 17082 9904 19200
rect 10048 17128 10100 17134
rect 9876 17054 9996 17082
rect 10048 17070 10100 17076
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9600 16590 9628 16730
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9876 16454 9904 16934
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9692 16114 9720 16186
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9692 15910 9720 16050
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9508 14618 9536 15370
rect 9784 14906 9812 15846
rect 9876 15178 9904 16390
rect 9968 16250 9996 17054
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10060 15314 10088 17070
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16250 10180 16390
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 15416 10272 19200
rect 10612 16998 10640 19200
rect 10980 17066 11008 19200
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 15910 10364 16050
rect 10324 15904 10376 15910
rect 10612 15892 10640 16390
rect 10612 15864 10732 15892
rect 10324 15846 10376 15852
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10704 15706 10732 15864
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10244 15388 10364 15416
rect 10060 15286 10272 15314
rect 9876 15150 10180 15178
rect 9784 14878 9996 14906
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9402 14512 9458 14521
rect 9402 14447 9458 14456
rect 9508 14074 9536 14554
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9416 12238 9444 14010
rect 9496 12640 9548 12646
rect 9494 12608 9496 12617
rect 9548 12608 9550 12617
rect 9494 12543 9550 12552
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9600 11778 9628 14282
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9324 11750 9628 11778
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9232 9994 9260 10202
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9324 9704 9352 11750
rect 9692 11694 9720 12038
rect 9496 11688 9548 11694
rect 9402 11656 9458 11665
rect 9680 11688 9732 11694
rect 9496 11630 9548 11636
rect 9600 11648 9680 11676
rect 9402 11591 9458 11600
rect 9416 10674 9444 11591
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9508 10470 9536 11630
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9232 9676 9352 9704
rect 9232 9500 9260 9676
rect 9508 9674 9536 10406
rect 9600 9897 9628 11648
rect 9680 11630 9732 11636
rect 9692 11565 9720 11630
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 9926 9720 11018
rect 9784 10538 9812 13738
rect 9876 13326 9904 14214
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9968 12434 9996 14878
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9876 12406 9996 12434
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9680 9920 9732 9926
rect 9586 9888 9642 9897
rect 9680 9862 9732 9868
rect 9586 9823 9642 9832
rect 9692 9722 9720 9862
rect 9680 9716 9732 9722
rect 9508 9646 9597 9674
rect 9680 9658 9732 9664
rect 9569 9500 9597 9646
rect 9678 9616 9734 9625
rect 9678 9551 9734 9560
rect 9232 9472 9352 9500
rect 9324 9382 9352 9472
rect 9508 9472 9597 9500
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9048 6254 9076 7822
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9048 5166 9076 6190
rect 9140 5817 9168 7414
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6798 9260 7142
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9126 5808 9182 5817
rect 9126 5743 9182 5752
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9048 4486 9076 4558
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 9140 4078 9168 5646
rect 9232 5574 9260 6734
rect 9324 6633 9352 9318
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9310 6624 9366 6633
rect 9310 6559 9366 6568
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9324 6254 9352 6394
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9416 6089 9444 7958
rect 9402 6080 9458 6089
rect 9402 6015 9458 6024
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9402 5808 9458 5817
rect 9508 5778 9536 9472
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9042 9628 9318
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9692 8090 9720 9551
rect 9784 8906 9812 10474
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9600 5953 9628 6394
rect 9586 5944 9642 5953
rect 9784 5914 9812 7754
rect 9586 5879 9642 5888
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9586 5808 9642 5817
rect 9402 5743 9458 5752
rect 9496 5772 9548 5778
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4690 9260 5510
rect 9324 5302 9352 5607
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9324 5030 9352 5238
rect 9416 5166 9444 5743
rect 9586 5743 9642 5752
rect 9496 5714 9548 5720
rect 9600 5710 9628 5743
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9600 4622 9628 5238
rect 9784 5166 9812 5510
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9876 5012 9904 12406
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9968 8634 9996 12106
rect 10060 11937 10088 13194
rect 10152 12986 10180 15150
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10046 11928 10102 11937
rect 10046 11863 10102 11872
rect 10152 11744 10180 12786
rect 10244 11830 10272 15286
rect 10336 15094 10364 15388
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10598 14376 10654 14385
rect 10598 14311 10654 14320
rect 10612 13716 10640 14311
rect 10704 14278 10732 14962
rect 10692 14272 10744 14278
rect 10690 14240 10692 14249
rect 10744 14240 10746 14249
rect 10690 14175 10746 14184
rect 10612 13688 10732 13716
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10322 11928 10378 11937
rect 10322 11863 10378 11872
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10060 11716 10180 11744
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10060 8430 10088 11716
rect 10336 11676 10364 11863
rect 10244 11648 10364 11676
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10152 9994 10180 11290
rect 10244 10810 10272 11648
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10060 7188 10088 8366
rect 10140 7200 10192 7206
rect 10060 7160 10140 7188
rect 10140 7142 10192 7148
rect 10244 7002 10272 10610
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 9654 10548 9862
rect 10704 9674 10732 13688
rect 10796 12442 10824 16526
rect 11348 15609 11376 19200
rect 11334 15600 11390 15609
rect 11334 15535 11390 15544
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10888 13326 10916 14962
rect 10980 14890 11008 15302
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11060 13864 11112 13870
rect 11058 13832 11060 13841
rect 11112 13832 11114 13841
rect 11058 13767 11114 13776
rect 11060 13456 11112 13462
rect 11058 13424 11060 13433
rect 11112 13424 11114 13433
rect 11058 13359 11114 13368
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10888 12782 10916 13262
rect 11072 13190 11100 13359
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11164 12782 11192 13874
rect 11348 13394 11376 15438
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 11150 10824 12378
rect 10888 12306 10916 12718
rect 10966 12472 11022 12481
rect 10966 12407 11022 12416
rect 10980 12322 11008 12407
rect 11164 12374 11192 12718
rect 11152 12368 11204 12374
rect 10876 12300 10928 12306
rect 10980 12294 11100 12322
rect 11152 12310 11204 12316
rect 10876 12242 10928 12248
rect 10888 11218 10916 12242
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10888 10674 10916 11154
rect 10980 10962 11008 11766
rect 11072 11354 11100 12294
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10980 10934 11100 10962
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10130 10916 10610
rect 10980 10130 11008 10746
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 10033 11008 10066
rect 10966 10024 11022 10033
rect 10966 9959 11022 9968
rect 10508 9648 10560 9654
rect 10704 9646 10824 9674
rect 10508 9590 10560 9596
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9876 4984 9996 5012
rect 9862 4856 9918 4865
rect 9862 4791 9864 4800
rect 9916 4791 9918 4800
rect 9864 4762 9916 4768
rect 9876 4622 9904 4762
rect 9588 4616 9640 4622
rect 9586 4584 9588 4593
rect 9864 4616 9916 4622
rect 9640 4584 9642 4593
rect 9586 4519 9642 4528
rect 9784 4564 9864 4570
rect 9784 4558 9916 4564
rect 9784 4542 9904 4558
rect 9600 4493 9628 4519
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9324 4146 9352 4247
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9404 3936 9456 3942
rect 8956 3896 9404 3924
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8446 3292 8754 3301
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8496 2514 8524 2994
rect 8942 2544 8998 2553
rect 8484 2508 8536 2514
rect 8942 2479 8998 2488
rect 8484 2450 8536 2456
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8666 2000 8722 2009
rect 8312 1958 8432 1986
rect 8404 800 8432 1958
rect 8666 1935 8722 1944
rect 8680 800 8708 1935
rect 8956 800 8984 2479
rect 9036 2440 9088 2446
rect 9088 2388 9168 2394
rect 9036 2382 9168 2388
rect 9048 2366 9168 2382
rect 9140 2310 9168 2366
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9232 800 9260 3896
rect 9404 3878 9456 3884
rect 9310 3768 9366 3777
rect 9310 3703 9312 3712
rect 9364 3703 9366 3712
rect 9588 3732 9640 3738
rect 9312 3674 9364 3680
rect 9588 3674 9640 3680
rect 9324 2446 9352 3674
rect 9600 3466 9628 3674
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9692 3369 9720 3606
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9508 2514 9536 2994
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2582 9720 2926
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9692 2310 9720 2518
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9494 1864 9550 1873
rect 9494 1799 9550 1808
rect 9508 800 9536 1799
rect 9784 800 9812 4542
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9876 4010 9904 4422
rect 9968 4282 9996 4984
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10060 4078 10088 6122
rect 10244 5760 10272 6938
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10324 5772 10376 5778
rect 10244 5732 10324 5760
rect 10796 5760 10824 9646
rect 11072 9625 11100 10934
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10324 5714 10376 5720
rect 10704 5732 10824 5760
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 10520 5370 10548 5471
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10152 5098 10180 5238
rect 10520 5234 10548 5306
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9876 1902 9904 3946
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9968 3398 9996 3606
rect 10060 3602 10088 4014
rect 10152 3738 10180 4150
rect 10336 3924 10364 4694
rect 10704 4146 10732 5732
rect 10980 5658 11008 9046
rect 11072 8974 11100 9454
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 7954 11100 8910
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 6458 11100 7754
rect 11164 6746 11192 11698
rect 11256 11014 11284 12786
rect 11348 12306 11376 13330
rect 11440 13258 11468 19230
rect 11624 19122 11652 19230
rect 11702 19200 11758 20000
rect 11808 19230 12020 19258
rect 11716 19122 11744 19200
rect 11624 19094 11744 19122
rect 11518 16280 11574 16289
rect 11808 16266 11836 19230
rect 11992 19122 12020 19230
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 14752 19230 14964 19258
rect 12084 19122 12112 19200
rect 11992 19094 12112 19122
rect 12072 17536 12124 17542
rect 12452 17524 12480 19200
rect 12452 17496 12572 17524
rect 12072 17478 12124 17484
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11518 16215 11574 16224
rect 11624 16238 11836 16266
rect 11992 16250 12020 17274
rect 12084 17270 12112 17478
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11980 16244 12032 16250
rect 11532 16046 11560 16215
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 13954 11560 15846
rect 11624 14074 11652 16238
rect 11980 16186 12032 16192
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11716 15638 11744 16050
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11808 15094 11836 15846
rect 11900 15570 11928 16050
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11992 15094 12020 15914
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11900 14482 11928 14894
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 12084 14362 12112 16594
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12176 15502 12204 16050
rect 12268 15706 12296 16118
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12360 15348 12388 15982
rect 12452 15745 12480 16186
rect 12544 15910 12572 17496
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12636 16998 12664 17070
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12438 15736 12494 15745
rect 12438 15671 12440 15680
rect 12492 15671 12494 15680
rect 12440 15642 12492 15648
rect 12360 15320 12572 15348
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12438 14648 12494 14657
rect 12438 14583 12494 14592
rect 12452 14385 12480 14583
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11992 14334 12112 14362
rect 12438 14376 12494 14385
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11532 13926 11652 13954
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13394 11560 13670
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11624 13274 11652 13926
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11532 13246 11652 13274
rect 11704 13252 11756 13258
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11440 12481 11468 12922
rect 11426 12472 11482 12481
rect 11426 12407 11482 12416
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11532 11762 11560 13246
rect 11704 13194 11756 13200
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11624 11694 11652 13126
rect 11716 12986 11744 13194
rect 11808 13190 11836 13738
rect 11900 13530 11928 14282
rect 11992 13530 12020 14334
rect 12438 14311 12494 14320
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11440 11234 11468 11494
rect 11532 11354 11560 11562
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11440 11206 11560 11234
rect 11624 11218 11652 11630
rect 11532 11098 11560 11206
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11428 11076 11480 11082
rect 11532 11070 11652 11098
rect 11428 11018 11480 11024
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11440 10266 11468 11018
rect 11518 10976 11574 10985
rect 11518 10911 11574 10920
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 7954 11284 8910
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7478 11284 7686
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11164 6718 11284 6746
rect 11150 6624 11206 6633
rect 11150 6559 11206 6568
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10784 5636 10836 5642
rect 10980 5630 11100 5658
rect 10784 5578 10836 5584
rect 10796 4758 10824 5578
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10888 4826 10916 5510
rect 10980 5370 11008 5510
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11072 5114 11100 5630
rect 10980 5086 11100 5114
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10980 4434 11008 5086
rect 10888 4406 11008 4434
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10244 3896 10364 3924
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10138 3632 10194 3641
rect 10048 3596 10100 3602
rect 10138 3567 10194 3576
rect 10048 3538 10100 3544
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3194 9996 3334
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 2038 9996 2246
rect 9956 2032 10008 2038
rect 9956 1974 10008 1980
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 10060 800 10088 3402
rect 10152 2258 10180 3567
rect 10244 3534 10272 3896
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10704 3398 10732 4082
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 3058 10732 3334
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10244 2446 10272 2994
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10704 2530 10732 2790
rect 10796 2650 10824 4150
rect 10888 3670 10916 4406
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10980 3738 11008 4218
rect 11164 4128 11192 6559
rect 11256 6322 11284 6718
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11348 5896 11376 8230
rect 11440 6798 11468 8774
rect 11532 8634 11560 10911
rect 11624 10266 11652 11070
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11716 9602 11744 12922
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11808 11354 11836 12106
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11992 10810 12020 13126
rect 12084 12442 12112 14214
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12268 13190 12296 14010
rect 12544 13938 12572 15320
rect 12636 15144 12664 16934
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12728 15706 12756 16662
rect 12820 15745 12848 19200
rect 13188 16946 13216 19200
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13188 16918 13308 16946
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12806 15736 12862 15745
rect 12716 15700 12768 15706
rect 12806 15671 12862 15680
rect 12716 15642 12768 15648
rect 12636 15116 12848 15144
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12636 14006 12664 14758
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12268 12306 12296 12582
rect 12728 12434 12756 14758
rect 12820 14362 12848 15116
rect 12912 14550 12940 16526
rect 13004 15570 13032 16594
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12820 14334 12940 14362
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 14074 12848 14214
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12912 13326 12940 14334
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12544 12406 12756 12434
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12254 12200 12310 12209
rect 12254 12135 12256 12144
rect 12308 12135 12310 12144
rect 12256 12106 12308 12112
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11898 12112 12038
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11624 9574 11744 9602
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 8090 11652 9574
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11716 8566 11744 9386
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11624 7342 11652 8026
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 6866 11560 7142
rect 11610 7032 11666 7041
rect 11610 6967 11666 6976
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11426 6352 11482 6361
rect 11426 6287 11482 6296
rect 11440 6254 11468 6287
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11348 5868 11468 5896
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11242 4856 11298 4865
rect 11242 4791 11298 4800
rect 11256 4622 11284 4791
rect 11348 4690 11376 5714
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4282 11284 4422
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11164 4100 11284 4128
rect 11256 4010 11284 4100
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11072 3670 11100 3878
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11256 3602 11284 3946
rect 11336 3936 11388 3942
rect 11334 3904 11336 3913
rect 11388 3904 11390 3913
rect 11334 3839 11390 3848
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11060 3528 11112 3534
rect 10874 3496 10930 3505
rect 11060 3470 11112 3476
rect 10874 3431 10930 3440
rect 10888 3233 10916 3431
rect 10874 3224 10930 3233
rect 10874 3159 10876 3168
rect 10928 3159 10930 3168
rect 10876 3130 10928 3136
rect 10888 3099 10916 3130
rect 11072 2990 11100 3470
rect 11336 3392 11388 3398
rect 11242 3360 11298 3369
rect 11336 3334 11388 3340
rect 11242 3295 11298 3304
rect 11256 3194 11284 3295
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11256 3058 11284 3130
rect 11348 3097 11376 3334
rect 11334 3088 11390 3097
rect 11244 3052 11296 3058
rect 11164 3012 11244 3040
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2774 11100 2926
rect 10888 2746 11100 2774
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10612 2502 10732 2530
rect 10796 2514 10824 2586
rect 10784 2508 10836 2514
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10152 2230 10364 2258
rect 10336 800 10364 2230
rect 10612 800 10640 2502
rect 10784 2450 10836 2456
rect 10888 800 10916 2746
rect 11164 800 11192 3012
rect 11334 3023 11390 3032
rect 11244 2994 11296 3000
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 1494 11284 2246
rect 11244 1488 11296 1494
rect 11244 1430 11296 1436
rect 11440 800 11468 5868
rect 11532 5778 11560 6598
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11624 5642 11652 6967
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11624 5370 11652 5578
rect 11612 5364 11664 5370
rect 11532 5324 11612 5352
rect 11532 2922 11560 5324
rect 11612 5306 11664 5312
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11624 4729 11652 5170
rect 11610 4720 11666 4729
rect 11610 4655 11666 4664
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11532 2650 11560 2751
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11624 1698 11652 4422
rect 11716 3942 11744 6054
rect 11808 5846 11836 9862
rect 11900 6662 11928 9862
rect 12084 9674 12112 11018
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12360 10266 12388 10746
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 11992 9646 12112 9674
rect 11992 9217 12020 9646
rect 12544 9518 12572 12406
rect 13004 12238 13032 15506
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14618 13124 14894
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13188 14074 13216 16730
rect 13280 15144 13308 16918
rect 13372 16726 13400 17070
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15502 13400 16390
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13280 15116 13400 15144
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14618 13308 14962
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13268 14272 13320 14278
rect 13266 14240 13268 14249
rect 13320 14240 13322 14249
rect 13266 14175 13322 14184
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11150 13032 12038
rect 13096 11354 13124 13942
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11978 9208 12034 9217
rect 11978 9143 12034 9152
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11992 7478 12020 8978
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 12084 7002 12112 9318
rect 12544 8974 12572 9454
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8537 12480 8570
rect 12438 8528 12494 8537
rect 12438 8463 12494 8472
rect 12452 7818 12480 8463
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11900 5522 11928 6054
rect 12084 5914 12112 6598
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12346 6352 12402 6361
rect 12452 6322 12480 6394
rect 12346 6287 12402 6296
rect 12440 6316 12492 6322
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12360 5778 12388 6287
rect 12440 6258 12492 6264
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12070 5672 12126 5681
rect 12070 5607 12072 5616
rect 12124 5607 12126 5616
rect 12072 5578 12124 5584
rect 11808 5494 11928 5522
rect 11808 5250 11836 5494
rect 11886 5400 11942 5409
rect 12084 5370 12112 5578
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12072 5364 12124 5370
rect 11942 5344 12020 5352
rect 11886 5335 11888 5344
rect 11940 5324 12020 5344
rect 11888 5306 11940 5312
rect 11808 5222 11928 5250
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11808 4078 11836 5102
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11704 3936 11756 3942
rect 11756 3896 11836 3924
rect 11704 3878 11756 3884
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 1692 11664 1698
rect 11612 1634 11664 1640
rect 11716 800 11744 3674
rect 11808 2774 11836 3896
rect 11900 3618 11928 5222
rect 11992 5030 12020 5324
rect 12072 5306 12124 5312
rect 12438 5264 12494 5273
rect 12072 5228 12124 5234
rect 12438 5199 12494 5208
rect 12072 5170 12124 5176
rect 12084 5098 12112 5170
rect 12162 5128 12218 5137
rect 12072 5092 12124 5098
rect 12162 5063 12218 5072
rect 12072 5034 12124 5040
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11992 4146 12020 4694
rect 12176 4690 12204 5063
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12452 4486 12480 5199
rect 12544 4842 12572 8910
rect 12636 7546 12664 10950
rect 13096 10810 13124 10950
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13188 10146 13216 11834
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 13096 10118 13216 10146
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9722 12756 9862
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12912 9654 12940 10066
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9722 13032 9862
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12900 9648 12952 9654
rect 13004 9625 13032 9658
rect 12900 9590 12952 9596
rect 12990 9616 13046 9625
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 6798 12756 9386
rect 12912 9042 12940 9590
rect 12990 9551 13046 9560
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12990 8936 13046 8945
rect 12990 8871 13046 8880
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8634 12848 8774
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 8090 12940 8434
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6322 12664 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12728 6118 12756 6394
rect 12820 6322 12848 7754
rect 12912 7342 12940 7890
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5953 12848 6054
rect 12806 5944 12862 5953
rect 12806 5879 12862 5888
rect 12714 5672 12770 5681
rect 12714 5607 12770 5616
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5030 12664 5510
rect 12728 5370 12756 5607
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12544 4814 12664 4842
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12084 3738 12112 4422
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12176 3942 12204 4150
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12452 3738 12480 4082
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11900 3590 12112 3618
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3194 12020 3334
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11808 2746 12020 2774
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11808 2106 11836 2246
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11900 1970 11928 2246
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11992 800 12020 2746
rect 12084 1986 12112 3590
rect 12452 3534 12480 3674
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12348 3120 12400 3126
rect 12162 3088 12218 3097
rect 12348 3062 12400 3068
rect 12162 3023 12218 3032
rect 12176 2825 12204 3023
rect 12360 2922 12388 3062
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12162 2816 12218 2825
rect 12162 2751 12218 2760
rect 12360 2650 12388 2858
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12452 2378 12480 2994
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12084 1958 12296 1986
rect 12268 800 12296 1958
rect 12544 800 12572 4694
rect 12636 2514 12664 4814
rect 12728 4672 12756 5306
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12820 4865 12848 5034
rect 12806 4856 12862 4865
rect 12806 4791 12862 4800
rect 12728 4644 12848 4672
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 4282 12756 4490
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12728 3777 12756 3878
rect 12714 3768 12770 3777
rect 12714 3703 12716 3712
rect 12768 3703 12770 3712
rect 12716 3674 12768 3680
rect 12728 2990 12756 3674
rect 12820 3097 12848 4644
rect 12912 4622 12940 6598
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12806 3088 12862 3097
rect 12806 3023 12862 3032
rect 12716 2984 12768 2990
rect 13004 2938 13032 8871
rect 13096 8838 13124 10118
rect 13176 9988 13228 9994
rect 13176 9930 13228 9936
rect 13188 9722 13216 9930
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13280 8650 13308 14010
rect 13372 13530 13400 15116
rect 13464 15094 13492 16594
rect 13556 15162 13584 19200
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13648 16289 13676 17002
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15570 13676 16050
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13464 13938 13492 14486
rect 13556 14260 13584 15098
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13648 14498 13676 15030
rect 13740 14657 13768 16186
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13832 14822 13860 15642
rect 13924 15609 13952 19200
rect 14292 17082 14320 19200
rect 14660 19122 14688 19200
rect 14752 19122 14780 19230
rect 14660 19094 14780 19122
rect 14292 17054 14504 17082
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14476 16182 14504 17054
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16658 14596 17002
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14752 16454 14780 16934
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14464 16176 14516 16182
rect 14278 16144 14334 16153
rect 14464 16118 14516 16124
rect 14278 16079 14280 16088
rect 14332 16079 14334 16088
rect 14280 16050 14332 16056
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 14476 15706 14504 16118
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 13910 15600 13966 15609
rect 13910 15535 13966 15544
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13726 14648 13782 14657
rect 13726 14583 13782 14592
rect 13648 14470 13768 14498
rect 13556 14232 13676 14260
rect 13542 14104 13598 14113
rect 13648 14074 13676 14232
rect 13542 14039 13598 14048
rect 13636 14068 13688 14074
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12850 13400 13330
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13372 10606 13400 12242
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 9654 13400 10542
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13096 8622 13308 8650
rect 13096 6866 13124 8622
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 13188 7546 13216 8502
rect 13372 8430 13400 9590
rect 13464 9586 13492 13874
rect 13556 12986 13584 14039
rect 13636 14010 13688 14016
rect 13740 13734 13768 14470
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13648 13190 13676 13466
rect 13740 13394 13768 13670
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13556 9994 13584 12718
rect 13648 12102 13676 13126
rect 13832 12986 13860 14282
rect 13924 14074 13952 15370
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 13924 13190 13952 13874
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 14094 13424 14150 13433
rect 14094 13359 14096 13368
rect 14148 13359 14150 13368
rect 14096 13330 14148 13336
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13924 12866 13952 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13832 12838 13952 12866
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11898 13676 12038
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13634 11792 13690 11801
rect 13634 11727 13636 11736
rect 13688 11727 13690 11736
rect 13636 11698 13688 11704
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 10742 13676 11494
rect 13740 11354 13768 12786
rect 13832 11830 13860 12838
rect 13910 12744 13966 12753
rect 13910 12679 13966 12688
rect 13924 12442 13952 12679
rect 14016 12646 14044 13262
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13726 11112 13782 11121
rect 13726 11047 13782 11056
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13740 9602 13768 11047
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13832 10130 13860 10678
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13648 9574 13768 9602
rect 13464 9110 13492 9522
rect 13648 9518 13676 9574
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9382 13676 9454
rect 13820 9444 13872 9450
rect 13740 9404 13820 9432
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13740 9110 13768 9404
rect 13820 9386 13872 9392
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13464 8106 13492 9046
rect 13740 8906 13768 9046
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13820 8832 13872 8838
rect 13924 8809 13952 12174
rect 14108 12170 14136 12378
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14002 11792 14058 11801
rect 14002 11727 14004 11736
rect 14056 11727 14058 11736
rect 14004 11698 14056 11704
rect 14200 11694 14228 12310
rect 14476 11778 14504 13874
rect 14568 13530 14596 14214
rect 14660 14006 14688 14962
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14752 13682 14780 16390
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14660 13654 14780 13682
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14660 13161 14688 13654
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14646 13152 14702 13161
rect 14646 13087 14702 13096
rect 14752 12918 14780 13330
rect 14844 13190 14872 15574
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14740 12776 14792 12782
rect 14792 12736 14872 12764
rect 14740 12718 14792 12724
rect 14844 12442 14872 12736
rect 14936 12442 14964 19230
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16854 19200 16910 20000
rect 15028 15858 15056 19200
rect 15108 16584 15160 16590
rect 15106 16552 15108 16561
rect 15160 16552 15162 16561
rect 15106 16487 15162 16496
rect 15028 15830 15148 15858
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 14074 15056 14758
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12850 15056 13126
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 12753 15056 12786
rect 15014 12744 15070 12753
rect 15014 12679 15070 12688
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14830 12336 14886 12345
rect 15028 12288 15056 12582
rect 14830 12271 14886 12280
rect 14384 11750 14504 11778
rect 14556 11756 14608 11762
rect 14188 11688 14240 11694
rect 14384 11665 14412 11750
rect 14556 11698 14608 11704
rect 14464 11688 14516 11694
rect 14188 11630 14240 11636
rect 14370 11656 14426 11665
rect 14464 11630 14516 11636
rect 14370 11591 14426 11600
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 14096 11280 14148 11286
rect 14372 11280 14424 11286
rect 14096 11222 14148 11228
rect 14186 11248 14242 11257
rect 14108 10810 14136 11222
rect 14186 11183 14242 11192
rect 14370 11248 14372 11257
rect 14424 11248 14426 11257
rect 14370 11183 14426 11192
rect 14200 11082 14228 11183
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10810 14412 10950
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14384 10452 14412 10746
rect 14476 10606 14504 11630
rect 14568 11014 14596 11698
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14384 10424 14504 10452
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10299 14376 10308
rect 14002 10160 14058 10169
rect 14476 10130 14504 10424
rect 14568 10266 14596 10678
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14002 10095 14058 10104
rect 14464 10124 14516 10130
rect 14016 9625 14044 10095
rect 14464 10066 14516 10072
rect 14476 9674 14504 10066
rect 14384 9646 14504 9674
rect 14002 9616 14058 9625
rect 14002 9551 14058 9560
rect 14384 9489 14412 9646
rect 14370 9480 14426 9489
rect 14370 9415 14426 9424
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 13820 8774 13872 8780
rect 13910 8800 13966 8809
rect 13372 8078 13492 8106
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13084 6860 13136 6866
rect 13136 6820 13216 6848
rect 13084 6802 13136 6808
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 4758 13124 6598
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13188 4214 13216 6820
rect 13280 5914 13308 7686
rect 13372 6798 13400 8078
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7274 13492 7890
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7546 13584 7686
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13648 7426 13676 8774
rect 13832 7478 13860 8774
rect 13910 8735 13966 8744
rect 14002 8664 14058 8673
rect 14002 8599 14004 8608
rect 14056 8599 14058 8608
rect 14004 8570 14056 8576
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13556 7398 13676 7426
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6458 13400 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13556 6338 13584 7398
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13648 7002 13676 7278
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13924 6866 13952 8502
rect 14016 8294 14044 8570
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14292 7546 14320 7754
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13372 6310 13584 6338
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5760 13400 6310
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13280 5732 13400 5760
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 13280 4146 13308 5732
rect 13358 5672 13414 5681
rect 13358 5607 13360 5616
rect 13412 5607 13414 5616
rect 13360 5578 13412 5584
rect 13464 5370 13492 6190
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5710 13584 6054
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13452 5160 13504 5166
rect 13372 5120 13452 5148
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13280 3194 13308 3674
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 12716 2926 12768 2932
rect 12820 2910 13032 2938
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12820 800 12848 2910
rect 13096 2774 13124 3062
rect 13372 2774 13400 5120
rect 13556 5148 13584 5238
rect 13504 5120 13584 5148
rect 13636 5160 13688 5166
rect 13452 5102 13504 5108
rect 13636 5102 13688 5108
rect 13648 4826 13676 5102
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13648 3738 13676 4762
rect 13740 4146 13768 6122
rect 13832 5846 13860 6802
rect 13924 5896 13952 6802
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 14016 6458 14044 6666
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14016 6254 14044 6394
rect 14108 6254 14136 6802
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 13924 5868 14044 5896
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13910 5808 13966 5817
rect 13832 4690 13860 5782
rect 13910 5743 13966 5752
rect 13924 5574 13952 5743
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13924 5370 13952 5510
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 14016 4978 14044 5868
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14384 5370 14412 5646
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14280 5228 14332 5234
rect 14384 5216 14412 5306
rect 14476 5250 14504 9318
rect 14568 8974 14596 9318
rect 14660 9178 14688 10610
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10062 14780 10406
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14738 9888 14794 9897
rect 14738 9823 14794 9832
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14752 9024 14780 9823
rect 14660 8996 14780 9024
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14660 7562 14688 8996
rect 14738 8936 14794 8945
rect 14738 8871 14794 8880
rect 14752 8430 14780 8871
rect 14844 8566 14872 12271
rect 14936 12260 15056 12288
rect 14936 8922 14964 12260
rect 15120 12186 15148 15830
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 13394 15240 14418
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15304 13394 15332 14214
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15212 13240 15240 13330
rect 15396 13326 15424 19200
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15212 13212 15332 13240
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15212 12434 15240 12922
rect 15304 12782 15332 13212
rect 15396 12986 15424 13262
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15212 12406 15424 12434
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15028 12158 15148 12186
rect 15028 9450 15056 12158
rect 15212 11626 15240 12242
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15212 11218 15240 11562
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 10124 15160 10130
rect 15212 10112 15240 11154
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15160 10084 15240 10112
rect 15108 10066 15160 10072
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15120 9110 15148 9959
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 14936 8894 15148 8922
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8634 14964 8774
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14568 7534 14688 7562
rect 14568 6662 14596 7534
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14660 7002 14688 7346
rect 14844 7342 14872 7890
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6390 14688 6802
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14660 5778 14688 6326
rect 14752 5914 14780 7278
rect 14844 6866 14872 7278
rect 15120 7002 15148 8894
rect 15212 8634 15240 9590
rect 15304 9178 15332 11086
rect 15396 9382 15424 12406
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15290 8936 15346 8945
rect 15290 8871 15292 8880
rect 15344 8871 15346 8880
rect 15292 8842 15344 8848
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15212 7546 15240 7686
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 15016 6792 15068 6798
rect 14830 6760 14886 6769
rect 15016 6734 15068 6740
rect 14830 6695 14886 6704
rect 14844 6662 14872 6695
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6118 14872 6598
rect 15028 6474 15056 6734
rect 14936 6446 15056 6474
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5370 14596 5510
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14476 5222 14596 5250
rect 14332 5188 14412 5216
rect 14280 5170 14332 5176
rect 13924 4950 14044 4978
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13726 3904 13782 3913
rect 13726 3839 13782 3848
rect 13740 3738 13768 3839
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13832 3534 13860 3946
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13924 3380 13952 4950
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14384 4078 14412 4655
rect 14568 4622 14596 5222
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4298 14596 4558
rect 14568 4270 14688 4298
rect 14660 4214 14688 4270
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 14476 3738 14504 4150
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13832 3352 13952 3380
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 12912 2746 13124 2774
rect 13280 2746 13400 2774
rect 12912 2650 12940 2746
rect 13280 2650 13308 2746
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12912 2310 12940 2586
rect 13280 2446 13308 2586
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13084 1828 13136 1834
rect 13084 1770 13136 1776
rect 13096 800 13124 1770
rect 13372 800 13400 2586
rect 13464 2310 13492 2994
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13740 2650 13768 2790
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13464 1834 13492 2246
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13648 800 13676 2450
rect 13832 2446 13860 3352
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13924 1578 13952 2926
rect 14016 2922 14044 3538
rect 14568 3398 14596 4014
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14464 3120 14516 3126
rect 14186 3088 14242 3097
rect 14464 3062 14516 3068
rect 14186 3023 14188 3032
rect 14240 3023 14242 3032
rect 14188 2994 14240 3000
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 14186 2408 14242 2417
rect 14186 2343 14242 2352
rect 14200 2310 14228 2343
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 13924 1550 14228 1578
rect 13912 1488 13964 1494
rect 13912 1430 13964 1436
rect 13924 800 13952 1430
rect 14200 800 14228 1550
rect 14476 800 14504 3062
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14568 2650 14596 2994
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14660 2394 14688 4150
rect 14752 3194 14780 5170
rect 14844 4146 14872 6054
rect 14936 4729 14964 6446
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15028 5234 15056 5306
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14922 4720 14978 4729
rect 15120 4690 15148 6190
rect 15212 5302 15240 7482
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 6798 15332 7142
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15290 6488 15346 6497
rect 15290 6423 15292 6432
rect 15344 6423 15346 6432
rect 15292 6394 15344 6400
rect 15304 5574 15332 6394
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15292 5160 15344 5166
rect 15396 5148 15424 9318
rect 15488 9110 15516 14282
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 6866 15516 8910
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15488 5778 15516 6802
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15488 5302 15516 5714
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 15396 5120 15516 5148
rect 15292 5102 15344 5108
rect 14922 4655 14978 4664
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3602 14872 3878
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 15120 3534 15148 4626
rect 15304 4622 15332 5102
rect 15292 4616 15344 4622
rect 15198 4584 15254 4593
rect 15292 4558 15344 4564
rect 15198 4519 15254 4528
rect 15212 4282 15240 4519
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15212 3602 15240 4218
rect 15488 4146 15516 5120
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14568 2378 14688 2394
rect 14556 2372 14688 2378
rect 14608 2366 14688 2372
rect 14556 2314 14608 2320
rect 14752 800 14780 2858
rect 15304 2582 15332 3878
rect 15488 3738 15516 4082
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3074 15608 17138
rect 15764 16250 15792 19200
rect 16132 17134 16160 19200
rect 16500 17338 16528 19200
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15672 14414 15700 15098
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15672 7206 15700 10950
rect 15764 10810 15792 14010
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15764 5710 15792 9930
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15488 3058 15608 3074
rect 15672 3058 15700 4558
rect 15764 3738 15792 5646
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15764 3398 15792 3674
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15476 3052 15608 3058
rect 15528 3046 15608 3052
rect 15660 3052 15712 3058
rect 15476 2994 15528 3000
rect 15660 2994 15712 3000
rect 15382 2952 15438 2961
rect 15382 2887 15384 2896
rect 15436 2887 15438 2896
rect 15384 2858 15436 2864
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15856 2446 15884 16390
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15948 5370 15976 15846
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16040 2514 16068 15914
rect 16132 7546 16160 17070
rect 16868 15162 16896 19200
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16132 4282 16160 5510
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16210 3360 16266 3369
rect 16316 3346 16344 14894
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16408 4622 16436 9046
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16266 3318 16344 3346
rect 16210 3295 16266 3304
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15028 800 15056 2314
rect 15212 1494 15240 2382
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15200 1488 15252 1494
rect 15200 1430 15252 1436
rect 15304 800 15332 2314
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
<< via2 >>
rect 1582 17992 1638 18048
rect 2778 18944 2834 19000
rect 1766 16224 1822 16280
rect 1674 15952 1730 16008
rect 2134 16088 2190 16144
rect 1398 14184 1454 14240
rect 1674 13232 1730 13288
rect 1582 11328 1638 11384
rect 1398 9424 1454 9480
rect 1582 7520 1638 7576
rect 2410 15444 2412 15464
rect 2412 15444 2464 15464
rect 2464 15444 2466 15464
rect 2410 15408 2466 15444
rect 2410 15136 2466 15192
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 2042 8880 2098 8936
rect 1950 8472 2006 8528
rect 2226 8472 2282 8528
rect 1766 7384 1822 7440
rect 2226 6568 2282 6624
rect 1582 4664 1638 4720
rect 1858 3712 1914 3768
rect 1858 2760 1914 2816
rect 1766 1808 1822 1864
rect 2318 3984 2374 4040
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 2962 11092 2964 11112
rect 2964 11092 3016 11112
rect 3016 11092 3018 11112
rect 2962 11056 3018 11092
rect 2686 10376 2742 10432
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2686 9016 2742 9072
rect 3606 14220 3608 14240
rect 3608 14220 3660 14240
rect 3660 14220 3662 14240
rect 3606 14184 3662 14220
rect 4158 17040 4214 17096
rect 4158 15564 4214 15600
rect 4158 15544 4160 15564
rect 4160 15544 4212 15564
rect 4212 15544 4214 15564
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 4066 13232 4122 13288
rect 3238 12280 3294 12336
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 3698 8608 3754 8664
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2686 5616 2742 5672
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 3330 4684 3386 4720
rect 3330 4664 3332 4684
rect 3332 4664 3384 4684
rect 3384 4664 3386 4684
rect 3238 4276 3294 4312
rect 3238 4256 3240 4276
rect 3240 4256 3292 4276
rect 3292 4256 3294 4276
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 3238 2796 3240 2816
rect 3240 2796 3292 2816
rect 3292 2796 3294 2816
rect 3238 2760 3294 2796
rect 3698 3576 3754 3632
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4986 15852 4988 15872
rect 4988 15852 5040 15872
rect 5040 15852 5042 15872
rect 4986 15816 5042 15852
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 5262 16088 5318 16144
rect 4342 12280 4398 12336
rect 3974 4528 4030 4584
rect 4158 3884 4160 3904
rect 4160 3884 4212 3904
rect 4212 3884 4214 3904
rect 4158 3848 4214 3884
rect 4158 3712 4214 3768
rect 4434 11872 4490 11928
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 5170 13096 5226 13152
rect 4710 12416 4766 12472
rect 5262 12552 5318 12608
rect 4710 12144 4766 12200
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4802 11736 4858 11792
rect 4710 11192 4766 11248
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 5170 12008 5226 12064
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4526 4936 4582 4992
rect 4158 3032 4214 3088
rect 3974 2760 4030 2816
rect 3790 856 3846 912
rect 4526 3984 4582 4040
rect 5078 5480 5134 5536
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 5078 4820 5134 4856
rect 5078 4800 5080 4820
rect 5080 4800 5132 4820
rect 5132 4800 5134 4820
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4710 3984 4766 4040
rect 4526 3440 4582 3496
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 4618 2760 4674 2816
rect 5078 2760 5134 2816
rect 5078 2488 5134 2544
rect 5354 5344 5410 5400
rect 5354 4936 5410 4992
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 6734 16668 6736 16688
rect 6736 16668 6788 16688
rect 6788 16668 6790 16688
rect 6734 16632 6790 16668
rect 7286 16632 7342 16688
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6918 15408 6974 15464
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6550 12688 6606 12744
rect 6366 12144 6422 12200
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6090 7792 6146 7848
rect 4618 2352 4674 2408
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6642 10648 6698 10704
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6642 9424 6698 9480
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 7286 13368 7342 13424
rect 7286 13268 7288 13288
rect 7288 13268 7340 13288
rect 7340 13268 7342 13288
rect 7286 13232 7342 13268
rect 7102 9968 7158 10024
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6458 7384 6514 7440
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6274 5072 6330 5128
rect 6734 5244 6736 5264
rect 6736 5244 6788 5264
rect 6788 5244 6790 5264
rect 6734 5208 6790 5244
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 7562 13232 7618 13288
rect 8206 15544 8262 15600
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8758 12416 8814 12472
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8298 11192 8354 11248
rect 6458 4664 6514 4720
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 7562 5480 7618 5536
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7010 2896 7066 2952
rect 7930 5616 7986 5672
rect 7654 4528 7710 4584
rect 7562 4120 7618 4176
rect 7562 3596 7618 3632
rect 7562 3576 7564 3596
rect 7564 3576 7616 3596
rect 7616 3576 7618 3596
rect 7930 5364 7986 5400
rect 7930 5344 7932 5364
rect 7932 5344 7984 5364
rect 7984 5344 7986 5364
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8298 10240 8354 10296
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8850 5344 8906 5400
rect 8850 5072 8906 5128
rect 8114 4120 8170 4176
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8022 3984 8078 4040
rect 9218 16224 9274 16280
rect 9126 16088 9182 16144
rect 9126 12416 9182 12472
rect 9402 16224 9458 16280
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 9402 14456 9458 14512
rect 9494 12588 9496 12608
rect 9496 12588 9548 12608
rect 9548 12588 9550 12608
rect 9494 12552 9550 12588
rect 9402 11600 9458 11656
rect 9586 9832 9642 9888
rect 9678 9560 9734 9616
rect 9126 5752 9182 5808
rect 9310 6568 9366 6624
rect 9402 6024 9458 6080
rect 9402 5752 9458 5808
rect 9586 5888 9642 5944
rect 9310 5616 9366 5672
rect 9586 5752 9642 5808
rect 10046 11872 10102 11928
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10598 14320 10654 14376
rect 10690 14220 10692 14240
rect 10692 14220 10744 14240
rect 10744 14220 10746 14240
rect 10690 14184 10746 14220
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10322 11872 10378 11928
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 11334 15544 11390 15600
rect 11058 13812 11060 13832
rect 11060 13812 11112 13832
rect 11112 13812 11114 13832
rect 11058 13776 11114 13812
rect 11058 13404 11060 13424
rect 11060 13404 11112 13424
rect 11112 13404 11114 13424
rect 11058 13368 11114 13404
rect 10966 12416 11022 12472
rect 10966 9968 11022 10024
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 9862 4820 9918 4856
rect 9862 4800 9864 4820
rect 9864 4800 9916 4820
rect 9916 4800 9918 4820
rect 9586 4564 9588 4584
rect 9588 4564 9640 4584
rect 9640 4564 9642 4584
rect 9586 4528 9642 4564
rect 9310 4256 9366 4312
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8942 2488 8998 2544
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 8666 1944 8722 2000
rect 9310 3732 9366 3768
rect 9310 3712 9312 3732
rect 9312 3712 9364 3732
rect 9364 3712 9366 3732
rect 9678 3304 9734 3360
rect 9494 1808 9550 1864
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 11058 9560 11114 9616
rect 10506 5480 10562 5536
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 11518 16224 11574 16280
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12438 15700 12494 15736
rect 12438 15680 12440 15700
rect 12440 15680 12492 15700
rect 12492 15680 12494 15700
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12438 14592 12494 14648
rect 11426 12416 11482 12472
rect 12438 14320 12494 14376
rect 11518 10920 11574 10976
rect 11150 6568 11206 6624
rect 10138 3576 10194 3632
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12806 15680 12862 15736
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12254 12164 12310 12200
rect 12254 12144 12256 12164
rect 12256 12144 12308 12164
rect 12308 12144 12310 12164
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 11610 6976 11666 7032
rect 11426 6296 11482 6352
rect 11242 4800 11298 4856
rect 11334 3884 11336 3904
rect 11336 3884 11388 3904
rect 11388 3884 11390 3904
rect 11334 3848 11390 3884
rect 10874 3440 10930 3496
rect 10874 3188 10930 3224
rect 10874 3168 10876 3188
rect 10876 3168 10928 3188
rect 10928 3168 10930 3188
rect 11242 3304 11298 3360
rect 11334 3032 11390 3088
rect 11610 4664 11666 4720
rect 11518 2760 11574 2816
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 13266 14220 13268 14240
rect 13268 14220 13320 14240
rect 13320 14220 13322 14240
rect 13266 14184 13322 14220
rect 11978 9152 12034 9208
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12438 8472 12494 8528
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12346 6296 12402 6352
rect 12070 5636 12126 5672
rect 12070 5616 12072 5636
rect 12072 5616 12124 5636
rect 12124 5616 12126 5636
rect 11886 5364 11942 5400
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 11886 5344 11888 5364
rect 11888 5344 11940 5364
rect 11940 5344 11942 5364
rect 12438 5208 12494 5264
rect 12162 5072 12218 5128
rect 12990 9560 13046 9616
rect 12990 8880 13046 8936
rect 12806 5888 12862 5944
rect 12714 5616 12770 5672
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12162 3032 12218 3088
rect 12162 2760 12218 2816
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12806 4800 12862 4856
rect 12714 3732 12770 3768
rect 12714 3712 12716 3732
rect 12716 3712 12768 3732
rect 12768 3712 12770 3732
rect 12806 3032 12862 3088
rect 13634 16224 13690 16280
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14278 16108 14334 16144
rect 14278 16088 14280 16108
rect 14280 16088 14332 16108
rect 14332 16088 14334 16108
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 13910 15544 13966 15600
rect 13726 14592 13782 14648
rect 13542 14048 13598 14104
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14094 13388 14150 13424
rect 14094 13368 14096 13388
rect 14096 13368 14148 13388
rect 14148 13368 14150 13388
rect 13634 11756 13690 11792
rect 13634 11736 13636 11756
rect 13636 11736 13688 11756
rect 13688 11736 13690 11756
rect 13910 12688 13966 12744
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 13726 11056 13782 11112
rect 14002 11756 14058 11792
rect 14002 11736 14004 11756
rect 14004 11736 14056 11756
rect 14056 11736 14058 11756
rect 14646 13096 14702 13152
rect 15106 16532 15108 16552
rect 15108 16532 15160 16552
rect 15160 16532 15162 16552
rect 15106 16496 15162 16532
rect 15014 12688 15070 12744
rect 14830 12280 14886 12336
rect 14370 11600 14426 11656
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14186 11192 14242 11248
rect 14370 11228 14372 11248
rect 14372 11228 14424 11248
rect 14424 11228 14426 11248
rect 14370 11192 14426 11228
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 14002 10104 14058 10160
rect 14002 9560 14058 9616
rect 14370 9424 14426 9480
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 13910 8744 13966 8800
rect 14002 8628 14058 8664
rect 14002 8608 14004 8628
rect 14004 8608 14056 8628
rect 14056 8608 14058 8628
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 13358 5636 13414 5672
rect 13358 5616 13360 5636
rect 13360 5616 13412 5636
rect 13412 5616 13414 5636
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 13910 5752 13966 5808
rect 14738 9832 14794 9888
rect 14738 8880 14794 8936
rect 15106 9968 15162 10024
rect 15290 8900 15346 8936
rect 15290 8880 15292 8900
rect 15292 8880 15344 8900
rect 15344 8880 15346 8900
rect 14830 6704 14886 6760
rect 13726 3848 13782 3904
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14370 4664 14426 4720
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14186 3052 14242 3088
rect 14186 3032 14188 3052
rect 14188 3032 14240 3052
rect 14240 3032 14242 3052
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 14186 2352 14242 2408
rect 14922 4664 14978 4720
rect 15290 6452 15346 6488
rect 15290 6432 15292 6452
rect 15292 6432 15344 6452
rect 15344 6432 15346 6452
rect 15198 4528 15254 4584
rect 15382 2916 15438 2952
rect 15382 2896 15384 2916
rect 15384 2896 15436 2916
rect 15436 2896 15438 2916
rect 16210 3304 16266 3360
<< metal3 >>
rect 0 19002 800 19032
rect 2773 19002 2839 19005
rect 0 19000 2839 19002
rect 0 18944 2778 19000
rect 2834 18944 2839 19000
rect 0 18942 2839 18944
rect 0 18912 800 18942
rect 2773 18939 2839 18942
rect 0 18050 800 18080
rect 1577 18050 1643 18053
rect 0 18048 1643 18050
rect 0 17992 1582 18048
rect 1638 17992 1643 18048
rect 0 17990 1643 17992
rect 0 17960 800 17990
rect 1577 17987 1643 17990
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 0 17008 800 17128
rect 3550 17036 3556 17100
rect 3620 17098 3626 17100
rect 4153 17098 4219 17101
rect 3620 17096 4219 17098
rect 3620 17040 4158 17096
rect 4214 17040 4219 17096
rect 3620 17038 4219 17040
rect 3620 17036 3626 17038
rect 4153 17035 4219 17038
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 6729 16690 6795 16693
rect 7281 16690 7347 16693
rect 6729 16688 7347 16690
rect 6729 16632 6734 16688
rect 6790 16632 7286 16688
rect 7342 16632 7347 16688
rect 6729 16630 7347 16632
rect 6729 16627 6795 16630
rect 7281 16627 7347 16630
rect 16400 16600 17200 16720
rect 15101 16554 15167 16557
rect 2730 16552 15167 16554
rect 2730 16496 15106 16552
rect 15162 16496 15167 16552
rect 2730 16494 15167 16496
rect 1761 16282 1827 16285
rect 1761 16280 2330 16282
rect 1761 16224 1766 16280
rect 1822 16224 2330 16280
rect 1761 16222 2330 16224
rect 1761 16219 1827 16222
rect 0 16146 800 16176
rect 2129 16146 2195 16149
rect 0 16144 2195 16146
rect 0 16088 2134 16144
rect 2190 16088 2195 16144
rect 0 16086 2195 16088
rect 2270 16146 2330 16222
rect 2730 16146 2790 16494
rect 15101 16491 15167 16494
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 9213 16282 9279 16285
rect 9397 16282 9463 16285
rect 11513 16282 11579 16285
rect 9213 16280 11579 16282
rect 9213 16224 9218 16280
rect 9274 16224 9402 16280
rect 9458 16224 11518 16280
rect 11574 16224 11579 16280
rect 9213 16222 11579 16224
rect 9213 16219 9279 16222
rect 9397 16219 9463 16222
rect 11513 16219 11579 16222
rect 13629 16284 13695 16285
rect 13629 16280 13676 16284
rect 13740 16282 13746 16284
rect 13629 16224 13634 16280
rect 13629 16220 13676 16224
rect 13740 16222 13786 16282
rect 13740 16220 13746 16222
rect 13629 16219 13695 16220
rect 2270 16086 2790 16146
rect 5257 16146 5323 16149
rect 9121 16146 9187 16149
rect 14273 16146 14339 16149
rect 5257 16144 9187 16146
rect 5257 16088 5262 16144
rect 5318 16088 9126 16144
rect 9182 16088 9187 16144
rect 5257 16086 9187 16088
rect 0 16056 800 16086
rect 2129 16083 2195 16086
rect 5257 16083 5323 16086
rect 9121 16083 9187 16086
rect 12390 16144 14339 16146
rect 12390 16088 14278 16144
rect 14334 16088 14339 16144
rect 12390 16086 14339 16088
rect 1669 16010 1735 16013
rect 12390 16010 12450 16086
rect 14273 16083 14339 16086
rect 1669 16008 12450 16010
rect 1669 15952 1674 16008
rect 1730 15952 12450 16008
rect 1669 15950 12450 15952
rect 1669 15947 1735 15950
rect 4981 15874 5047 15877
rect 5206 15874 5212 15876
rect 4981 15872 5212 15874
rect 4981 15816 4986 15872
rect 5042 15816 5212 15872
rect 4981 15814 5212 15816
rect 4981 15811 5047 15814
rect 5206 15812 5212 15814
rect 5276 15812 5282 15876
rect 2820 15808 3136 15809
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 12433 15738 12499 15741
rect 12566 15738 12572 15740
rect 12433 15736 12572 15738
rect 12433 15680 12438 15736
rect 12494 15680 12572 15736
rect 12433 15678 12572 15680
rect 12433 15675 12499 15678
rect 12566 15676 12572 15678
rect 12636 15676 12642 15740
rect 12801 15738 12867 15741
rect 12934 15738 12940 15740
rect 12801 15736 12940 15738
rect 12801 15680 12806 15736
rect 12862 15680 12940 15736
rect 12801 15678 12940 15680
rect 12801 15675 12867 15678
rect 12934 15676 12940 15678
rect 13004 15676 13010 15740
rect 4153 15602 4219 15605
rect 8201 15602 8267 15605
rect 4153 15600 8267 15602
rect 4153 15544 4158 15600
rect 4214 15544 8206 15600
rect 8262 15544 8267 15600
rect 4153 15542 8267 15544
rect 4153 15539 4219 15542
rect 8201 15539 8267 15542
rect 9070 15540 9076 15604
rect 9140 15602 9146 15604
rect 11329 15602 11395 15605
rect 9140 15600 11395 15602
rect 9140 15544 11334 15600
rect 11390 15544 11395 15600
rect 9140 15542 11395 15544
rect 9140 15540 9146 15542
rect 11329 15539 11395 15542
rect 13905 15602 13971 15605
rect 14774 15602 14780 15604
rect 13905 15600 14780 15602
rect 13905 15544 13910 15600
rect 13966 15544 14780 15600
rect 13905 15542 14780 15544
rect 13905 15539 13971 15542
rect 14774 15540 14780 15542
rect 14844 15540 14850 15604
rect 2405 15466 2471 15469
rect 6913 15466 6979 15469
rect 2405 15464 6979 15466
rect 2405 15408 2410 15464
rect 2466 15408 6918 15464
rect 6974 15408 6979 15464
rect 2405 15406 6979 15408
rect 2405 15403 2471 15406
rect 6913 15403 6979 15406
rect 4694 15264 5010 15265
rect 0 15194 800 15224
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 2405 15194 2471 15197
rect 0 15192 2471 15194
rect 0 15136 2410 15192
rect 2466 15136 2471 15192
rect 0 15134 2471 15136
rect 0 15104 800 15134
rect 2405 15131 2471 15134
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 12433 14650 12499 14653
rect 13721 14650 13787 14653
rect 12433 14648 13787 14650
rect 12433 14592 12438 14648
rect 12494 14592 13726 14648
rect 13782 14592 13787 14648
rect 12433 14590 13787 14592
rect 12433 14587 12499 14590
rect 13721 14587 13787 14590
rect 9397 14514 9463 14517
rect 13854 14514 13860 14516
rect 9397 14512 13860 14514
rect 9397 14456 9402 14512
rect 9458 14456 13860 14512
rect 9397 14454 13860 14456
rect 9397 14451 9463 14454
rect 13854 14452 13860 14454
rect 13924 14452 13930 14516
rect 10593 14378 10659 14381
rect 12433 14378 12499 14381
rect 10593 14376 12499 14378
rect 10593 14320 10598 14376
rect 10654 14320 12438 14376
rect 12494 14320 12499 14376
rect 10593 14318 12499 14320
rect 10593 14315 10659 14318
rect 12433 14315 12499 14318
rect 0 14242 800 14272
rect 1393 14242 1459 14245
rect 0 14240 1459 14242
rect 0 14184 1398 14240
rect 1454 14184 1459 14240
rect 0 14182 1459 14184
rect 0 14152 800 14182
rect 1393 14179 1459 14182
rect 3366 14180 3372 14244
rect 3436 14242 3442 14244
rect 3601 14242 3667 14245
rect 3436 14240 3667 14242
rect 3436 14184 3606 14240
rect 3662 14184 3667 14240
rect 3436 14182 3667 14184
rect 3436 14180 3442 14182
rect 3601 14179 3667 14182
rect 9438 14180 9444 14244
rect 9508 14242 9514 14244
rect 10685 14242 10751 14245
rect 9508 14240 10751 14242
rect 9508 14184 10690 14240
rect 10746 14184 10751 14240
rect 9508 14182 10751 14184
rect 9508 14180 9514 14182
rect 10685 14179 10751 14182
rect 13261 14242 13327 14245
rect 13261 14240 13554 14242
rect 13261 14184 13266 14240
rect 13322 14184 13554 14240
rect 13261 14182 13554 14184
rect 13261 14179 13327 14182
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 13494 14109 13554 14182
rect 13494 14104 13603 14109
rect 13494 14048 13542 14104
rect 13598 14048 13603 14104
rect 13494 14046 13603 14048
rect 13537 14043 13603 14046
rect 9622 13772 9628 13836
rect 9692 13834 9698 13836
rect 11053 13834 11119 13837
rect 9692 13832 11119 13834
rect 9692 13776 11058 13832
rect 11114 13776 11119 13832
rect 9692 13774 11119 13776
rect 9692 13772 9698 13774
rect 11053 13771 11119 13774
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 7281 13426 7347 13429
rect 11053 13426 11119 13429
rect 11646 13426 11652 13428
rect 7281 13424 11652 13426
rect 7281 13368 7286 13424
rect 7342 13368 11058 13424
rect 11114 13368 11652 13424
rect 7281 13366 11652 13368
rect 7281 13363 7347 13366
rect 11053 13363 11119 13366
rect 11646 13364 11652 13366
rect 11716 13364 11722 13428
rect 13854 13364 13860 13428
rect 13924 13426 13930 13428
rect 14089 13426 14155 13429
rect 13924 13424 14155 13426
rect 13924 13368 14094 13424
rect 14150 13368 14155 13424
rect 13924 13366 14155 13368
rect 13924 13364 13930 13366
rect 14089 13363 14155 13366
rect 0 13290 800 13320
rect 1669 13290 1735 13293
rect 0 13288 1735 13290
rect 0 13232 1674 13288
rect 1730 13232 1735 13288
rect 0 13230 1735 13232
rect 0 13200 800 13230
rect 1669 13227 1735 13230
rect 4061 13290 4127 13293
rect 7281 13290 7347 13293
rect 7557 13290 7623 13293
rect 4061 13288 7623 13290
rect 4061 13232 4066 13288
rect 4122 13232 7286 13288
rect 7342 13232 7562 13288
rect 7618 13232 7623 13288
rect 4061 13230 7623 13232
rect 4061 13227 4127 13230
rect 7281 13227 7347 13230
rect 7557 13227 7623 13230
rect 5165 13154 5231 13157
rect 14641 13154 14707 13157
rect 5165 13152 5274 13154
rect 5165 13096 5170 13152
rect 5226 13096 5274 13152
rect 5165 13091 5274 13096
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 5214 12613 5274 13091
rect 14598 13152 14707 13154
rect 14598 13096 14646 13152
rect 14702 13096 14707 13152
rect 14598 13091 14707 13096
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 6545 12746 6611 12749
rect 9806 12746 9812 12748
rect 6545 12744 9812 12746
rect 6545 12688 6550 12744
rect 6606 12688 9812 12744
rect 6545 12686 9812 12688
rect 6545 12683 6611 12686
rect 9806 12684 9812 12686
rect 9876 12746 9882 12748
rect 13905 12746 13971 12749
rect 14598 12746 14658 13091
rect 15009 12748 15075 12749
rect 9876 12744 14658 12746
rect 9876 12688 13910 12744
rect 13966 12688 14658 12744
rect 9876 12686 14658 12688
rect 9876 12684 9882 12686
rect 13905 12683 13971 12686
rect 14958 12684 14964 12748
rect 15028 12746 15075 12748
rect 15028 12744 15120 12746
rect 15070 12688 15120 12744
rect 15028 12686 15120 12688
rect 15028 12684 15075 12686
rect 15009 12683 15075 12684
rect 5214 12608 5323 12613
rect 5214 12552 5262 12608
rect 5318 12552 5323 12608
rect 5214 12550 5323 12552
rect 5257 12547 5323 12550
rect 8150 12548 8156 12612
rect 8220 12610 8226 12612
rect 9489 12610 9555 12613
rect 8220 12608 9555 12610
rect 8220 12552 9494 12608
rect 9550 12552 9555 12608
rect 8220 12550 9555 12552
rect 8220 12548 8226 12550
rect 9489 12547 9555 12550
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 4705 12474 4771 12477
rect 4478 12472 4771 12474
rect 4478 12416 4710 12472
rect 4766 12416 4771 12472
rect 4478 12414 4771 12416
rect 0 12338 800 12368
rect 3233 12338 3299 12341
rect 0 12336 3299 12338
rect 0 12280 3238 12336
rect 3294 12280 3299 12336
rect 0 12278 3299 12280
rect 0 12248 800 12278
rect 3233 12275 3299 12278
rect 4337 12338 4403 12341
rect 4478 12338 4538 12414
rect 4705 12411 4771 12414
rect 8753 12474 8819 12477
rect 9121 12474 9187 12477
rect 8753 12472 9187 12474
rect 8753 12416 8758 12472
rect 8814 12416 9126 12472
rect 9182 12416 9187 12472
rect 8753 12414 9187 12416
rect 8753 12411 8819 12414
rect 9121 12411 9187 12414
rect 10961 12474 11027 12477
rect 11421 12474 11487 12477
rect 10961 12472 11487 12474
rect 10961 12416 10966 12472
rect 11022 12416 11426 12472
rect 11482 12416 11487 12472
rect 10961 12414 11487 12416
rect 10961 12411 11027 12414
rect 11421 12411 11487 12414
rect 14825 12340 14891 12341
rect 4337 12336 4538 12338
rect 4337 12280 4342 12336
rect 4398 12280 4538 12336
rect 4337 12278 4538 12280
rect 4337 12275 4403 12278
rect 14774 12276 14780 12340
rect 14844 12338 14891 12340
rect 14844 12336 14936 12338
rect 14886 12280 14936 12336
rect 14844 12278 14936 12280
rect 14844 12276 14891 12278
rect 14825 12275 14891 12276
rect 4705 12202 4771 12205
rect 6361 12202 6427 12205
rect 12014 12202 12020 12204
rect 4705 12200 5274 12202
rect 4705 12144 4710 12200
rect 4766 12144 5274 12200
rect 4705 12142 5274 12144
rect 4705 12139 4771 12142
rect 5214 12069 5274 12142
rect 6361 12200 12020 12202
rect 6361 12144 6366 12200
rect 6422 12144 12020 12200
rect 6361 12142 12020 12144
rect 6361 12139 6427 12142
rect 12014 12140 12020 12142
rect 12084 12202 12090 12204
rect 12249 12202 12315 12205
rect 12084 12200 12315 12202
rect 12084 12144 12254 12200
rect 12310 12144 12315 12200
rect 12084 12142 12315 12144
rect 12084 12140 12090 12142
rect 12249 12139 12315 12142
rect 5165 12064 5274 12069
rect 5165 12008 5170 12064
rect 5226 12008 5274 12064
rect 5165 12006 5274 12008
rect 5165 12003 5231 12006
rect 4694 12000 5010 12001
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 4429 11930 4495 11933
rect 10041 11930 10107 11933
rect 10317 11930 10383 11933
rect 4429 11928 4538 11930
rect 4429 11872 4434 11928
rect 4490 11872 4538 11928
rect 4429 11867 4538 11872
rect 10041 11928 10383 11930
rect 10041 11872 10046 11928
rect 10102 11872 10322 11928
rect 10378 11872 10383 11928
rect 10041 11870 10383 11872
rect 10041 11867 10107 11870
rect 10317 11867 10383 11870
rect 4478 11794 4538 11867
rect 4797 11794 4863 11797
rect 13629 11796 13695 11797
rect 13629 11794 13676 11796
rect 4478 11792 4863 11794
rect 4478 11736 4802 11792
rect 4858 11736 4863 11792
rect 4478 11734 4863 11736
rect 13584 11792 13676 11794
rect 13740 11794 13746 11796
rect 13997 11794 14063 11797
rect 13740 11792 14063 11794
rect 13584 11736 13634 11792
rect 13740 11736 14002 11792
rect 14058 11736 14063 11792
rect 13584 11734 13676 11736
rect 4797 11731 4863 11734
rect 13629 11732 13676 11734
rect 13740 11734 14063 11736
rect 13740 11732 13746 11734
rect 13629 11731 13695 11732
rect 13997 11731 14063 11734
rect 9397 11658 9463 11661
rect 14365 11658 14431 11661
rect 9397 11656 14431 11658
rect 9397 11600 9402 11656
rect 9458 11600 14370 11656
rect 14426 11600 14431 11656
rect 9397 11598 14431 11600
rect 9397 11595 9463 11598
rect 14365 11595 14431 11598
rect 2820 11456 3136 11457
rect 0 11386 800 11416
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 1577 11386 1643 11389
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 4705 11250 4771 11253
rect 8293 11250 8359 11253
rect 4705 11248 8359 11250
rect 4705 11192 4710 11248
rect 4766 11192 8298 11248
rect 8354 11192 8359 11248
rect 4705 11190 8359 11192
rect 4705 11187 4771 11190
rect 8293 11187 8359 11190
rect 8886 11188 8892 11252
rect 8956 11250 8962 11252
rect 9622 11250 9628 11252
rect 8956 11190 9628 11250
rect 8956 11188 8962 11190
rect 9622 11188 9628 11190
rect 9692 11188 9698 11252
rect 13670 11188 13676 11252
rect 13740 11250 13746 11252
rect 14181 11250 14247 11253
rect 14365 11250 14431 11253
rect 13740 11248 14431 11250
rect 13740 11192 14186 11248
rect 14242 11192 14370 11248
rect 14426 11192 14431 11248
rect 13740 11190 14431 11192
rect 13740 11188 13746 11190
rect 14181 11187 14247 11190
rect 14365 11187 14431 11190
rect 2957 11114 3023 11117
rect 2957 11112 9690 11114
rect 2957 11056 2962 11112
rect 3018 11056 9690 11112
rect 2957 11054 9690 11056
rect 2957 11051 3023 11054
rect 9630 10978 9690 11054
rect 12566 11052 12572 11116
rect 12636 11114 12642 11116
rect 13721 11114 13787 11117
rect 12636 11112 13787 11114
rect 12636 11056 13726 11112
rect 13782 11056 13787 11112
rect 12636 11054 13787 11056
rect 12636 11052 12642 11054
rect 13721 11051 13787 11054
rect 11513 10978 11579 10981
rect 9630 10976 11579 10978
rect 9630 10920 11518 10976
rect 11574 10920 11579 10976
rect 9630 10918 11579 10920
rect 11513 10915 11579 10918
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 3550 10644 3556 10708
rect 3620 10706 3626 10708
rect 6637 10706 6703 10709
rect 3620 10704 6703 10706
rect 3620 10648 6642 10704
rect 6698 10648 6703 10704
rect 3620 10646 6703 10648
rect 3620 10644 3626 10646
rect 6637 10643 6703 10646
rect 0 10434 800 10464
rect 2681 10434 2747 10437
rect 0 10432 2747 10434
rect 0 10376 2686 10432
rect 2742 10376 2747 10432
rect 0 10374 2747 10376
rect 0 10344 800 10374
rect 2681 10371 2747 10374
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 8293 10298 8359 10301
rect 9070 10298 9076 10300
rect 8293 10296 9076 10298
rect 8293 10240 8298 10296
rect 8354 10240 9076 10296
rect 8293 10238 9076 10240
rect 8293 10235 8359 10238
rect 9070 10236 9076 10238
rect 9140 10236 9146 10300
rect 13670 10100 13676 10164
rect 13740 10162 13746 10164
rect 13997 10162 14063 10165
rect 13740 10160 14063 10162
rect 13740 10104 14002 10160
rect 14058 10104 14063 10160
rect 13740 10102 14063 10104
rect 13740 10100 13746 10102
rect 13997 10099 14063 10102
rect 7097 10026 7163 10029
rect 10961 10026 11027 10029
rect 7097 10024 11027 10026
rect 7097 9968 7102 10024
rect 7158 9968 10966 10024
rect 11022 9968 11027 10024
rect 7097 9966 11027 9968
rect 7097 9963 7163 9966
rect 10961 9963 11027 9966
rect 15101 10026 15167 10029
rect 16400 10026 17200 10056
rect 15101 10024 17200 10026
rect 15101 9968 15106 10024
rect 15162 9968 17200 10024
rect 15101 9966 17200 9968
rect 15101 9963 15167 9966
rect 16400 9936 17200 9966
rect 9581 9890 9647 9893
rect 14733 9890 14799 9893
rect 14958 9890 14964 9892
rect 9581 9888 9690 9890
rect 9581 9832 9586 9888
rect 9642 9832 9690 9888
rect 9581 9827 9690 9832
rect 14733 9888 14964 9890
rect 14733 9832 14738 9888
rect 14794 9832 14964 9888
rect 14733 9830 14964 9832
rect 14733 9827 14799 9830
rect 14958 9828 14964 9830
rect 15028 9828 15034 9892
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 9630 9621 9690 9827
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 9630 9616 9739 9621
rect 9630 9560 9678 9616
rect 9734 9560 9739 9616
rect 9630 9558 9739 9560
rect 9673 9555 9739 9558
rect 11053 9618 11119 9621
rect 11278 9618 11284 9620
rect 11053 9616 11284 9618
rect 11053 9560 11058 9616
rect 11114 9560 11284 9616
rect 11053 9558 11284 9560
rect 11053 9555 11119 9558
rect 11278 9556 11284 9558
rect 11348 9618 11354 9620
rect 12985 9618 13051 9621
rect 11348 9616 13051 9618
rect 11348 9560 12990 9616
rect 13046 9560 13051 9616
rect 11348 9558 13051 9560
rect 11348 9556 11354 9558
rect 12985 9555 13051 9558
rect 13997 9618 14063 9621
rect 14774 9618 14780 9620
rect 13997 9616 14780 9618
rect 13997 9560 14002 9616
rect 14058 9560 14780 9616
rect 13997 9558 14780 9560
rect 13997 9555 14063 9558
rect 14774 9556 14780 9558
rect 14844 9556 14850 9620
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 6637 9482 6703 9485
rect 12566 9482 12572 9484
rect 6637 9480 12572 9482
rect 6637 9424 6642 9480
rect 6698 9424 12572 9480
rect 6637 9422 12572 9424
rect 6637 9419 6703 9422
rect 12566 9420 12572 9422
rect 12636 9420 12642 9484
rect 14365 9482 14431 9485
rect 14590 9482 14596 9484
rect 14365 9480 14596 9482
rect 14365 9424 14370 9480
rect 14426 9424 14596 9480
rect 14365 9422 14596 9424
rect 14365 9419 14431 9422
rect 14590 9420 14596 9422
rect 14660 9420 14666 9484
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 11830 9148 11836 9212
rect 11900 9210 11906 9212
rect 11973 9210 12039 9213
rect 11900 9208 12039 9210
rect 11900 9152 11978 9208
rect 12034 9152 12039 9208
rect 11900 9150 12039 9152
rect 11900 9148 11906 9150
rect 11973 9147 12039 9150
rect 2681 9074 2747 9077
rect 8150 9074 8156 9076
rect 2681 9072 8156 9074
rect 2681 9016 2686 9072
rect 2742 9016 8156 9072
rect 2681 9014 8156 9016
rect 2681 9011 2747 9014
rect 8150 9012 8156 9014
rect 8220 9074 8226 9076
rect 9622 9074 9628 9076
rect 8220 9014 9628 9074
rect 8220 9012 8226 9014
rect 9622 9012 9628 9014
rect 9692 9012 9698 9076
rect 2037 8938 2103 8941
rect 12985 8938 13051 8941
rect 14733 8938 14799 8941
rect 15285 8938 15351 8941
rect 2037 8936 15351 8938
rect 2037 8880 2042 8936
rect 2098 8880 12990 8936
rect 13046 8880 14738 8936
rect 14794 8880 15290 8936
rect 15346 8880 15351 8936
rect 2037 8878 15351 8880
rect 2037 8875 2103 8878
rect 12985 8875 13051 8878
rect 14733 8875 14799 8878
rect 15285 8875 15351 8878
rect 13905 8802 13971 8805
rect 13678 8800 13971 8802
rect 13678 8744 13910 8800
rect 13966 8744 13971 8800
rect 13678 8742 13971 8744
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 3550 8604 3556 8668
rect 3620 8666 3626 8668
rect 3693 8666 3759 8669
rect 3620 8664 3759 8666
rect 3620 8608 3698 8664
rect 3754 8608 3759 8664
rect 3620 8606 3759 8608
rect 3620 8604 3626 8606
rect 3693 8603 3759 8606
rect 0 8530 800 8560
rect 1945 8530 2011 8533
rect 0 8528 2011 8530
rect 0 8472 1950 8528
rect 2006 8472 2011 8528
rect 0 8470 2011 8472
rect 0 8440 800 8470
rect 1945 8467 2011 8470
rect 2221 8530 2287 8533
rect 3550 8530 3556 8532
rect 2221 8528 3556 8530
rect 2221 8472 2226 8528
rect 2282 8472 3556 8528
rect 2221 8470 3556 8472
rect 2221 8467 2287 8470
rect 3550 8468 3556 8470
rect 3620 8530 3626 8532
rect 8886 8530 8892 8532
rect 3620 8470 8892 8530
rect 3620 8468 3626 8470
rect 8886 8468 8892 8470
rect 8956 8468 8962 8532
rect 12433 8530 12499 8533
rect 13678 8530 13738 8742
rect 13905 8739 13971 8742
rect 13854 8604 13860 8668
rect 13924 8666 13930 8668
rect 13997 8666 14063 8669
rect 13924 8664 14063 8666
rect 13924 8608 14002 8664
rect 14058 8608 14063 8664
rect 13924 8606 14063 8608
rect 13924 8604 13930 8606
rect 13997 8603 14063 8606
rect 12433 8528 13738 8530
rect 12433 8472 12438 8528
rect 12494 8472 13738 8528
rect 12433 8470 13738 8472
rect 12433 8467 12499 8470
rect 2820 8192 3136 8193
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 6085 7850 6151 7853
rect 13854 7850 13860 7852
rect 6085 7848 13860 7850
rect 6085 7792 6090 7848
rect 6146 7792 13860 7848
rect 6085 7790 13860 7792
rect 6085 7787 6151 7790
rect 13854 7788 13860 7790
rect 13924 7788 13930 7852
rect 4694 7648 5010 7649
rect 0 7578 800 7608
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 1761 7442 1827 7445
rect 6453 7442 6519 7445
rect 1761 7440 6519 7442
rect 1761 7384 1766 7440
rect 1822 7384 6458 7440
rect 6514 7384 6519 7440
rect 1761 7382 6519 7384
rect 1761 7379 1827 7382
rect 6453 7379 6519 7382
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 11605 7036 11671 7037
rect 11605 7034 11652 7036
rect 11560 7032 11652 7034
rect 11560 6976 11610 7032
rect 11560 6974 11652 6976
rect 11605 6972 11652 6974
rect 11716 6972 11722 7036
rect 11605 6971 11671 6972
rect 14825 6764 14891 6765
rect 14774 6762 14780 6764
rect 14734 6702 14780 6762
rect 14844 6760 14891 6764
rect 14886 6704 14891 6760
rect 14774 6700 14780 6702
rect 14844 6700 14891 6704
rect 14825 6699 14891 6700
rect 0 6626 800 6656
rect 2221 6626 2287 6629
rect 0 6624 2287 6626
rect 0 6568 2226 6624
rect 2282 6568 2287 6624
rect 0 6566 2287 6568
rect 0 6536 800 6566
rect 2221 6563 2287 6566
rect 9305 6626 9371 6629
rect 11145 6626 11211 6629
rect 9305 6624 11211 6626
rect 9305 6568 9310 6624
rect 9366 6568 11150 6624
rect 11206 6568 11211 6624
rect 9305 6566 11211 6568
rect 9305 6563 9371 6566
rect 11145 6563 11211 6566
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 14590 6428 14596 6492
rect 14660 6490 14666 6492
rect 15285 6490 15351 6493
rect 14660 6488 15351 6490
rect 14660 6432 15290 6488
rect 15346 6432 15351 6488
rect 14660 6430 15351 6432
rect 14660 6428 14666 6430
rect 15285 6427 15351 6430
rect 9622 6292 9628 6356
rect 9692 6354 9698 6356
rect 11421 6354 11487 6357
rect 12341 6354 12407 6357
rect 9692 6352 12407 6354
rect 9692 6296 11426 6352
rect 11482 6296 12346 6352
rect 12402 6296 12407 6352
rect 9692 6294 12407 6296
rect 9692 6292 9698 6294
rect 11421 6291 11487 6294
rect 12341 6291 12407 6294
rect 9070 6020 9076 6084
rect 9140 6082 9146 6084
rect 9397 6082 9463 6085
rect 9140 6080 9463 6082
rect 9140 6024 9402 6080
rect 9458 6024 9463 6080
rect 9140 6022 9463 6024
rect 9140 6020 9146 6022
rect 9397 6019 9463 6022
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 14064 5951 14380 5952
rect 9254 5884 9260 5948
rect 9324 5946 9330 5948
rect 9581 5946 9647 5949
rect 12801 5946 12867 5949
rect 9324 5944 9647 5946
rect 9324 5888 9586 5944
rect 9642 5888 9647 5944
rect 9324 5886 9647 5888
rect 9324 5884 9330 5886
rect 9581 5883 9647 5886
rect 10734 5944 12867 5946
rect 10734 5888 12806 5944
rect 12862 5888 12867 5944
rect 10734 5886 12867 5888
rect 9121 5810 9187 5813
rect 9397 5810 9463 5813
rect 9121 5808 9463 5810
rect 9121 5752 9126 5808
rect 9182 5752 9402 5808
rect 9458 5752 9463 5808
rect 9121 5750 9463 5752
rect 9121 5747 9187 5750
rect 9397 5747 9463 5750
rect 9581 5810 9647 5813
rect 10734 5810 10794 5886
rect 12801 5883 12867 5886
rect 9581 5808 10794 5810
rect 9581 5752 9586 5808
rect 9642 5752 10794 5808
rect 9581 5750 10794 5752
rect 9581 5747 9647 5750
rect 12014 5748 12020 5812
rect 12084 5810 12090 5812
rect 13905 5810 13971 5813
rect 12084 5808 13971 5810
rect 12084 5752 13910 5808
rect 13966 5752 13971 5808
rect 12084 5750 13971 5752
rect 12084 5748 12090 5750
rect 13905 5747 13971 5750
rect 0 5674 800 5704
rect 2681 5674 2747 5677
rect 7925 5676 7991 5677
rect 0 5672 2747 5674
rect 0 5616 2686 5672
rect 2742 5616 2747 5672
rect 0 5614 2747 5616
rect 0 5584 800 5614
rect 2681 5611 2747 5614
rect 5206 5612 5212 5676
rect 5276 5674 5282 5676
rect 7925 5674 7972 5676
rect 5276 5672 7972 5674
rect 5276 5616 7930 5672
rect 5276 5614 7972 5616
rect 5276 5612 5282 5614
rect 7925 5612 7972 5614
rect 8036 5612 8042 5676
rect 9305 5674 9371 5677
rect 11830 5674 11836 5676
rect 8158 5614 8954 5674
rect 7925 5611 7991 5612
rect 5073 5538 5139 5541
rect 7557 5538 7623 5541
rect 8158 5538 8218 5614
rect 5073 5536 8218 5538
rect 5073 5480 5078 5536
rect 5134 5480 7562 5536
rect 7618 5480 8218 5536
rect 5073 5478 8218 5480
rect 8894 5538 8954 5614
rect 9305 5672 11836 5674
rect 9305 5616 9310 5672
rect 9366 5616 11836 5672
rect 9305 5614 11836 5616
rect 9305 5611 9371 5614
rect 11830 5612 11836 5614
rect 11900 5674 11906 5676
rect 12065 5674 12131 5677
rect 11900 5672 12131 5674
rect 11900 5616 12070 5672
rect 12126 5616 12131 5672
rect 11900 5614 12131 5616
rect 11900 5612 11906 5614
rect 12065 5611 12131 5614
rect 12709 5674 12775 5677
rect 12934 5674 12940 5676
rect 12709 5672 12940 5674
rect 12709 5616 12714 5672
rect 12770 5616 12940 5672
rect 12709 5614 12940 5616
rect 12709 5611 12775 5614
rect 12934 5612 12940 5614
rect 13004 5674 13010 5676
rect 13353 5674 13419 5677
rect 13004 5672 13419 5674
rect 13004 5616 13358 5672
rect 13414 5616 13419 5672
rect 13004 5614 13419 5616
rect 13004 5612 13010 5614
rect 13353 5611 13419 5614
rect 10501 5538 10567 5541
rect 8894 5536 10567 5538
rect 8894 5480 10506 5536
rect 10562 5480 10567 5536
rect 8894 5478 10567 5480
rect 5073 5475 5139 5478
rect 7557 5475 7623 5478
rect 10501 5475 10567 5478
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 5349 5402 5415 5405
rect 7925 5402 7991 5405
rect 5349 5400 7991 5402
rect 5349 5344 5354 5400
rect 5410 5344 7930 5400
rect 7986 5344 7991 5400
rect 5349 5342 7991 5344
rect 5349 5339 5415 5342
rect 7925 5339 7991 5342
rect 8845 5402 8911 5405
rect 11881 5402 11947 5405
rect 8845 5400 11947 5402
rect 8845 5344 8850 5400
rect 8906 5344 11886 5400
rect 11942 5344 11947 5400
rect 8845 5342 11947 5344
rect 8845 5339 8911 5342
rect 11881 5339 11947 5342
rect 6729 5266 6795 5269
rect 12433 5266 12499 5269
rect 6729 5264 12499 5266
rect 6729 5208 6734 5264
rect 6790 5208 12438 5264
rect 12494 5208 12499 5264
rect 6729 5206 12499 5208
rect 6729 5203 6795 5206
rect 12433 5203 12499 5206
rect 6269 5130 6335 5133
rect 8845 5130 8911 5133
rect 6269 5128 8911 5130
rect 6269 5072 6274 5128
rect 6330 5072 8850 5128
rect 8906 5072 8911 5128
rect 6269 5070 8911 5072
rect 6269 5067 6335 5070
rect 8845 5067 8911 5070
rect 9438 5068 9444 5132
rect 9508 5130 9514 5132
rect 12157 5130 12223 5133
rect 9508 5128 12223 5130
rect 9508 5072 12162 5128
rect 12218 5072 12223 5128
rect 9508 5070 12223 5072
rect 9508 5068 9514 5070
rect 12157 5067 12223 5070
rect 4521 4994 4587 4997
rect 5349 4994 5415 4997
rect 4521 4992 5415 4994
rect 4521 4936 4526 4992
rect 4582 4936 5354 4992
rect 5410 4936 5415 4992
rect 4521 4934 5415 4936
rect 4521 4931 4587 4934
rect 5349 4931 5415 4934
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 5073 4858 5139 4861
rect 9857 4860 9923 4861
rect 5206 4858 5212 4860
rect 5073 4856 5212 4858
rect 5073 4800 5078 4856
rect 5134 4800 5212 4856
rect 5073 4798 5212 4800
rect 5073 4795 5139 4798
rect 5206 4796 5212 4798
rect 5276 4796 5282 4860
rect 9806 4796 9812 4860
rect 9876 4858 9923 4860
rect 11237 4858 11303 4861
rect 12801 4858 12867 4861
rect 9876 4856 9968 4858
rect 9918 4800 9968 4856
rect 9876 4798 9968 4800
rect 11237 4856 12867 4858
rect 11237 4800 11242 4856
rect 11298 4800 12806 4856
rect 12862 4800 12867 4856
rect 11237 4798 12867 4800
rect 9876 4796 9923 4798
rect 9857 4795 9923 4796
rect 11237 4795 11303 4798
rect 12801 4795 12867 4798
rect 0 4722 800 4752
rect 1577 4722 1643 4725
rect 3325 4724 3391 4725
rect 3325 4722 3372 4724
rect 0 4720 1643 4722
rect 0 4664 1582 4720
rect 1638 4664 1643 4720
rect 0 4662 1643 4664
rect 3280 4720 3372 4722
rect 3436 4722 3442 4724
rect 6453 4722 6519 4725
rect 3436 4720 6519 4722
rect 3280 4664 3330 4720
rect 3436 4664 6458 4720
rect 6514 4664 6519 4720
rect 3280 4662 3372 4664
rect 0 4632 800 4662
rect 1577 4659 1643 4662
rect 3325 4660 3372 4662
rect 3436 4662 6519 4664
rect 3436 4660 3442 4662
rect 3325 4659 3391 4660
rect 6453 4659 6519 4662
rect 11605 4722 11671 4725
rect 14365 4722 14431 4725
rect 14917 4722 14983 4725
rect 11605 4720 14983 4722
rect 11605 4664 11610 4720
rect 11666 4664 14370 4720
rect 14426 4664 14922 4720
rect 14978 4664 14983 4720
rect 11605 4662 14983 4664
rect 11605 4659 11671 4662
rect 14365 4659 14431 4662
rect 14917 4659 14983 4662
rect 3969 4586 4035 4589
rect 7649 4586 7715 4589
rect 3969 4584 7715 4586
rect 3969 4528 3974 4584
rect 4030 4528 7654 4584
rect 7710 4528 7715 4584
rect 3969 4526 7715 4528
rect 3969 4523 4035 4526
rect 7649 4523 7715 4526
rect 9581 4586 9647 4589
rect 15193 4586 15259 4589
rect 9581 4584 15259 4586
rect 9581 4528 9586 4584
rect 9642 4528 15198 4584
rect 15254 4528 15259 4584
rect 9581 4526 15259 4528
rect 9581 4523 9647 4526
rect 15193 4523 15259 4526
rect 4694 4384 5010 4385
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 3233 4314 3299 4317
rect 3550 4314 3556 4316
rect 3233 4312 3556 4314
rect 3233 4256 3238 4312
rect 3294 4256 3556 4312
rect 3233 4254 3556 4256
rect 3233 4251 3299 4254
rect 3550 4252 3556 4254
rect 3620 4252 3626 4316
rect 9070 4252 9076 4316
rect 9140 4314 9146 4316
rect 9305 4314 9371 4317
rect 9140 4312 9371 4314
rect 9140 4256 9310 4312
rect 9366 4256 9371 4312
rect 9140 4254 9371 4256
rect 9140 4252 9146 4254
rect 3558 4178 3618 4252
rect 9305 4251 9371 4254
rect 7557 4178 7623 4181
rect 8109 4178 8175 4181
rect 3558 4118 4768 4178
rect 4708 4045 4768 4118
rect 7557 4176 8175 4178
rect 7557 4120 7562 4176
rect 7618 4120 8114 4176
rect 8170 4120 8175 4176
rect 7557 4118 8175 4120
rect 7557 4115 7623 4118
rect 8109 4115 8175 4118
rect 2313 4042 2379 4045
rect 4521 4042 4587 4045
rect 2313 4040 4587 4042
rect 2313 3984 2318 4040
rect 2374 3984 4526 4040
rect 4582 3984 4587 4040
rect 2313 3982 4587 3984
rect 2313 3979 2379 3982
rect 4521 3979 4587 3982
rect 4705 4040 4771 4045
rect 8017 4042 8083 4045
rect 4705 3984 4710 4040
rect 4766 3984 4771 4040
rect 4705 3979 4771 3984
rect 5398 4040 8083 4042
rect 5398 3984 8022 4040
rect 8078 3984 8083 4040
rect 5398 3982 8083 3984
rect 4153 3906 4219 3909
rect 5206 3906 5212 3908
rect 4153 3904 5212 3906
rect 4153 3848 4158 3904
rect 4214 3848 5212 3904
rect 4153 3846 5212 3848
rect 4153 3843 4219 3846
rect 5206 3844 5212 3846
rect 5276 3844 5282 3908
rect 2820 3840 3136 3841
rect 0 3770 800 3800
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 1853 3770 1919 3773
rect 0 3768 1919 3770
rect 0 3712 1858 3768
rect 1914 3712 1919 3768
rect 0 3710 1919 3712
rect 0 3680 800 3710
rect 1853 3707 1919 3710
rect 4153 3770 4219 3773
rect 5398 3770 5458 3982
rect 8017 3979 8083 3982
rect 11329 3906 11395 3909
rect 13721 3906 13787 3909
rect 11329 3904 13787 3906
rect 11329 3848 11334 3904
rect 11390 3848 13726 3904
rect 13782 3848 13787 3904
rect 11329 3846 13787 3848
rect 11329 3843 11395 3846
rect 13721 3843 13787 3846
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 9305 3772 9371 3773
rect 4153 3768 5458 3770
rect 4153 3712 4158 3768
rect 4214 3712 5458 3768
rect 4153 3710 5458 3712
rect 4153 3707 4219 3710
rect 9254 3708 9260 3772
rect 9324 3770 9371 3772
rect 9324 3768 9416 3770
rect 9366 3712 9416 3768
rect 9324 3710 9416 3712
rect 9324 3708 9371 3710
rect 12566 3708 12572 3772
rect 12636 3770 12642 3772
rect 12709 3770 12775 3773
rect 12636 3768 12775 3770
rect 12636 3712 12714 3768
rect 12770 3712 12775 3768
rect 12636 3710 12775 3712
rect 12636 3708 12642 3710
rect 9305 3707 9371 3708
rect 12709 3707 12775 3710
rect 3693 3634 3759 3637
rect 7557 3634 7623 3637
rect 3693 3632 7623 3634
rect 3693 3576 3698 3632
rect 3754 3576 7562 3632
rect 7618 3576 7623 3632
rect 3693 3574 7623 3576
rect 3693 3571 3759 3574
rect 7557 3571 7623 3574
rect 10133 3634 10199 3637
rect 12014 3634 12020 3636
rect 10133 3632 12020 3634
rect 10133 3576 10138 3632
rect 10194 3576 12020 3632
rect 10133 3574 12020 3576
rect 10133 3571 10199 3574
rect 12014 3572 12020 3574
rect 12084 3572 12090 3636
rect 4521 3498 4587 3501
rect 10869 3498 10935 3501
rect 4521 3496 10935 3498
rect 4521 3440 4526 3496
rect 4582 3440 10874 3496
rect 10930 3440 10935 3496
rect 4521 3438 10935 3440
rect 4521 3435 4587 3438
rect 10869 3435 10935 3438
rect 9673 3362 9739 3365
rect 11237 3364 11303 3365
rect 11237 3362 11284 3364
rect 9673 3360 11284 3362
rect 9673 3304 9678 3360
rect 9734 3304 11242 3360
rect 9673 3302 11284 3304
rect 9673 3299 9739 3302
rect 11237 3300 11284 3302
rect 11348 3300 11354 3364
rect 16205 3362 16271 3365
rect 16400 3362 17200 3392
rect 16205 3360 17200 3362
rect 16205 3304 16210 3360
rect 16266 3304 17200 3360
rect 16205 3302 17200 3304
rect 11237 3299 11303 3300
rect 16205 3299 16271 3302
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 16400 3272 17200 3302
rect 12190 3231 12506 3232
rect 10869 3226 10935 3229
rect 10869 3224 12082 3226
rect 10869 3168 10874 3224
rect 10930 3168 12082 3224
rect 10869 3166 12082 3168
rect 10869 3163 10935 3166
rect 4153 3090 4219 3093
rect 11329 3090 11395 3093
rect 4153 3088 11395 3090
rect 4153 3032 4158 3088
rect 4214 3032 11334 3088
rect 11390 3032 11395 3088
rect 4153 3030 11395 3032
rect 12022 3090 12082 3166
rect 12157 3090 12223 3093
rect 12801 3090 12867 3093
rect 12022 3088 12867 3090
rect 12022 3032 12162 3088
rect 12218 3032 12806 3088
rect 12862 3032 12867 3088
rect 12022 3030 12867 3032
rect 4153 3027 4219 3030
rect 11329 3027 11395 3030
rect 12157 3027 12223 3030
rect 12801 3027 12867 3030
rect 13854 3028 13860 3092
rect 13924 3090 13930 3092
rect 14181 3090 14247 3093
rect 13924 3088 14247 3090
rect 13924 3032 14186 3088
rect 14242 3032 14247 3088
rect 13924 3030 14247 3032
rect 13924 3028 13930 3030
rect 14181 3027 14247 3030
rect 7005 2954 7071 2957
rect 15377 2954 15443 2957
rect 7005 2952 15443 2954
rect 7005 2896 7010 2952
rect 7066 2896 15382 2952
rect 15438 2896 15443 2952
rect 7005 2894 15443 2896
rect 7005 2891 7071 2894
rect 15377 2891 15443 2894
rect 0 2818 800 2848
rect 1853 2818 1919 2821
rect 0 2816 1919 2818
rect 0 2760 1858 2816
rect 1914 2760 1919 2816
rect 0 2758 1919 2760
rect 0 2728 800 2758
rect 1853 2755 1919 2758
rect 3233 2818 3299 2821
rect 3969 2818 4035 2821
rect 3233 2816 4035 2818
rect 3233 2760 3238 2816
rect 3294 2760 3974 2816
rect 4030 2760 4035 2816
rect 3233 2758 4035 2760
rect 3233 2755 3299 2758
rect 3969 2755 4035 2758
rect 4613 2818 4679 2821
rect 5073 2818 5139 2821
rect 4613 2816 5139 2818
rect 4613 2760 4618 2816
rect 4674 2760 5078 2816
rect 5134 2760 5139 2816
rect 4613 2758 5139 2760
rect 4613 2755 4679 2758
rect 5073 2755 5139 2758
rect 11513 2818 11579 2821
rect 12157 2818 12223 2821
rect 11513 2816 12223 2818
rect 11513 2760 11518 2816
rect 11574 2760 12162 2816
rect 12218 2760 12223 2816
rect 11513 2758 12223 2760
rect 11513 2755 11579 2758
rect 12157 2755 12223 2758
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 5073 2546 5139 2549
rect 8937 2546 9003 2549
rect 5073 2544 9003 2546
rect 5073 2488 5078 2544
rect 5134 2488 8942 2544
rect 8998 2488 9003 2544
rect 5073 2486 9003 2488
rect 5073 2483 5139 2486
rect 8937 2483 9003 2486
rect 4613 2410 4679 2413
rect 14181 2410 14247 2413
rect 4613 2408 14247 2410
rect 4613 2352 4618 2408
rect 4674 2352 14186 2408
rect 14242 2352 14247 2408
rect 4613 2350 14247 2352
rect 4613 2347 4679 2350
rect 14181 2347 14247 2350
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 5206 1940 5212 2004
rect 5276 2002 5282 2004
rect 8661 2002 8727 2005
rect 5276 2000 8727 2002
rect 5276 1944 8666 2000
rect 8722 1944 8727 2000
rect 5276 1942 8727 1944
rect 5276 1940 5282 1942
rect 8661 1939 8727 1942
rect 0 1866 800 1896
rect 1761 1866 1827 1869
rect 0 1864 1827 1866
rect 0 1808 1766 1864
rect 1822 1808 1827 1864
rect 0 1806 1827 1808
rect 0 1776 800 1806
rect 1761 1803 1827 1806
rect 7966 1804 7972 1868
rect 8036 1866 8042 1868
rect 9489 1866 9555 1869
rect 8036 1864 9555 1866
rect 8036 1808 9494 1864
rect 9550 1808 9555 1864
rect 8036 1806 9555 1808
rect 8036 1804 8042 1806
rect 9489 1803 9555 1806
rect 0 914 800 944
rect 3785 914 3851 917
rect 0 912 3851 914
rect 0 856 3790 912
rect 3846 856 3851 912
rect 0 854 3851 856
rect 0 824 800 854
rect 3785 851 3851 854
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 3556 17036 3620 17100
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 13676 16280 13740 16284
rect 13676 16224 13690 16280
rect 13690 16224 13740 16280
rect 13676 16220 13740 16224
rect 5212 15812 5276 15876
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 12572 15676 12636 15740
rect 12940 15676 13004 15740
rect 9076 15540 9140 15604
rect 14780 15540 14844 15604
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 13860 14452 13924 14516
rect 3372 14180 3436 14244
rect 9444 14180 9508 14244
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 9628 13772 9692 13836
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 11652 13364 11716 13428
rect 13860 13364 13924 13428
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 9812 12684 9876 12748
rect 14964 12744 15028 12748
rect 14964 12688 15014 12744
rect 15014 12688 15028 12744
rect 14964 12684 15028 12688
rect 8156 12548 8220 12612
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 14780 12336 14844 12340
rect 14780 12280 14830 12336
rect 14830 12280 14844 12336
rect 14780 12276 14844 12280
rect 12020 12140 12084 12204
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 13676 11792 13740 11796
rect 13676 11736 13690 11792
rect 13690 11736 13740 11792
rect 13676 11732 13740 11736
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 8892 11188 8956 11252
rect 9628 11188 9692 11252
rect 13676 11188 13740 11252
rect 12572 11052 12636 11116
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 3556 10644 3620 10708
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 9076 10236 9140 10300
rect 13676 10100 13740 10164
rect 14964 9828 15028 9892
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 11284 9556 11348 9620
rect 14780 9556 14844 9620
rect 12572 9420 12636 9484
rect 14596 9420 14660 9484
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 11836 9148 11900 9212
rect 8156 9012 8220 9076
rect 9628 9012 9692 9076
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 3556 8604 3620 8668
rect 3556 8468 3620 8532
rect 8892 8468 8956 8532
rect 13860 8604 13924 8668
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 13860 7788 13924 7852
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 11652 7032 11716 7036
rect 11652 6976 11666 7032
rect 11666 6976 11716 7032
rect 11652 6972 11716 6976
rect 14780 6760 14844 6764
rect 14780 6704 14830 6760
rect 14830 6704 14844 6760
rect 14780 6700 14844 6704
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 14596 6428 14660 6492
rect 9628 6292 9692 6356
rect 9076 6020 9140 6084
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 9260 5884 9324 5948
rect 12020 5748 12084 5812
rect 5212 5612 5276 5676
rect 7972 5672 8036 5676
rect 7972 5616 7986 5672
rect 7986 5616 8036 5672
rect 7972 5612 8036 5616
rect 11836 5612 11900 5676
rect 12940 5612 13004 5676
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 9444 5068 9508 5132
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 5212 4796 5276 4860
rect 9812 4856 9876 4860
rect 9812 4800 9862 4856
rect 9862 4800 9876 4856
rect 9812 4796 9876 4800
rect 3372 4720 3436 4724
rect 3372 4664 3386 4720
rect 3386 4664 3436 4720
rect 3372 4660 3436 4664
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 3556 4252 3620 4316
rect 9076 4252 9140 4316
rect 5212 3844 5276 3908
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 9260 3768 9324 3772
rect 9260 3712 9310 3768
rect 9310 3712 9324 3768
rect 9260 3708 9324 3712
rect 12572 3708 12636 3772
rect 12020 3572 12084 3636
rect 11284 3360 11348 3364
rect 11284 3304 11298 3360
rect 11298 3304 11348 3360
rect 11284 3300 11348 3304
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 13860 3028 13924 3092
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
rect 5212 1940 5276 2004
rect 7972 1804 8036 1868
<< metal4 >>
rect 2818 16896 3138 17456
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 3555 17100 3621 17101
rect 3555 17036 3556 17100
rect 3620 17036 3621 17100
rect 3555 17035 3621 17036
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 3371 14244 3437 14245
rect 3371 14180 3372 14244
rect 3436 14180 3437 14244
rect 3371 14179 3437 14180
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 3374 4725 3434 14179
rect 3558 10709 3618 17035
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 5211 15876 5277 15877
rect 5211 15812 5212 15876
rect 5276 15812 5277 15876
rect 5211 15811 5277 15812
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 3555 10708 3621 10709
rect 3555 10644 3556 10708
rect 3620 10644 3621 10708
rect 3555 10643 3621 10644
rect 3558 8669 3618 10643
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 3555 8668 3621 8669
rect 3555 8604 3556 8668
rect 3620 8604 3621 8668
rect 3555 8603 3621 8604
rect 3555 8532 3621 8533
rect 3555 8468 3556 8532
rect 3620 8468 3621 8532
rect 3555 8467 3621 8468
rect 3371 4724 3437 4725
rect 3371 4660 3372 4724
rect 3436 4660 3437 4724
rect 3371 4659 3437 4660
rect 3558 4317 3618 8467
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 5214 5677 5274 15811
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 10314 16896 10634 17456
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 9075 15604 9141 15605
rect 9075 15540 9076 15604
rect 9140 15540 9141 15604
rect 9075 15539 9141 15540
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8155 12612 8221 12613
rect 8155 12548 8156 12612
rect 8220 12548 8221 12612
rect 8155 12547 8221 12548
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 8158 9077 8218 12547
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8891 11252 8957 11253
rect 8891 11188 8892 11252
rect 8956 11188 8957 11252
rect 8891 11187 8957 11188
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8155 9076 8221 9077
rect 8155 9012 8156 9076
rect 8220 9012 8221 9076
rect 8155 9011 8221 9012
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 5211 5676 5277 5677
rect 5211 5612 5212 5676
rect 5276 5612 5277 5676
rect 5211 5611 5277 5612
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 5214 4861 5274 5611
rect 6566 4928 6886 5952
rect 8440 8736 8760 9760
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8894 8533 8954 11187
rect 9078 10301 9138 15539
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 9443 14244 9509 14245
rect 9443 14180 9444 14244
rect 9508 14180 9509 14244
rect 9443 14179 9509 14180
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 8891 8532 8957 8533
rect 8891 8468 8892 8532
rect 8956 8468 8957 8532
rect 8891 8467 8957 8468
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 7971 5676 8037 5677
rect 7971 5612 7972 5676
rect 8036 5612 8037 5676
rect 7971 5611 8037 5612
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 5211 4860 5277 4861
rect 5211 4796 5212 4860
rect 5276 4796 5277 4860
rect 5211 4795 5277 4796
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 3555 4316 3621 4317
rect 3555 4252 3556 4316
rect 3620 4252 3621 4316
rect 3555 4251 3621 4252
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 4692 3296 5012 4320
rect 5211 3908 5277 3909
rect 5211 3844 5212 3908
rect 5276 3844 5277 3908
rect 5211 3843 5277 3844
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 2208 5012 3232
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 5214 2005 5274 3843
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2128 6886 2688
rect 5211 2004 5277 2005
rect 5211 1940 5212 2004
rect 5276 1940 5277 2004
rect 5211 1939 5277 1940
rect 7974 1869 8034 5611
rect 8440 5472 8760 6496
rect 9075 6084 9141 6085
rect 9075 6020 9076 6084
rect 9140 6020 9141 6084
rect 9075 6019 9141 6020
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 9078 4317 9138 6019
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 9075 4316 9141 4317
rect 9075 4252 9076 4316
rect 9140 4252 9141 4316
rect 9075 4251 9141 4252
rect 9262 3773 9322 5883
rect 9446 5133 9506 14179
rect 9627 13836 9693 13837
rect 9627 13772 9628 13836
rect 9692 13772 9693 13836
rect 9627 13771 9693 13772
rect 9630 11253 9690 13771
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 9811 12748 9877 12749
rect 9811 12684 9812 12748
rect 9876 12684 9877 12748
rect 9811 12683 9877 12684
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 9630 6357 9690 9011
rect 9627 6356 9693 6357
rect 9627 6292 9628 6356
rect 9692 6292 9693 6356
rect 9627 6291 9693 6292
rect 9443 5132 9509 5133
rect 9443 5068 9444 5132
rect 9508 5068 9509 5132
rect 9443 5067 9509 5068
rect 9814 4861 9874 12683
rect 10314 12544 10634 13568
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 13675 16284 13741 16285
rect 13675 16220 13676 16284
rect 13740 16220 13741 16284
rect 13675 16219 13741 16220
rect 12571 15740 12637 15741
rect 12571 15676 12572 15740
rect 12636 15676 12637 15740
rect 12571 15675 12637 15676
rect 12939 15740 13005 15741
rect 12939 15676 12940 15740
rect 13004 15676 13005 15740
rect 12939 15675 13005 15676
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 11651 13428 11717 13429
rect 11651 13364 11652 13428
rect 11716 13364 11717 13428
rect 11651 13363 11717 13364
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 9280 10634 10304
rect 11283 9620 11349 9621
rect 11283 9556 11284 9620
rect 11348 9556 11349 9620
rect 11283 9555 11349 9556
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 9259 3772 9325 3773
rect 9259 3708 9260 3772
rect 9324 3708 9325 3772
rect 9259 3707 9325 3708
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2752 10634 3776
rect 11286 3365 11346 9555
rect 11654 7037 11714 13363
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12019 12204 12085 12205
rect 12019 12140 12020 12204
rect 12084 12140 12085 12204
rect 12019 12139 12085 12140
rect 11835 9212 11901 9213
rect 11835 9148 11836 9212
rect 11900 9148 11901 9212
rect 11835 9147 11901 9148
rect 11651 7036 11717 7037
rect 11651 6972 11652 7036
rect 11716 6972 11717 7036
rect 11651 6971 11717 6972
rect 11838 5677 11898 9147
rect 12022 5813 12082 12139
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12574 11117 12634 15675
rect 12571 11116 12637 11117
rect 12571 11052 12572 11116
rect 12636 11052 12637 11116
rect 12571 11051 12637 11052
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12571 9484 12637 9485
rect 12571 9420 12572 9484
rect 12636 9420 12637 9484
rect 12571 9419 12637 9420
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12019 5812 12085 5813
rect 12019 5748 12020 5812
rect 12084 5748 12085 5812
rect 12019 5747 12085 5748
rect 11835 5676 11901 5677
rect 11835 5612 11836 5676
rect 11900 5612 11901 5676
rect 11835 5611 11901 5612
rect 12022 3637 12082 5747
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12019 3636 12085 3637
rect 12019 3572 12020 3636
rect 12084 3572 12085 3636
rect 12019 3571 12085 3572
rect 11283 3364 11349 3365
rect 11283 3300 11284 3364
rect 11348 3300 11349 3364
rect 11283 3299 11349 3300
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 3296 12508 4320
rect 12574 3773 12634 9419
rect 12942 5677 13002 15675
rect 13678 11797 13738 16219
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14779 15604 14845 15605
rect 14779 15540 14780 15604
rect 14844 15540 14845 15604
rect 14779 15539 14845 15540
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 13859 14516 13925 14517
rect 13859 14452 13860 14516
rect 13924 14452 13925 14516
rect 13859 14451 13925 14452
rect 13862 13429 13922 14451
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 13859 13428 13925 13429
rect 13859 13364 13860 13428
rect 13924 13364 13925 13428
rect 13859 13363 13925 13364
rect 13675 11796 13741 11797
rect 13675 11732 13676 11796
rect 13740 11732 13741 11796
rect 13675 11731 13741 11732
rect 13678 11253 13738 11731
rect 13675 11252 13741 11253
rect 13675 11188 13676 11252
rect 13740 11188 13741 11252
rect 13675 11187 13741 11188
rect 13678 10165 13738 11187
rect 13675 10164 13741 10165
rect 13675 10100 13676 10164
rect 13740 10100 13741 10164
rect 13675 10099 13741 10100
rect 13862 8669 13922 13363
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14782 12341 14842 15539
rect 14963 12748 15029 12749
rect 14963 12684 14964 12748
rect 15028 12684 15029 12748
rect 14963 12683 15029 12684
rect 14779 12340 14845 12341
rect 14779 12276 14780 12340
rect 14844 12276 14845 12340
rect 14779 12275 14845 12276
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 9280 14382 10304
rect 14966 9893 15026 12683
rect 14963 9892 15029 9893
rect 14963 9828 14964 9892
rect 15028 9828 15029 9892
rect 14963 9827 15029 9828
rect 14779 9620 14845 9621
rect 14779 9556 14780 9620
rect 14844 9556 14845 9620
rect 14779 9555 14845 9556
rect 14595 9484 14661 9485
rect 14595 9420 14596 9484
rect 14660 9420 14661 9484
rect 14595 9419 14661 9420
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 13859 8668 13925 8669
rect 13859 8604 13860 8668
rect 13924 8604 13925 8668
rect 13859 8603 13925 8604
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 13859 7852 13925 7853
rect 13859 7788 13860 7852
rect 13924 7788 13925 7852
rect 13859 7787 13925 7788
rect 12939 5676 13005 5677
rect 12939 5612 12940 5676
rect 13004 5612 13005 5676
rect 12939 5611 13005 5612
rect 12571 3772 12637 3773
rect 12571 3708 12572 3772
rect 12636 3708 12637 3772
rect 12571 3707 12637 3708
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 13862 3093 13922 7787
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14598 6493 14658 9419
rect 14782 6765 14842 9555
rect 14779 6764 14845 6765
rect 14779 6700 14780 6764
rect 14844 6700 14845 6764
rect 14779 6699 14845 6700
rect 14595 6492 14661 6493
rect 14595 6428 14596 6492
rect 14660 6428 14661 6492
rect 14595 6427 14661 6428
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 13859 3092 13925 3093
rect 13859 3028 13860 3092
rect 13924 3028 13925 3092
rect 13859 3027 13925 3028
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
rect 7971 1868 8037 1869
rect 7971 1804 7972 1868
rect 8036 1804 8037 1868
rect 7971 1803 8037 1804
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1649977179
transform 1 0 3128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1649977179
transform -1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform 1 0 2576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform -1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform -1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform -1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform -1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 6164 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 7176 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_S_FTB01_A
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 12696 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_S_FTB01_A
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform -1 0 7544 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3864 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4968 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5152 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 10396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15732 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13248 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1649977179
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform -1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1649977179
transform -1 0 15640 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_S_FTB01_A
timestamp 1649977179
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1649977179
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1649977179
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_104
timestamp 1649977179
transform 1 0 10672 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 1649977179
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_46
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_91
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_132
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_42
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_68
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_121
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_138
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_31
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_111
timestamp 1649977179
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_130
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_81
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_16
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_104
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_140
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_154
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_67
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1649977179
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1649977179
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_76
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1649977179
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1649977179
transform 1 0 5428 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_151
timestamp 1649977179
transform 1 0 14996 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_18
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1649977179
transform 1 0 12788 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_130
timestamp 1649977179
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_49
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_72
timestamp 1649977179
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_10
timestamp 1649977179
transform 1 0 2024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_14
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_42
timestamp 1649977179
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_54
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_66
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_156
timestamp 1649977179
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_16
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_77
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_101
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_122
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_13
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_87
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_124
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_132
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_142
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_154
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_158
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_128
timestamp 1649977179
transform 1 0 12880 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_10
timestamp 1649977179
transform 1 0 2024 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_36
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_68
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_109
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_31
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_43
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_18
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_37
timestamp 1649977179
transform 1 0 4508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_122
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_142
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_105
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1649977179
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1649977179
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_61
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_70
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1649977179
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_91
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_102
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1649977179
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_21
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_39
timestamp 1649977179
transform 1 0 4692 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1649977179
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_20
timestamp 1649977179
transform 1 0 2944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_41
timestamp 1649977179
transform 1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_63
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_98
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_128
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_143
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1649977179
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1649977179
transform -1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1649977179
transform -1 0 1932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _16_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1649977179
transform -1 0 13984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform -1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _32_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1649977179
transform -1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform -1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 4692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform -1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform -1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform -1 0 5980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform -1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform -1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform -1 0 6992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform -1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform -1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform -1 0 10304 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform -1 0 11868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform -1 0 11776 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 12512 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5796 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8740 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 4324 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9476 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4876 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7728 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10948 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8188 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2944 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4324 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10672 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5244 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3956 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4324 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6716 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3312 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8832 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6900 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11132 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10856 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8832 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4324 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9292 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7636 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10120 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8096 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3864 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5244 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2944 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13156 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11960 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12420 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13064 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5336 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 4968 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8280 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10764 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12788 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 1472 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2392 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13892 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13248 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1564 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1472 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14996 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11776 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11960 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13248 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2760 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14536 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12880 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform -1 0 2024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform -1 0 14628 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 15456 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 590 592
<< labels >>
flabel metal3 s 16400 16600 17200 16720 0 FreeSans 480 0 0 0 Test_en_E_in
port 0 nsew signal input
flabel metal3 s 16400 9936 17200 10056 0 FreeSans 480 0 0 0 Test_en_E_out
port 1 nsew signal tristate
flabel metal2 s 2134 19200 2190 20000 0 FreeSans 224 90 0 0 Test_en_N_out
port 2 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 3 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 Test_en_W_in
port 4 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 Test_en_W_out
port 5 nsew signal tristate
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 6 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 7 nsew power bidirectional
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 ccff_head
port 8 nsew signal input
flabel metal3 s 16400 3272 17200 3392 0 FreeSans 480 0 0 0 ccff_tail
port 9 nsew signal tristate
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 10 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 11 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 12 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 13 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 14 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 15 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 16 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 17 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 18 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 19 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 20 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 21 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 22 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 23 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 24 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 25 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 26 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 27 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 28 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 29 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 30 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 31 nsew signal tristate
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 32 nsew signal tristate
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 33 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 34 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 35 nsew signal tristate
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 36 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 37 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 38 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 39 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 40 nsew signal tristate
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 41 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 42 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 43 nsew signal tristate
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 44 nsew signal tristate
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 45 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 46 nsew signal tristate
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 47 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 48 nsew signal tristate
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 49 nsew signal tristate
flabel metal2 s 9862 19200 9918 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 50 nsew signal input
flabel metal2 s 13542 19200 13598 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 51 nsew signal input
flabel metal2 s 13910 19200 13966 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 52 nsew signal input
flabel metal2 s 14278 19200 14334 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 53 nsew signal input
flabel metal2 s 14646 19200 14702 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 54 nsew signal input
flabel metal2 s 15014 19200 15070 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 55 nsew signal input
flabel metal2 s 15382 19200 15438 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 56 nsew signal input
flabel metal2 s 15750 19200 15806 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 57 nsew signal input
flabel metal2 s 16118 19200 16174 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 58 nsew signal input
flabel metal2 s 16486 19200 16542 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 59 nsew signal input
flabel metal2 s 16854 19200 16910 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 60 nsew signal input
flabel metal2 s 10230 19200 10286 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 61 nsew signal input
flabel metal2 s 10598 19200 10654 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 62 nsew signal input
flabel metal2 s 10966 19200 11022 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 63 nsew signal input
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 64 nsew signal input
flabel metal2 s 11702 19200 11758 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 65 nsew signal input
flabel metal2 s 12070 19200 12126 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 66 nsew signal input
flabel metal2 s 12438 19200 12494 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 67 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 68 nsew signal input
flabel metal2 s 13174 19200 13230 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 69 nsew signal input
flabel metal2 s 2502 19200 2558 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 70 nsew signal tristate
flabel metal2 s 6182 19200 6238 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 71 nsew signal tristate
flabel metal2 s 6550 19200 6606 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 72 nsew signal tristate
flabel metal2 s 6918 19200 6974 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 73 nsew signal tristate
flabel metal2 s 7286 19200 7342 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 74 nsew signal tristate
flabel metal2 s 7654 19200 7710 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 75 nsew signal tristate
flabel metal2 s 8022 19200 8078 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 76 nsew signal tristate
flabel metal2 s 8390 19200 8446 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 77 nsew signal tristate
flabel metal2 s 8758 19200 8814 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 78 nsew signal tristate
flabel metal2 s 9126 19200 9182 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 79 nsew signal tristate
flabel metal2 s 9494 19200 9550 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 80 nsew signal tristate
flabel metal2 s 2870 19200 2926 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 81 nsew signal tristate
flabel metal2 s 3238 19200 3294 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 82 nsew signal tristate
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 83 nsew signal tristate
flabel metal2 s 3974 19200 4030 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 84 nsew signal tristate
flabel metal2 s 4342 19200 4398 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 85 nsew signal tristate
flabel metal2 s 4710 19200 4766 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 86 nsew signal tristate
flabel metal2 s 5078 19200 5134 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 87 nsew signal tristate
flabel metal2 s 5446 19200 5502 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 88 nsew signal tristate
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 89 nsew signal tristate
flabel metal2 s 294 19200 350 20000 0 FreeSans 224 90 0 0 clk_2_N_out
port 90 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 clk_2_S_in
port 91 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 clk_2_S_out
port 92 nsew signal tristate
flabel metal2 s 662 19200 718 20000 0 FreeSans 224 90 0 0 clk_3_N_out
port 93 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 clk_3_S_in
port 94 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 clk_3_S_out
port 95 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_grid_pin_16_
port 96 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 left_grid_pin_17_
port 97 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_grid_pin_18_
port 98 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 left_grid_pin_19_
port 99 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 left_grid_pin_20_
port 100 nsew signal tristate
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 left_grid_pin_21_
port 101 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 left_grid_pin_22_
port 102 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 left_grid_pin_23_
port 103 nsew signal tristate
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 left_grid_pin_24_
port 104 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 left_grid_pin_25_
port 105 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 left_grid_pin_26_
port 106 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 left_grid_pin_27_
port 107 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 left_grid_pin_28_
port 108 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 left_grid_pin_29_
port 109 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 left_grid_pin_30_
port 110 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 left_grid_pin_31_
port 111 nsew signal tristate
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 112 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 113 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 prog_clk_0_W_in
port 114 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 prog_clk_2_N_out
port 115 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 prog_clk_2_S_in
port 116 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 prog_clk_2_S_out
port 117 nsew signal tristate
flabel metal2 s 1766 19200 1822 20000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 118 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 prog_clk_3_S_in
port 119 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 prog_clk_3_S_out
port 120 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
