magic
tech sky130A
magscale 1 2
timestamp 1682507234
<< viali >>
rect 1777 24361 1811 24395
rect 24409 24361 24443 24395
rect 18153 24293 18187 24327
rect 3249 24225 3283 24259
rect 6561 24225 6595 24259
rect 8217 24225 8251 24259
rect 12817 24225 12851 24259
rect 18705 24225 18739 24259
rect 25053 24225 25087 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9873 24157 9907 24191
rect 10977 24157 11011 24191
rect 12357 24157 12391 24191
rect 14289 24157 14323 24191
rect 15393 24157 15427 24191
rect 16865 24157 16899 24191
rect 18613 24157 18647 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 24961 24157 24995 24191
rect 1593 24089 1627 24123
rect 5825 24089 5859 24123
rect 9045 24089 9079 24123
rect 17509 24089 17543 24123
rect 18521 24089 18555 24123
rect 21005 24089 21039 24123
rect 21925 24089 21959 24123
rect 22477 24089 22511 24123
rect 3985 24021 4019 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14933 24021 14967 24055
rect 16037 24021 16071 24055
rect 16313 24021 16347 24055
rect 17785 24021 17819 24055
rect 19441 24021 19475 24055
rect 22109 24021 22143 24055
rect 23949 24021 23983 24055
rect 24593 24021 24627 24055
rect 6561 23817 6595 23851
rect 14105 23817 14139 23851
rect 14565 23817 14599 23851
rect 20361 23817 20395 23851
rect 20729 23817 20763 23851
rect 22201 23817 22235 23851
rect 24409 23817 24443 23851
rect 25053 23817 25087 23851
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 16221 23749 16255 23783
rect 21557 23749 21591 23783
rect 21833 23749 21867 23783
rect 22569 23749 22603 23783
rect 24961 23749 24995 23783
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 6825 23681 6859 23715
rect 7481 23681 7515 23715
rect 7941 23681 7975 23715
rect 9781 23681 9815 23715
rect 12081 23681 12115 23715
rect 14473 23681 14507 23715
rect 15577 23681 15611 23715
rect 16957 23681 16991 23715
rect 1777 23613 1811 23647
rect 5825 23613 5859 23647
rect 12541 23613 12575 23647
rect 14749 23613 14783 23647
rect 18061 23613 18095 23647
rect 18337 23613 18371 23647
rect 20821 23613 20855 23647
rect 20913 23613 20947 23647
rect 22293 23613 22327 23647
rect 25145 23613 25179 23647
rect 2329 23545 2363 23579
rect 11529 23477 11563 23511
rect 11805 23477 11839 23511
rect 13829 23477 13863 23511
rect 15209 23477 15243 23511
rect 17601 23477 17635 23511
rect 19809 23477 19843 23511
rect 21373 23477 21407 23511
rect 24041 23477 24075 23511
rect 24593 23477 24627 23511
rect 9321 23273 9355 23307
rect 14473 23273 14507 23307
rect 18337 23273 18371 23307
rect 18613 23273 18647 23307
rect 21189 23205 21223 23239
rect 3249 23137 3283 23171
rect 6561 23137 6595 23171
rect 8217 23137 8251 23171
rect 10517 23137 10551 23171
rect 15301 23137 15335 23171
rect 17785 23137 17819 23171
rect 19717 23137 19751 23171
rect 21649 23137 21683 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 4261 23069 4295 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 9965 23069 9999 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 1593 23001 1627 23035
rect 9229 23001 9263 23035
rect 12633 23001 12667 23035
rect 14381 23001 14415 23035
rect 17693 23001 17727 23035
rect 18521 23001 18555 23035
rect 21925 23001 21959 23035
rect 24961 23001 24995 23035
rect 1777 22933 1811 22967
rect 3893 22933 3927 22967
rect 4905 22933 4939 22967
rect 13553 22933 13587 22967
rect 16773 22933 16807 22967
rect 17233 22933 17267 22967
rect 18981 22933 19015 22967
rect 23397 22933 23431 22967
rect 23857 22933 23891 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 13093 22729 13127 22763
rect 15393 22729 15427 22763
rect 20269 22729 20303 22763
rect 21465 22729 21499 22763
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 8769 22661 8803 22695
rect 15945 22661 15979 22695
rect 17141 22661 17175 22695
rect 19441 22661 19475 22695
rect 22385 22661 22419 22695
rect 23581 22661 23615 22695
rect 1685 22593 1719 22627
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6653 22593 6687 22627
rect 7297 22593 7331 22627
rect 7573 22593 7607 22627
rect 12081 22593 12115 22627
rect 12173 22593 12207 22627
rect 13001 22593 13035 22627
rect 13645 22593 13679 22627
rect 16865 22593 16899 22627
rect 19533 22593 19567 22627
rect 20637 22593 20671 22627
rect 2329 22525 2363 22559
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 11161 22525 11195 22559
rect 12265 22525 12299 22559
rect 13921 22525 13955 22559
rect 19625 22525 19659 22559
rect 20729 22525 20763 22559
rect 20821 22525 20855 22559
rect 22477 22525 22511 22559
rect 22569 22525 22603 22559
rect 23305 22525 23339 22559
rect 11529 22457 11563 22491
rect 16129 22457 16163 22491
rect 19073 22457 19107 22491
rect 25053 22457 25087 22491
rect 6745 22389 6779 22423
rect 11713 22389 11747 22423
rect 16405 22389 16439 22423
rect 18613 22389 18647 22423
rect 21373 22389 21407 22423
rect 22017 22389 22051 22423
rect 25329 22389 25363 22423
rect 14552 22185 14586 22219
rect 18705 22185 18739 22219
rect 20618 22185 20652 22219
rect 16037 22117 16071 22151
rect 1685 22049 1719 22083
rect 2881 22049 2915 22083
rect 6101 22049 6135 22083
rect 8309 22049 8343 22083
rect 10057 22049 10091 22083
rect 10977 22049 11011 22083
rect 14289 22049 14323 22083
rect 17049 22049 17083 22083
rect 18245 22049 18279 22083
rect 23213 22049 23247 22083
rect 24041 22049 24075 22083
rect 25237 22049 25271 22083
rect 2237 21981 2271 22015
rect 4261 21981 4295 22015
rect 5365 21981 5399 22015
rect 7389 21981 7423 22015
rect 10701 21981 10735 22015
rect 13093 21981 13127 22015
rect 18153 21981 18187 22015
rect 19533 21981 19567 22015
rect 20361 21981 20395 22015
rect 23857 21981 23891 22015
rect 24961 21981 24995 22015
rect 9873 21913 9907 21947
rect 16957 21913 16991 21947
rect 18889 21913 18923 21947
rect 19993 21913 20027 21947
rect 23029 21913 23063 21947
rect 1593 21845 1627 21879
rect 3893 21845 3927 21879
rect 4905 21845 4939 21879
rect 8953 21845 8987 21879
rect 9229 21845 9263 21879
rect 9505 21845 9539 21879
rect 9965 21845 9999 21879
rect 12449 21845 12483 21879
rect 12725 21845 12759 21879
rect 13737 21845 13771 21879
rect 16497 21845 16531 21879
rect 16865 21845 16899 21879
rect 17693 21845 17727 21879
rect 18061 21845 18095 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 22569 21845 22603 21879
rect 22937 21845 22971 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 2329 21641 2363 21675
rect 11897 21641 11931 21675
rect 12173 21641 12207 21675
rect 13277 21641 13311 21675
rect 14197 21641 14231 21675
rect 14289 21641 14323 21675
rect 25145 21641 25179 21675
rect 25513 21641 25547 21675
rect 9321 21573 9355 21607
rect 11069 21573 11103 21607
rect 13553 21573 13587 21607
rect 16405 21573 16439 21607
rect 17417 21573 17451 21607
rect 1685 21505 1719 21539
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 7205 21505 7239 21539
rect 9045 21505 9079 21539
rect 11253 21505 11287 21539
rect 11713 21505 11747 21539
rect 12633 21505 12667 21539
rect 15393 21505 15427 21539
rect 16221 21505 16255 21539
rect 16773 21505 16807 21539
rect 18245 21505 18279 21539
rect 20821 21505 20855 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 6561 21437 6595 21471
rect 7665 21437 7699 21471
rect 12725 21437 12759 21471
rect 12817 21437 12851 21471
rect 14473 21437 14507 21471
rect 15485 21437 15519 21471
rect 15577 21437 15611 21471
rect 17509 21437 17543 21471
rect 17601 21437 17635 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 22477 21437 22511 21471
rect 22569 21437 22603 21471
rect 23673 21437 23707 21471
rect 10793 21369 10827 21403
rect 11621 21369 11655 21403
rect 23213 21369 23247 21403
rect 12265 21301 12299 21335
rect 13829 21301 13863 21335
rect 15025 21301 15059 21335
rect 16129 21301 16163 21335
rect 17049 21301 17083 21335
rect 19533 21301 19567 21335
rect 20453 21301 20487 21335
rect 21557 21301 21591 21335
rect 22017 21301 22051 21335
rect 23121 21301 23155 21335
rect 13645 21097 13679 21131
rect 16681 21097 16715 21131
rect 17877 21097 17911 21131
rect 22845 21097 22879 21131
rect 6469 21029 6503 21063
rect 12909 21029 12943 21063
rect 15485 21029 15519 21063
rect 4905 20961 4939 20995
rect 7389 20961 7423 20995
rect 11161 20961 11195 20995
rect 15945 20961 15979 20995
rect 16129 20961 16163 20995
rect 17233 20961 17267 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 21189 20961 21223 20995
rect 22201 20961 22235 20995
rect 23305 20961 23339 20995
rect 23397 20961 23431 20995
rect 25053 20961 25087 20995
rect 25237 20961 25271 20995
rect 2237 20893 2271 20927
rect 2973 20893 3007 20927
rect 4077 20893 4111 20927
rect 5825 20893 5859 20927
rect 7113 20893 7147 20927
rect 8769 20893 8803 20927
rect 9137 20893 9171 20927
rect 9413 20893 9447 20927
rect 10609 20893 10643 20927
rect 13553 20893 13587 20927
rect 14289 20893 14323 20927
rect 19441 20893 19475 20927
rect 22109 20893 22143 20927
rect 23213 20893 23247 20927
rect 1593 20825 1627 20859
rect 11437 20825 11471 20859
rect 18245 20825 18279 20859
rect 19717 20825 19751 20859
rect 24961 20825 24995 20859
rect 1685 20757 1719 20791
rect 10425 20757 10459 20791
rect 14933 20757 14967 20791
rect 15853 20757 15887 20791
rect 17049 20757 17083 20791
rect 17141 20757 17175 20791
rect 18889 20757 18923 20791
rect 21649 20757 21683 20791
rect 22017 20757 22051 20791
rect 23949 20757 23983 20791
rect 24041 20757 24075 20791
rect 24593 20757 24627 20791
rect 6009 20553 6043 20587
rect 7481 20553 7515 20587
rect 18705 20553 18739 20587
rect 23121 20553 23155 20587
rect 8585 20485 8619 20519
rect 11161 20485 11195 20519
rect 11345 20485 11379 20519
rect 11713 20485 11747 20519
rect 12449 20485 12483 20519
rect 16313 20485 16347 20519
rect 17233 20485 17267 20519
rect 22477 20485 22511 20519
rect 1869 20417 1903 20451
rect 3065 20417 3099 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 6469 20417 6503 20451
rect 6837 20417 6871 20451
rect 7929 20417 7963 20451
rect 9045 20417 9079 20451
rect 13185 20417 13219 20451
rect 13553 20417 13587 20451
rect 16129 20417 16163 20451
rect 16957 20417 16991 20451
rect 22569 20417 22603 20451
rect 23489 20417 23523 20451
rect 1593 20349 1627 20383
rect 3341 20349 3375 20383
rect 9321 20349 9355 20383
rect 12541 20349 12575 20383
rect 12633 20349 12667 20383
rect 13829 20349 13863 20383
rect 15301 20349 15335 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 21281 20349 21315 20383
rect 22661 20349 22695 20383
rect 23765 20349 23799 20383
rect 15577 20281 15611 20315
rect 4721 20213 4755 20247
rect 10793 20213 10827 20247
rect 11529 20213 11563 20247
rect 12081 20213 12115 20247
rect 21005 20213 21039 20247
rect 21557 20213 21591 20247
rect 22109 20213 22143 20247
rect 25237 20213 25271 20247
rect 1593 20009 1627 20043
rect 7481 20009 7515 20043
rect 8953 20009 8987 20043
rect 14933 20009 14967 20043
rect 17693 20009 17727 20043
rect 20453 20009 20487 20043
rect 20913 20009 20947 20043
rect 21354 20009 21388 20043
rect 22845 20009 22879 20043
rect 24593 20009 24627 20043
rect 17049 19941 17083 19975
rect 17325 19941 17359 19975
rect 2513 19873 2547 19907
rect 3985 19873 4019 19907
rect 10885 19873 10919 19907
rect 10977 19873 11011 19907
rect 13369 19873 13403 19907
rect 15485 19873 15519 19907
rect 18245 19873 18279 19907
rect 19993 19873 20027 19907
rect 21097 19873 21131 19907
rect 23765 19873 23799 19907
rect 23949 19873 23983 19907
rect 25145 19873 25179 19907
rect 2145 19805 2179 19839
rect 4629 19805 4663 19839
rect 4905 19805 4939 19839
rect 6837 19805 6871 19839
rect 7941 19805 7975 19839
rect 9321 19805 9355 19839
rect 11621 19805 11655 19839
rect 13921 19805 13955 19839
rect 16129 19805 16163 19839
rect 19901 19805 19935 19839
rect 6561 19737 6595 19771
rect 9965 19737 9999 19771
rect 11897 19737 11931 19771
rect 23673 19737 23707 19771
rect 1685 19669 1719 19703
rect 5917 19669 5951 19703
rect 8585 19669 8619 19703
rect 10425 19669 10459 19703
rect 10793 19669 10827 19703
rect 13645 19669 13679 19703
rect 14289 19669 14323 19703
rect 15301 19669 15335 19703
rect 15393 19669 15427 19703
rect 16773 19669 16807 19703
rect 17509 19669 17543 19703
rect 18061 19669 18095 19703
rect 18153 19669 18187 19703
rect 18705 19669 18739 19703
rect 18981 19669 19015 19703
rect 19441 19669 19475 19703
rect 19809 19669 19843 19703
rect 20729 19669 20763 19703
rect 23305 19669 23339 19703
rect 24961 19669 24995 19703
rect 25053 19669 25087 19703
rect 1501 19465 1535 19499
rect 3893 19465 3927 19499
rect 4537 19465 4571 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 19625 19465 19659 19499
rect 20453 19465 20487 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 22477 19465 22511 19499
rect 25053 19465 25087 19499
rect 7481 19397 7515 19431
rect 9321 19397 9355 19431
rect 15393 19397 15427 19431
rect 20821 19397 20855 19431
rect 1961 19329 1995 19363
rect 4077 19329 4111 19363
rect 4721 19329 4755 19363
rect 6009 19329 6043 19363
rect 7941 19329 7975 19363
rect 9045 19329 9079 19363
rect 12081 19329 12115 19363
rect 12725 19329 12759 19363
rect 16129 19329 16163 19363
rect 17049 19329 17083 19363
rect 19717 19329 19751 19363
rect 23305 19329 23339 19363
rect 2237 19261 2271 19295
rect 3617 19261 3651 19295
rect 5365 19261 5399 19295
rect 6929 19261 6963 19295
rect 11621 19261 11655 19295
rect 12265 19261 12299 19295
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 17325 19261 17359 19295
rect 18797 19261 18831 19295
rect 19901 19261 19935 19295
rect 20913 19261 20947 19295
rect 21097 19261 21131 19295
rect 22569 19261 22603 19295
rect 23581 19261 23615 19295
rect 25421 19261 25455 19295
rect 8585 19193 8619 19227
rect 5089 19125 5123 19159
rect 6561 19125 6595 19159
rect 10793 19125 10827 19159
rect 11069 19125 11103 19159
rect 11345 19125 11379 19159
rect 16681 19125 16715 19159
rect 19257 19125 19291 19159
rect 21465 19125 21499 19159
rect 2605 18921 2639 18955
rect 5457 18921 5491 18955
rect 7481 18921 7515 18955
rect 14289 18921 14323 18955
rect 1685 18853 1719 18887
rect 13001 18853 13035 18887
rect 17233 18853 17267 18887
rect 19717 18853 19751 18887
rect 22569 18853 22603 18887
rect 24593 18853 24627 18887
rect 3249 18785 3283 18819
rect 3985 18785 4019 18819
rect 4261 18785 4295 18819
rect 5825 18785 5859 18819
rect 9873 18785 9907 18819
rect 12449 18785 12483 18819
rect 13645 18785 13679 18819
rect 14749 18785 14783 18819
rect 14933 18785 14967 18819
rect 15761 18785 15795 18819
rect 18613 18785 18647 18819
rect 23121 18785 23155 18819
rect 25237 18785 25271 18819
rect 2145 18717 2179 18751
rect 2789 18717 2823 18751
rect 6837 18717 6871 18751
rect 7941 18717 7975 18751
rect 10425 18717 10459 18751
rect 13369 18717 13403 18751
rect 15485 18717 15519 18751
rect 17693 18717 17727 18751
rect 18429 18717 18463 18751
rect 20361 18717 20395 18751
rect 23857 18717 23891 18751
rect 13461 18649 13495 18683
rect 18521 18649 18555 18683
rect 19533 18649 19567 18683
rect 20637 18649 20671 18683
rect 23029 18649 23063 18683
rect 25053 18649 25087 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 5181 18581 5215 18615
rect 6377 18581 6411 18615
rect 8585 18581 8619 18615
rect 9229 18581 9263 18615
rect 9597 18581 9631 18615
rect 9689 18581 9723 18615
rect 11713 18581 11747 18615
rect 12725 18581 12759 18615
rect 14657 18581 14691 18615
rect 17509 18581 17543 18615
rect 18061 18581 18095 18615
rect 20085 18581 20119 18615
rect 22109 18581 22143 18615
rect 22937 18581 22971 18615
rect 23949 18581 23983 18615
rect 24961 18581 24995 18615
rect 10701 18377 10735 18411
rect 11069 18377 11103 18411
rect 11253 18377 11287 18411
rect 14289 18377 14323 18411
rect 15209 18377 15243 18411
rect 23305 18377 23339 18411
rect 25329 18377 25363 18411
rect 5825 18309 5859 18343
rect 6193 18309 6227 18343
rect 9229 18309 9263 18343
rect 13001 18309 13035 18343
rect 15669 18309 15703 18343
rect 16221 18309 16255 18343
rect 18429 18309 18463 18343
rect 20821 18309 20855 18343
rect 21465 18309 21499 18343
rect 22017 18309 22051 18343
rect 24869 18309 24903 18343
rect 25237 18309 25271 18343
rect 1593 18241 1627 18275
rect 2789 18241 2823 18275
rect 3617 18241 3651 18275
rect 4261 18241 4295 18275
rect 4721 18241 4755 18275
rect 4997 18241 5031 18275
rect 6469 18241 6503 18275
rect 6745 18241 6779 18275
rect 7849 18241 7883 18275
rect 8953 18241 8987 18275
rect 12173 18241 12207 18275
rect 15577 18241 15611 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 19625 18241 19659 18275
rect 24225 18241 24259 18275
rect 1869 18173 1903 18207
rect 2973 18173 3007 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 15761 18173 15795 18207
rect 17509 18173 17543 18207
rect 18521 18173 18555 18207
rect 18613 18173 18647 18207
rect 19717 18173 19751 18207
rect 19901 18173 19935 18207
rect 20913 18173 20947 18207
rect 21097 18173 21131 18207
rect 3157 18105 3191 18139
rect 4077 18105 4111 18139
rect 3433 18037 3467 18071
rect 7389 18037 7423 18071
rect 8493 18037 8527 18071
rect 11805 18037 11839 18071
rect 16405 18037 16439 18071
rect 16865 18037 16899 18071
rect 18061 18037 18095 18071
rect 19257 18037 19291 18071
rect 20453 18037 20487 18071
rect 17141 17833 17175 17867
rect 3249 17765 3283 17799
rect 6009 17765 6043 17799
rect 11529 17765 11563 17799
rect 13737 17765 13771 17799
rect 18613 17765 18647 17799
rect 22477 17765 22511 17799
rect 23121 17765 23155 17799
rect 1869 17697 1903 17731
rect 4813 17697 4847 17731
rect 9781 17697 9815 17731
rect 11989 17697 12023 17731
rect 14197 17697 14231 17731
rect 14289 17697 14323 17731
rect 14933 17697 14967 17731
rect 17693 17697 17727 17731
rect 20085 17697 20119 17731
rect 20729 17697 20763 17731
rect 23765 17697 23799 17731
rect 23857 17697 23891 17731
rect 1593 17629 1627 17663
rect 3433 17629 3467 17663
rect 3893 17629 3927 17663
rect 4537 17629 4571 17663
rect 5733 17629 5767 17663
rect 6193 17629 6227 17663
rect 6837 17629 6871 17663
rect 7481 17629 7515 17663
rect 7941 17629 7975 17663
rect 17509 17629 17543 17663
rect 19901 17629 19935 17663
rect 22845 17629 22879 17663
rect 23673 17629 23707 17663
rect 24593 17629 24627 17663
rect 2881 17561 2915 17595
rect 8585 17561 8619 17595
rect 10057 17561 10091 17595
rect 12265 17561 12299 17595
rect 15209 17561 15243 17595
rect 18429 17561 18463 17595
rect 19809 17561 19843 17595
rect 21005 17561 21039 17595
rect 25237 17561 25271 17595
rect 2789 17493 2823 17527
rect 3985 17493 4019 17527
rect 4261 17493 4295 17527
rect 6653 17493 6687 17527
rect 7297 17493 7331 17527
rect 9137 17493 9171 17527
rect 16681 17493 16715 17527
rect 17601 17493 17635 17527
rect 18889 17493 18923 17527
rect 19441 17493 19475 17527
rect 23029 17493 23063 17527
rect 23305 17493 23339 17527
rect 1685 17289 1719 17323
rect 3479 17289 3513 17323
rect 7665 17289 7699 17323
rect 8769 17289 8803 17323
rect 13461 17289 13495 17323
rect 14105 17289 14139 17323
rect 15025 17289 15059 17323
rect 15853 17289 15887 17323
rect 21189 17289 21223 17323
rect 25421 17289 25455 17323
rect 1501 17221 1535 17255
rect 11989 17221 12023 17255
rect 21557 17221 21591 17255
rect 22017 17221 22051 17255
rect 22201 17221 22235 17255
rect 2237 17153 2271 17187
rect 3249 17153 3283 17187
rect 4813 17153 4847 17187
rect 6561 17153 6595 17187
rect 8125 17153 8159 17187
rect 9229 17153 9263 17187
rect 11253 17153 11287 17187
rect 11713 17153 11747 17187
rect 14381 17153 14415 17187
rect 17233 17153 17267 17187
rect 17325 17153 17359 17187
rect 18337 17153 18371 17187
rect 20545 17153 20579 17187
rect 21833 17153 21867 17187
rect 22569 17153 22603 17187
rect 24869 17153 24903 17187
rect 1961 17085 1995 17119
rect 4537 17085 4571 17119
rect 5825 17085 5859 17119
rect 6837 17085 6871 17119
rect 9505 17085 9539 17119
rect 10977 17085 11011 17119
rect 13829 17085 13863 17119
rect 15945 17085 15979 17119
rect 16037 17085 16071 17119
rect 17417 17085 17451 17119
rect 20085 17085 20119 17119
rect 22845 17085 22879 17119
rect 25053 17017 25087 17051
rect 15485 16949 15519 16983
rect 16865 16949 16899 16983
rect 17877 16949 17911 16983
rect 18600 16949 18634 16983
rect 24317 16949 24351 16983
rect 7573 16745 7607 16779
rect 9045 16745 9079 16779
rect 9413 16745 9447 16779
rect 16037 16745 16071 16779
rect 3893 16677 3927 16711
rect 4169 16677 4203 16711
rect 21649 16677 21683 16711
rect 2605 16609 2639 16643
rect 2881 16609 2915 16643
rect 3985 16609 4019 16643
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 6745 16609 6779 16643
rect 8585 16609 8619 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 12265 16609 12299 16643
rect 14289 16609 14323 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 19717 16609 19751 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 1685 16541 1719 16575
rect 2145 16541 2179 16575
rect 4721 16541 4755 16575
rect 6469 16541 6503 16575
rect 8217 16541 8251 16575
rect 8769 16541 8803 16575
rect 9689 16541 9723 16575
rect 11989 16541 12023 16575
rect 16681 16541 16715 16575
rect 17141 16541 17175 16575
rect 21833 16541 21867 16575
rect 24593 16541 24627 16575
rect 14565 16473 14599 16507
rect 1961 16405 1995 16439
rect 4537 16405 4571 16439
rect 8033 16405 8067 16439
rect 9137 16405 9171 16439
rect 10333 16405 10367 16439
rect 10793 16405 10827 16439
rect 11161 16405 11195 16439
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18889 16405 18923 16439
rect 21189 16405 21223 16439
rect 24041 16405 24075 16439
rect 25237 16405 25271 16439
rect 5825 16201 5859 16235
rect 9965 16201 9999 16235
rect 13921 16201 13955 16235
rect 14381 16201 14415 16235
rect 19349 16201 19383 16235
rect 21005 16201 21039 16235
rect 23213 16201 23247 16235
rect 23765 16201 23799 16235
rect 23857 16201 23891 16235
rect 2973 16133 3007 16167
rect 6653 16133 6687 16167
rect 11989 16133 12023 16167
rect 15209 16133 15243 16167
rect 15945 16133 15979 16167
rect 21557 16133 21591 16167
rect 1869 16065 1903 16099
rect 3249 16065 3283 16099
rect 4537 16065 4571 16099
rect 4813 16065 4847 16099
rect 6009 16065 6043 16099
rect 6469 16065 6503 16099
rect 7297 16065 7331 16099
rect 8309 16065 8343 16099
rect 8861 16065 8895 16099
rect 9321 16065 9355 16099
rect 10793 16065 10827 16099
rect 14289 16065 14323 16099
rect 14933 16065 14967 16099
rect 15853 16065 15887 16099
rect 17141 16065 17175 16099
rect 19717 16065 19751 16099
rect 19809 16065 19843 16099
rect 20913 16065 20947 16099
rect 22385 16065 22419 16099
rect 23029 16065 23063 16099
rect 24593 16065 24627 16099
rect 1593 15997 1627 16031
rect 2789 15997 2823 16031
rect 3525 15997 3559 16031
rect 7021 15997 7055 16031
rect 10885 15997 10919 16031
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 14565 15997 14599 16031
rect 16037 15997 16071 16031
rect 18889 15997 18923 16031
rect 19993 15997 20027 16031
rect 21189 15997 21223 16031
rect 22477 15997 22511 16031
rect 22569 15997 22603 16031
rect 24041 15997 24075 16031
rect 10425 15929 10459 15963
rect 15485 15929 15519 15963
rect 25237 15929 25271 15963
rect 8125 15861 8159 15895
rect 8677 15861 8711 15895
rect 13461 15861 13495 15895
rect 16681 15861 16715 15895
rect 20545 15861 20579 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 1961 15657 1995 15691
rect 5825 15657 5859 15691
rect 6469 15657 6503 15691
rect 7113 15657 7147 15691
rect 23673 15657 23707 15691
rect 24225 15657 24259 15691
rect 16681 15589 16715 15623
rect 2881 15521 2915 15555
rect 4813 15521 4847 15555
rect 8401 15521 8435 15555
rect 10793 15521 10827 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 18705 15521 18739 15555
rect 19993 15521 20027 15555
rect 20177 15521 20211 15555
rect 21189 15521 21223 15555
rect 21373 15521 21407 15555
rect 2145 15453 2179 15487
rect 2605 15453 2639 15487
rect 4537 15453 4571 15487
rect 6009 15453 6043 15487
rect 6653 15453 6687 15487
rect 7297 15453 7331 15487
rect 7941 15453 7975 15487
rect 9965 15453 9999 15487
rect 10517 15453 10551 15487
rect 13093 15453 13127 15487
rect 21925 15453 21959 15487
rect 23029 15453 23063 15487
rect 24593 15453 24627 15487
rect 14565 15385 14599 15419
rect 21097 15385 21131 15419
rect 23949 15385 23983 15419
rect 3893 15317 3927 15351
rect 7757 15317 7791 15351
rect 9137 15317 9171 15351
rect 9781 15317 9815 15351
rect 12265 15317 12299 15351
rect 12725 15317 12759 15351
rect 13737 15317 13771 15351
rect 16037 15317 16071 15351
rect 16313 15317 16347 15351
rect 18981 15317 19015 15351
rect 19533 15317 19567 15351
rect 19901 15317 19935 15351
rect 20729 15317 20763 15351
rect 22569 15317 22603 15351
rect 25237 15317 25271 15351
rect 1777 15113 1811 15147
rect 1961 15113 1995 15147
rect 2605 15113 2639 15147
rect 3801 15113 3835 15147
rect 5825 15113 5859 15147
rect 9229 15113 9263 15147
rect 9873 15113 9907 15147
rect 13461 15113 13495 15147
rect 13737 15113 13771 15147
rect 16313 15113 16347 15147
rect 18981 15113 19015 15147
rect 5549 15045 5583 15079
rect 11989 15045 12023 15079
rect 15301 15045 15335 15079
rect 17141 15045 17175 15079
rect 21649 15045 21683 15079
rect 22109 15045 22143 15079
rect 25145 15045 25179 15079
rect 2789 14977 2823 15011
rect 3433 14977 3467 15011
rect 6009 14977 6043 15011
rect 6837 14977 6871 15011
rect 8493 14977 8527 15011
rect 8769 14977 8803 15011
rect 9413 14977 9447 15011
rect 10057 14977 10091 15011
rect 10517 14977 10551 15011
rect 11713 14977 11747 15011
rect 14197 14977 14231 15011
rect 15669 14977 15703 15011
rect 16865 14977 16899 15011
rect 22845 14977 22879 15011
rect 4077 14909 4111 14943
rect 4353 14909 4387 14943
rect 6561 14909 6595 14943
rect 7941 14909 7975 14943
rect 19349 14909 19383 14943
rect 19625 14909 19659 14943
rect 21097 14909 21131 14943
rect 23121 14909 23155 14943
rect 24593 14909 24627 14943
rect 3249 14841 3283 14875
rect 18613 14841 18647 14875
rect 7849 14773 7883 14807
rect 8585 14773 8619 14807
rect 11161 14773 11195 14807
rect 14841 14773 14875 14807
rect 15209 14773 15243 14807
rect 21373 14773 21407 14807
rect 22201 14773 22235 14807
rect 25237 14773 25271 14807
rect 2881 14569 2915 14603
rect 4169 14569 4203 14603
rect 4721 14569 4755 14603
rect 9321 14569 9355 14603
rect 13553 14569 13587 14603
rect 18245 14569 18279 14603
rect 18705 14569 18739 14603
rect 20545 14569 20579 14603
rect 22293 14569 22327 14603
rect 25237 14569 25271 14603
rect 3249 14501 3283 14535
rect 7849 14501 7883 14535
rect 10057 14501 10091 14535
rect 12449 14501 12483 14535
rect 13829 14501 13863 14535
rect 10977 14433 11011 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16497 14433 16531 14467
rect 16773 14433 16807 14467
rect 19901 14433 19935 14467
rect 19993 14433 20027 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 2329 14365 2363 14399
rect 2789 14365 2823 14399
rect 3433 14365 3467 14399
rect 4077 14365 4111 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 6009 14365 6043 14399
rect 6285 14365 6319 14399
rect 7481 14365 7515 14399
rect 8401 14365 8435 14399
rect 9505 14365 9539 14399
rect 10241 14365 10275 14399
rect 10701 14365 10735 14399
rect 12909 14365 12943 14399
rect 18889 14365 18923 14399
rect 20821 14365 20855 14399
rect 24593 14365 24627 14399
rect 22937 14297 22971 14331
rect 2145 14229 2179 14263
rect 5365 14229 5399 14263
rect 7297 14229 7331 14263
rect 7941 14229 7975 14263
rect 9045 14229 9079 14263
rect 16037 14229 16071 14263
rect 19441 14229 19475 14263
rect 19809 14229 19843 14263
rect 23305 14229 23339 14263
rect 23673 14229 23707 14263
rect 2145 14025 2179 14059
rect 2605 14025 2639 14059
rect 3249 14025 3283 14059
rect 4537 14025 4571 14059
rect 5181 14025 5215 14059
rect 5641 14025 5675 14059
rect 5917 14025 5951 14059
rect 7297 14025 7331 14059
rect 8769 14025 8803 14059
rect 9229 14025 9263 14059
rect 9413 14025 9447 14059
rect 10977 14025 11011 14059
rect 13277 14025 13311 14059
rect 15485 14025 15519 14059
rect 16681 14025 16715 14059
rect 17509 14025 17543 14059
rect 19533 14025 19567 14059
rect 20361 14025 20395 14059
rect 21189 14025 21223 14059
rect 10333 13957 10367 13991
rect 11713 13957 11747 13991
rect 18245 13957 18279 13991
rect 22109 13957 22143 13991
rect 24961 13957 24995 13991
rect 25145 13957 25179 13991
rect 1869 13889 1903 13923
rect 2329 13889 2363 13923
rect 2973 13889 3007 13923
rect 3433 13889 3467 13923
rect 4077 13889 4111 13923
rect 5365 13889 5399 13923
rect 6745 13889 6779 13923
rect 7481 13889 7515 13923
rect 7849 13889 7883 13923
rect 9045 13889 9079 13923
rect 9873 13889 9907 13923
rect 11161 13889 11195 13923
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 13737 13889 13771 13923
rect 16129 13889 16163 13923
rect 17417 13889 17451 13923
rect 20545 13889 20579 13923
rect 21097 13889 21131 13923
rect 22845 13889 22879 13923
rect 16313 13821 16347 13855
rect 17601 13821 17635 13855
rect 21373 13821 21407 13855
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 25329 13821 25363 13855
rect 3893 13753 3927 13787
rect 17049 13753 17083 13787
rect 22293 13753 22327 13787
rect 6561 13685 6595 13719
rect 9689 13685 9723 13719
rect 14000 13685 14034 13719
rect 20729 13685 20763 13719
rect 2605 13481 2639 13515
rect 3249 13481 3283 13515
rect 7113 13481 7147 13515
rect 13553 13481 13587 13515
rect 18245 13481 18279 13515
rect 21465 13481 21499 13515
rect 23673 13481 23707 13515
rect 1593 13413 1627 13447
rect 24041 13413 24075 13447
rect 24225 13413 24259 13447
rect 2145 13345 2179 13379
rect 11805 13345 11839 13379
rect 13829 13345 13863 13379
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 16773 13345 16807 13379
rect 18705 13345 18739 13379
rect 21925 13345 21959 13379
rect 25145 13345 25179 13379
rect 1777 13277 1811 13311
rect 2797 13277 2831 13311
rect 3433 13277 3467 13311
rect 4629 13277 4663 13311
rect 19717 13277 19751 13311
rect 2329 13209 2363 13243
rect 3985 13209 4019 13243
rect 9597 13209 9631 13243
rect 12081 13209 12115 13243
rect 14565 13209 14599 13243
rect 19993 13209 20027 13243
rect 22201 13209 22235 13243
rect 24961 13209 24995 13243
rect 6561 13141 6595 13175
rect 10885 13141 10919 13175
rect 16037 13141 16071 13175
rect 19349 13141 19383 13175
rect 24593 13141 24627 13175
rect 25053 13141 25087 13175
rect 1961 12937 1995 12971
rect 2605 12937 2639 12971
rect 10609 12937 10643 12971
rect 11529 12937 11563 12971
rect 12541 12937 12575 12971
rect 14289 12937 14323 12971
rect 15117 12937 15151 12971
rect 19533 12937 19567 12971
rect 24869 12937 24903 12971
rect 13001 12869 13035 12903
rect 16313 12869 16347 12903
rect 20729 12869 20763 12903
rect 1685 12801 1719 12835
rect 2145 12801 2179 12835
rect 2789 12801 2823 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 15301 12801 15335 12835
rect 15669 12801 15703 12835
rect 16865 12801 16899 12835
rect 19441 12801 19475 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 24225 12801 24259 12835
rect 25145 12801 25179 12835
rect 25329 12801 25363 12835
rect 3157 12733 3191 12767
rect 3249 12733 3283 12767
rect 17141 12733 17175 12767
rect 19625 12733 19659 12767
rect 20821 12733 20855 12767
rect 21557 12733 21591 12767
rect 22293 12733 22327 12767
rect 23765 12733 23799 12767
rect 18613 12665 18647 12699
rect 10977 12597 11011 12631
rect 19073 12597 19107 12631
rect 20269 12597 20303 12631
rect 21373 12597 21407 12631
rect 11529 12393 11563 12427
rect 11713 12393 11747 12427
rect 13737 12393 13771 12427
rect 25237 12393 25271 12427
rect 18613 12325 18647 12359
rect 15393 12257 15427 12291
rect 15761 12257 15795 12291
rect 19441 12257 19475 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 11989 12189 12023 12223
rect 13093 12189 13127 12223
rect 14289 12189 14323 12223
rect 17969 12189 18003 12223
rect 21649 12189 21683 12223
rect 24593 12189 24627 12223
rect 15301 12121 15335 12155
rect 16037 12121 16071 12155
rect 18889 12121 18923 12155
rect 19717 12121 19751 12155
rect 1961 12053 1995 12087
rect 12633 12053 12667 12087
rect 14933 12053 14967 12087
rect 17509 12053 17543 12087
rect 21189 12053 21223 12087
rect 24041 12053 24075 12087
rect 11897 11849 11931 11883
rect 12265 11849 12299 11883
rect 16497 11849 16531 11883
rect 16773 11849 16807 11883
rect 18889 11849 18923 11883
rect 13093 11781 13127 11815
rect 23305 11781 23339 11815
rect 25145 11781 25179 11815
rect 12817 11713 12851 11747
rect 19441 11713 19475 11747
rect 22201 11713 22235 11747
rect 23949 11713 23983 11747
rect 12541 11645 12575 11679
rect 14565 11645 14599 11679
rect 15025 11645 15059 11679
rect 15301 11645 15335 11679
rect 17141 11645 17175 11679
rect 17417 11645 17451 11679
rect 19717 11645 19751 11679
rect 16313 11577 16347 11611
rect 21189 11509 21223 11543
rect 21649 11509 21683 11543
rect 22293 11305 22327 11339
rect 25237 11305 25271 11339
rect 13185 11237 13219 11271
rect 14197 11237 14231 11271
rect 14473 11237 14507 11271
rect 15393 11237 15427 11271
rect 16313 11237 16347 11271
rect 16681 11237 16715 11271
rect 17969 11237 18003 11271
rect 20085 11237 20119 11271
rect 21189 11237 21223 11271
rect 23857 11169 23891 11203
rect 13737 11101 13771 11135
rect 14657 11101 14691 11135
rect 15669 11101 15703 11135
rect 16773 11101 16807 11135
rect 16957 11101 16991 11135
rect 17325 11101 17359 11135
rect 19441 11101 19475 11135
rect 20545 11101 20579 11135
rect 21741 11101 21775 11135
rect 22753 11101 22787 11135
rect 24593 11101 24627 11135
rect 15209 11033 15243 11067
rect 18337 11033 18371 11067
rect 18705 11033 18739 11067
rect 18889 11033 18923 11067
rect 21925 11033 21959 11067
rect 13553 10965 13587 10999
rect 14933 10965 14967 10999
rect 13645 10761 13679 10795
rect 13921 10761 13955 10795
rect 16129 10761 16163 10795
rect 16773 10761 16807 10795
rect 17969 10761 18003 10795
rect 19073 10761 19107 10795
rect 20361 10761 20395 10795
rect 23305 10693 23339 10727
rect 14381 10625 14415 10659
rect 15117 10625 15151 10659
rect 16313 10625 16347 10659
rect 17325 10625 17359 10659
rect 18429 10625 18463 10659
rect 19717 10625 19751 10659
rect 20821 10625 20855 10659
rect 21465 10625 21499 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 14841 10557 14875 10591
rect 24777 10557 24811 10591
rect 14197 10421 14231 10455
rect 17049 10421 17083 10455
rect 19441 10421 19475 10455
rect 14473 10217 14507 10251
rect 15117 10217 15151 10251
rect 15761 10217 15795 10251
rect 17049 10217 17083 10251
rect 17601 10217 17635 10251
rect 18705 10217 18739 10251
rect 20913 10217 20947 10251
rect 17969 10081 18003 10115
rect 19625 10081 19659 10115
rect 21373 10081 21407 10115
rect 25145 10081 25179 10115
rect 14657 10013 14691 10047
rect 15301 10013 15335 10047
rect 15945 10013 15979 10047
rect 16589 10013 16623 10047
rect 17233 10013 17267 10047
rect 18889 10013 18923 10047
rect 20269 10013 20303 10047
rect 23857 10013 23891 10047
rect 25053 10013 25087 10047
rect 19349 9945 19383 9979
rect 21649 9945 21683 9979
rect 24961 9945 24995 9979
rect 16405 9877 16439 9911
rect 23121 9877 23155 9911
rect 23949 9877 23983 9911
rect 24593 9877 24627 9911
rect 14749 9673 14783 9707
rect 15393 9673 15427 9707
rect 20177 9673 20211 9707
rect 15669 9605 15703 9639
rect 18153 9605 18187 9639
rect 23305 9605 23339 9639
rect 25145 9605 25179 9639
rect 15853 9537 15887 9571
rect 16313 9537 16347 9571
rect 17049 9537 17083 9571
rect 17693 9537 17727 9571
rect 18981 9537 19015 9571
rect 19625 9537 19659 9571
rect 20729 9537 20763 9571
rect 21373 9537 21407 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 19993 9469 20027 9503
rect 16129 9401 16163 9435
rect 18797 9401 18831 9435
rect 19441 9401 19475 9435
rect 20545 9401 20579 9435
rect 16865 9333 16899 9367
rect 17509 9333 17543 9367
rect 21189 9333 21223 9367
rect 11805 9129 11839 9163
rect 18061 9129 18095 9163
rect 19441 9129 19475 9163
rect 22109 9129 22143 9163
rect 25237 9129 25271 9163
rect 20085 9061 20119 9095
rect 10057 8993 10091 9027
rect 16129 8993 16163 9027
rect 16405 8993 16439 9027
rect 23857 8993 23891 9027
rect 17601 8925 17635 8959
rect 18245 8925 18279 8959
rect 18889 8925 18923 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20821 8925 20855 8959
rect 21465 8925 21499 8959
rect 22661 8925 22695 8959
rect 24593 8925 24627 8959
rect 10333 8857 10367 8891
rect 12173 8857 12207 8891
rect 17417 8789 17451 8823
rect 18705 8789 18739 8823
rect 19165 8585 19199 8619
rect 19809 8585 19843 8619
rect 20913 8585 20947 8619
rect 21281 8585 21315 8619
rect 17417 8449 17451 8483
rect 19349 8449 19383 8483
rect 19993 8449 20027 8483
rect 20637 8449 20671 8483
rect 22293 8449 22327 8483
rect 24041 8449 24075 8483
rect 17877 8381 17911 8415
rect 18153 8381 18187 8415
rect 23305 8381 23339 8415
rect 24777 8381 24811 8415
rect 17233 8313 17267 8347
rect 20453 8313 20487 8347
rect 19441 8041 19475 8075
rect 20545 8041 20579 8075
rect 20821 8041 20855 8075
rect 25237 8041 25271 8075
rect 17417 7905 17451 7939
rect 17693 7905 17727 7939
rect 18705 7905 18739 7939
rect 23857 7905 23891 7939
rect 19625 7837 19659 7871
rect 21281 7837 21315 7871
rect 22109 7837 22143 7871
rect 22661 7837 22695 7871
rect 24593 7837 24627 7871
rect 20085 7769 20119 7803
rect 21005 7701 21039 7735
rect 21925 7701 21959 7735
rect 17417 7497 17451 7531
rect 17969 7497 18003 7531
rect 18521 7497 18555 7531
rect 23305 7429 23339 7463
rect 25145 7429 25179 7463
rect 17601 7361 17635 7395
rect 18705 7361 18739 7395
rect 19165 7361 19199 7395
rect 19441 7361 19475 7395
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 20269 7293 20303 7327
rect 20637 7157 20671 7191
rect 21281 7157 21315 7191
rect 20729 6885 20763 6919
rect 24501 6817 24535 6851
rect 24685 6817 24719 6851
rect 19625 6749 19659 6783
rect 20269 6749 20303 6783
rect 20913 6749 20947 6783
rect 22661 6749 22695 6783
rect 23857 6749 23891 6783
rect 25145 6749 25179 6783
rect 21465 6681 21499 6715
rect 21649 6681 21683 6715
rect 22017 6681 22051 6715
rect 24869 6681 24903 6715
rect 25329 6681 25363 6715
rect 19441 6613 19475 6647
rect 20085 6613 20119 6647
rect 21189 6613 21223 6647
rect 22109 6613 22143 6647
rect 19717 6409 19751 6443
rect 20177 6409 20211 6443
rect 20913 6409 20947 6443
rect 21281 6409 21315 6443
rect 23305 6341 23339 6375
rect 20637 6273 20671 6307
rect 21465 6273 21499 6307
rect 22201 6273 22235 6307
rect 23949 6273 23983 6307
rect 24777 6205 24811 6239
rect 20453 6137 20487 6171
rect 25513 5865 25547 5899
rect 21097 5797 21131 5831
rect 25329 5797 25363 5831
rect 22017 5729 22051 5763
rect 20637 5661 20671 5695
rect 21281 5661 21315 5695
rect 22845 5661 22879 5695
rect 24869 5661 24903 5695
rect 23857 5593 23891 5627
rect 20453 5525 20487 5559
rect 24685 5525 24719 5559
rect 23305 5253 23339 5287
rect 21465 5185 21499 5219
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 24685 5117 24719 5151
rect 21281 4981 21315 5015
rect 22017 4777 22051 4811
rect 25513 4777 25547 4811
rect 25237 4709 25271 4743
rect 21741 4573 21775 4607
rect 22201 4573 22235 4607
rect 22845 4573 22879 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 24685 4437 24719 4471
rect 20269 4097 20303 4131
rect 22109 4097 22143 4131
rect 23949 4097 23983 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 25237 3689 25271 3723
rect 21005 3485 21039 3519
rect 22845 3485 22879 3519
rect 24869 3485 24903 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 24685 3349 24719 3383
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 23949 3009 23983 3043
rect 19441 2941 19475 2975
rect 21281 2941 21315 2975
rect 6837 2601 6871 2635
rect 21281 2465 21315 2499
rect 7021 2397 7055 2431
rect 7297 2397 7331 2431
rect 20269 2397 20303 2431
rect 22845 2397 22879 2431
rect 24777 2397 24811 2431
rect 23857 2329 23891 2363
rect 24593 2261 24627 2295
<< metal1 >>
rect 5626 26324 5632 26376
rect 5684 26364 5690 26376
rect 22370 26364 22376 26376
rect 5684 26336 22376 26364
rect 5684 26324 5690 26336
rect 22370 26324 22376 26336
rect 22428 26324 22434 26376
rect 3602 26256 3608 26308
rect 3660 26296 3666 26308
rect 19610 26296 19616 26308
rect 3660 26268 19616 26296
rect 3660 26256 3666 26268
rect 19610 26256 19616 26268
rect 19668 26256 19674 26308
rect 3694 26188 3700 26240
rect 3752 26228 3758 26240
rect 17954 26228 17960 26240
rect 3752 26200 17960 26228
rect 3752 26188 3758 26200
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 6270 26120 6276 26172
rect 6328 26160 6334 26172
rect 19794 26160 19800 26172
rect 6328 26132 19800 26160
rect 6328 26120 6334 26132
rect 19794 26120 19800 26132
rect 19852 26120 19858 26172
rect 3142 25644 3148 25696
rect 3200 25684 3206 25696
rect 10686 25684 10692 25696
rect 3200 25656 10692 25684
rect 3200 25644 3206 25656
rect 10686 25644 10692 25656
rect 10744 25644 10750 25696
rect 7374 25508 7380 25560
rect 7432 25548 7438 25560
rect 23750 25548 23756 25560
rect 7432 25520 23756 25548
rect 7432 25508 7438 25520
rect 23750 25508 23756 25520
rect 23808 25508 23814 25560
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 20806 25480 20812 25492
rect 4120 25452 20812 25480
rect 4120 25440 4126 25452
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 6546 25372 6552 25424
rect 6604 25412 6610 25424
rect 22554 25412 22560 25424
rect 6604 25384 22560 25412
rect 6604 25372 6610 25384
rect 22554 25372 22560 25384
rect 22612 25372 22618 25424
rect 3786 25304 3792 25356
rect 3844 25344 3850 25356
rect 23842 25344 23848 25356
rect 3844 25316 23848 25344
rect 3844 25304 3850 25316
rect 23842 25304 23848 25316
rect 23900 25304 23906 25356
rect 5258 25236 5264 25288
rect 5316 25276 5322 25288
rect 18598 25276 18604 25288
rect 5316 25248 18604 25276
rect 5316 25236 5322 25248
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 6178 25168 6184 25220
rect 6236 25208 6242 25220
rect 24394 25208 24400 25220
rect 6236 25180 24400 25208
rect 6236 25168 6242 25180
rect 24394 25168 24400 25180
rect 24452 25168 24458 25220
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 24210 25140 24216 25152
rect 7340 25112 24216 25140
rect 7340 25100 7346 25112
rect 24210 25100 24216 25112
rect 24268 25100 24274 25152
rect 14366 25032 14372 25084
rect 14424 25072 14430 25084
rect 20714 25072 20720 25084
rect 14424 25044 20720 25072
rect 14424 25032 14430 25044
rect 20714 25032 20720 25044
rect 20772 25032 20778 25084
rect 13538 24964 13544 25016
rect 13596 25004 13602 25016
rect 23474 25004 23480 25016
rect 13596 24976 23480 25004
rect 13596 24964 13602 24976
rect 23474 24964 23480 24976
rect 23532 24964 23538 25016
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 22278 24936 22284 24948
rect 7248 24908 22284 24936
rect 7248 24896 7254 24908
rect 22278 24896 22284 24908
rect 22336 24896 22342 24948
rect 9490 24828 9496 24880
rect 9548 24868 9554 24880
rect 22462 24868 22468 24880
rect 9548 24840 22468 24868
rect 9548 24828 9554 24840
rect 22462 24828 22468 24840
rect 22520 24828 22526 24880
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 19978 24800 19984 24812
rect 7800 24772 19984 24800
rect 7800 24760 7806 24772
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 3970 24624 3976 24676
rect 4028 24664 4034 24676
rect 11238 24664 11244 24676
rect 4028 24636 11244 24664
rect 4028 24624 4034 24636
rect 11238 24624 11244 24636
rect 11296 24624 11302 24676
rect 12158 24624 12164 24676
rect 12216 24664 12222 24676
rect 16390 24664 16396 24676
rect 12216 24636 16396 24664
rect 12216 24624 12222 24636
rect 16390 24624 16396 24636
rect 16448 24624 16454 24676
rect 4154 24556 4160 24608
rect 4212 24596 4218 24608
rect 14734 24596 14740 24608
rect 4212 24568 14740 24596
rect 4212 24556 4218 24568
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 22370 24556 22376 24608
rect 22428 24596 22434 24608
rect 24762 24596 24768 24608
rect 22428 24568 24768 24596
rect 22428 24556 22434 24568
rect 24762 24556 24768 24568
rect 24820 24556 24826 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 1765 24395 1823 24401
rect 1765 24361 1777 24395
rect 1811 24392 1823 24395
rect 3326 24392 3332 24404
rect 1811 24364 3332 24392
rect 1811 24361 1823 24364
rect 1765 24355 1823 24361
rect 3326 24352 3332 24364
rect 3384 24392 3390 24404
rect 4062 24392 4068 24404
rect 3384 24364 4068 24392
rect 3384 24352 3390 24364
rect 4062 24352 4068 24364
rect 4120 24352 4126 24404
rect 12618 24392 12624 24404
rect 6564 24364 12624 24392
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6454 24256 6460 24268
rect 3283 24228 6460 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6454 24216 6460 24228
rect 6512 24216 6518 24268
rect 6564 24265 6592 24364
rect 12618 24352 12624 24364
rect 12676 24352 12682 24404
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 15286 24392 15292 24404
rect 14516 24364 15292 24392
rect 14516 24352 14522 24364
rect 15286 24352 15292 24364
rect 15344 24392 15350 24404
rect 19610 24392 19616 24404
rect 15344 24364 19616 24392
rect 15344 24352 15350 24364
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 20714 24352 20720 24404
rect 20772 24392 20778 24404
rect 24397 24395 24455 24401
rect 24397 24392 24409 24395
rect 20772 24364 24409 24392
rect 20772 24352 20778 24364
rect 24397 24361 24409 24364
rect 24443 24392 24455 24395
rect 24443 24364 25084 24392
rect 24443 24361 24455 24364
rect 24397 24355 24455 24361
rect 11514 24324 11520 24336
rect 6656 24296 11520 24324
rect 6549 24259 6607 24265
rect 6549 24225 6561 24259
rect 6595 24225 6607 24259
rect 6549 24219 6607 24225
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2271 24160 3556 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 1581 24123 1639 24129
rect 1581 24089 1593 24123
rect 1627 24120 1639 24123
rect 2682 24120 2688 24132
rect 1627 24092 2688 24120
rect 1627 24089 1639 24092
rect 1581 24083 1639 24089
rect 2682 24080 2688 24092
rect 2740 24080 2746 24132
rect 3528 24120 3556 24160
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 3528 24092 4200 24120
rect 4172 24064 4200 24092
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 4062 24052 4068 24064
rect 4019 24024 4068 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 4154 24012 4160 24064
rect 4212 24012 4218 24064
rect 4816 24052 4844 24151
rect 4890 24148 4896 24200
rect 4948 24188 4954 24200
rect 6656 24188 6684 24296
rect 11514 24284 11520 24296
rect 11572 24284 11578 24336
rect 12342 24284 12348 24336
rect 12400 24324 12406 24336
rect 12400 24284 12434 24324
rect 12526 24284 12532 24336
rect 12584 24324 12590 24336
rect 18141 24327 18199 24333
rect 18141 24324 18153 24327
rect 12584 24296 18153 24324
rect 12584 24284 12590 24296
rect 18141 24293 18153 24296
rect 18187 24293 18199 24327
rect 22094 24324 22100 24336
rect 18141 24287 18199 24293
rect 18432 24296 22100 24324
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 12406 24256 12434 24284
rect 12805 24259 12863 24265
rect 12805 24256 12817 24259
rect 12406 24228 12817 24256
rect 12805 24225 12817 24228
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 13722 24216 13728 24268
rect 13780 24256 13786 24268
rect 18322 24256 18328 24268
rect 13780 24228 18328 24256
rect 13780 24216 13786 24228
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 4948 24160 6684 24188
rect 4948 24148 4954 24160
rect 7098 24148 7104 24200
rect 7156 24188 7162 24200
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 7156 24160 7205 24188
rect 7156 24148 7162 24160
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8662 24120 8668 24132
rect 5859 24092 8668 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 9033 24123 9091 24129
rect 9033 24089 9045 24123
rect 9079 24120 9091 24123
rect 9324 24120 9352 24151
rect 9858 24148 9864 24200
rect 9916 24148 9922 24200
rect 10962 24148 10968 24200
rect 11020 24148 11026 24200
rect 12345 24191 12403 24197
rect 12345 24188 12357 24191
rect 11440 24160 12357 24188
rect 9674 24120 9680 24132
rect 9079 24092 9680 24120
rect 9079 24089 9091 24092
rect 9033 24083 9091 24089
rect 9674 24080 9680 24092
rect 9732 24080 9738 24132
rect 11440 24120 11468 24160
rect 12345 24157 12357 24160
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 15194 24188 15200 24200
rect 14323 24160 15200 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 16758 24188 16764 24200
rect 15427 24160 16764 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 16850 24148 16856 24200
rect 16908 24148 16914 24200
rect 18432 24188 18460 24296
rect 22094 24284 22100 24296
rect 22152 24284 22158 24336
rect 18690 24216 18696 24268
rect 18748 24216 18754 24268
rect 18782 24216 18788 24268
rect 18840 24256 18846 24268
rect 22830 24256 22836 24268
rect 18840 24228 22836 24256
rect 18840 24216 18846 24228
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 23658 24216 23664 24268
rect 23716 24216 23722 24268
rect 25056 24265 25084 24364
rect 25041 24259 25099 24265
rect 25041 24225 25053 24259
rect 25087 24225 25099 24259
rect 25041 24219 25099 24225
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 17604 24160 18460 24188
rect 18601 24191 18659 24197
rect 17497 24123 17555 24129
rect 17497 24120 17509 24123
rect 10980 24092 11468 24120
rect 11532 24092 17509 24120
rect 10980 24064 11008 24092
rect 8386 24052 8392 24064
rect 4816 24024 8392 24052
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 10962 24012 10968 24064
rect 11020 24012 11026 24064
rect 11054 24012 11060 24064
rect 11112 24052 11118 24064
rect 11532 24052 11560 24092
rect 17497 24089 17509 24092
rect 17543 24089 17555 24123
rect 17497 24083 17555 24089
rect 11112 24024 11560 24052
rect 11701 24055 11759 24061
rect 11112 24012 11118 24024
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 13998 24052 14004 24064
rect 11747 24024 14004 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 14918 24012 14924 24064
rect 14976 24012 14982 24064
rect 15102 24012 15108 24064
rect 15160 24052 15166 24064
rect 16025 24055 16083 24061
rect 16025 24052 16037 24055
rect 15160 24024 16037 24052
rect 15160 24012 15166 24024
rect 16025 24021 16037 24024
rect 16071 24021 16083 24055
rect 16025 24015 16083 24021
rect 16298 24012 16304 24064
rect 16356 24012 16362 24064
rect 16482 24012 16488 24064
rect 16540 24052 16546 24064
rect 17604 24052 17632 24160
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 19518 24188 19524 24200
rect 18647 24160 19524 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19610 24148 19616 24200
rect 19668 24148 19674 24200
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 22186 24148 22192 24200
rect 22244 24148 22250 24200
rect 23676 24188 23704 24216
rect 23598 24160 23704 24188
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 18509 24123 18567 24129
rect 18509 24089 18521 24123
rect 18555 24120 18567 24123
rect 18555 24092 18828 24120
rect 18555 24089 18567 24092
rect 18509 24083 18567 24089
rect 18800 24064 18828 24092
rect 20898 24080 20904 24132
rect 20956 24120 20962 24132
rect 20993 24123 21051 24129
rect 20993 24120 21005 24123
rect 20956 24092 21005 24120
rect 20956 24080 20962 24092
rect 20993 24089 21005 24092
rect 21039 24089 21051 24123
rect 20993 24083 21051 24089
rect 21913 24123 21971 24129
rect 21913 24089 21925 24123
rect 21959 24120 21971 24123
rect 22370 24120 22376 24132
rect 21959 24092 22376 24120
rect 21959 24089 21971 24092
rect 21913 24083 21971 24089
rect 22370 24080 22376 24092
rect 22428 24080 22434 24132
rect 22465 24123 22523 24129
rect 22465 24089 22477 24123
rect 22511 24089 22523 24123
rect 25148 24120 25176 24219
rect 22465 24083 22523 24089
rect 24136 24092 25176 24120
rect 16540 24024 17632 24052
rect 16540 24012 16546 24024
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 17773 24055 17831 24061
rect 17773 24052 17785 24055
rect 17736 24024 17785 24052
rect 17736 24012 17742 24024
rect 17773 24021 17785 24024
rect 17819 24021 17831 24055
rect 17773 24015 17831 24021
rect 18782 24012 18788 24064
rect 18840 24012 18846 24064
rect 19150 24012 19156 24064
rect 19208 24052 19214 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 19208 24024 19441 24052
rect 19208 24012 19214 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 22094 24012 22100 24064
rect 22152 24052 22158 24064
rect 22480 24052 22508 24083
rect 24136 24064 24164 24092
rect 22152 24024 22508 24052
rect 23937 24055 23995 24061
rect 22152 24012 22158 24024
rect 23937 24021 23949 24055
rect 23983 24052 23995 24055
rect 24118 24052 24124 24064
rect 23983 24024 24124 24052
rect 23983 24021 23995 24024
rect 23937 24015 23995 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 24854 24052 24860 24064
rect 24627 24024 24860 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25498 24052 25504 24064
rect 25004 24024 25504 24052
rect 25004 24012 25010 24024
rect 25498 24012 25504 24024
rect 25556 24012 25562 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 6546 23808 6552 23860
rect 6604 23808 6610 23860
rect 6840 23820 11192 23848
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5350 23780 5356 23792
rect 4019 23752 5356 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 2958 23672 2964 23724
rect 3016 23672 3022 23724
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 4890 23712 4896 23724
rect 4847 23684 4896 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 6840 23721 6868 23820
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 10134 23780 10140 23792
rect 9171 23752 10140 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 11164 23780 11192 23820
rect 11330 23808 11336 23860
rect 11388 23848 11394 23860
rect 11388 23820 13860 23848
rect 11388 23808 11394 23820
rect 13630 23780 13636 23792
rect 11164 23752 13636 23780
rect 13630 23740 13636 23752
rect 13688 23740 13694 23792
rect 13832 23780 13860 23820
rect 14090 23808 14096 23860
rect 14148 23808 14154 23860
rect 14553 23851 14611 23857
rect 14553 23817 14565 23851
rect 14599 23848 14611 23851
rect 14599 23820 17540 23848
rect 14599 23817 14611 23820
rect 14553 23811 14611 23817
rect 13832 23752 14596 23780
rect 6813 23715 6871 23721
rect 6813 23681 6825 23715
rect 6859 23681 6871 23715
rect 6813 23675 6871 23681
rect 7469 23715 7527 23721
rect 7469 23681 7481 23715
rect 7515 23712 7527 23715
rect 7515 23684 7880 23712
rect 7515 23681 7527 23684
rect 7469 23675 7527 23681
rect 1765 23647 1823 23653
rect 1765 23613 1777 23647
rect 1811 23644 1823 23647
rect 1946 23644 1952 23656
rect 1811 23616 1952 23644
rect 1811 23613 1823 23616
rect 1765 23607 1823 23613
rect 1946 23604 1952 23616
rect 2004 23604 2010 23656
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 7558 23644 7564 23656
rect 5859 23616 7564 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7852 23644 7880 23684
rect 7926 23672 7932 23724
rect 7984 23672 7990 23724
rect 9766 23672 9772 23724
rect 9824 23672 9830 23724
rect 10042 23672 10048 23724
rect 10100 23712 10106 23724
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 10100 23684 12081 23712
rect 10100 23672 10106 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 13814 23672 13820 23724
rect 13872 23712 13878 23724
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 13872 23684 14473 23712
rect 13872 23672 13878 23684
rect 14461 23681 14473 23684
rect 14507 23681 14519 23715
rect 14568 23712 14596 23752
rect 15010 23740 15016 23792
rect 15068 23780 15074 23792
rect 16209 23783 16267 23789
rect 16209 23780 16221 23783
rect 15068 23752 16221 23780
rect 15068 23740 15074 23752
rect 16209 23749 16221 23752
rect 16255 23749 16267 23783
rect 17512 23780 17540 23820
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 20349 23851 20407 23857
rect 20349 23848 20361 23851
rect 17644 23820 20361 23848
rect 17644 23808 17650 23820
rect 20349 23817 20361 23820
rect 20395 23817 20407 23851
rect 20349 23811 20407 23817
rect 20717 23851 20775 23857
rect 20717 23817 20729 23851
rect 20763 23848 20775 23851
rect 20806 23848 20812 23860
rect 20763 23820 20812 23848
rect 20763 23817 20775 23820
rect 20717 23811 20775 23817
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 22278 23848 22284 23860
rect 22235 23820 22284 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 22278 23808 22284 23820
rect 22336 23848 22342 23860
rect 22336 23820 22600 23848
rect 22336 23808 22342 23820
rect 18414 23780 18420 23792
rect 17512 23752 18420 23780
rect 16209 23743 16267 23749
rect 18414 23740 18420 23752
rect 18472 23740 18478 23792
rect 20898 23780 20904 23792
rect 19550 23752 20904 23780
rect 20898 23740 20904 23752
rect 20956 23780 20962 23792
rect 21545 23783 21603 23789
rect 21545 23780 21557 23783
rect 20956 23752 21557 23780
rect 20956 23740 20962 23752
rect 21545 23749 21557 23752
rect 21591 23780 21603 23783
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 21591 23752 21833 23780
rect 21591 23749 21603 23752
rect 21545 23743 21603 23749
rect 21821 23749 21833 23752
rect 21867 23780 21879 23783
rect 22002 23780 22008 23792
rect 21867 23752 22008 23780
rect 21867 23749 21879 23752
rect 21821 23743 21879 23749
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 22572 23789 22600 23820
rect 22830 23808 22836 23860
rect 22888 23848 22894 23860
rect 24397 23851 24455 23857
rect 24397 23848 24409 23851
rect 22888 23820 24409 23848
rect 22888 23808 22894 23820
rect 24397 23817 24409 23820
rect 24443 23848 24455 23851
rect 25041 23851 25099 23857
rect 25041 23848 25053 23851
rect 24443 23820 25053 23848
rect 24443 23817 24455 23820
rect 24397 23811 24455 23817
rect 25041 23817 25053 23820
rect 25087 23817 25099 23851
rect 25041 23811 25099 23817
rect 22557 23783 22615 23789
rect 22557 23749 22569 23783
rect 22603 23749 22615 23783
rect 22557 23743 22615 23749
rect 24762 23740 24768 23792
rect 24820 23780 24826 23792
rect 24949 23783 25007 23789
rect 24949 23780 24961 23783
rect 24820 23752 24961 23780
rect 24820 23740 24826 23752
rect 24949 23749 24961 23752
rect 24995 23749 25007 23783
rect 24949 23743 25007 23749
rect 15286 23712 15292 23724
rect 14568 23684 15292 23712
rect 14461 23675 14519 23681
rect 15286 23672 15292 23684
rect 15344 23672 15350 23724
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23712 15623 23715
rect 16022 23712 16028 23724
rect 15611 23684 16028 23712
rect 15611 23681 15623 23684
rect 15565 23675 15623 23681
rect 16022 23672 16028 23684
rect 16080 23672 16086 23724
rect 16482 23712 16488 23724
rect 16132 23684 16488 23712
rect 11330 23644 11336 23656
rect 7852 23616 11336 23644
rect 11330 23604 11336 23616
rect 11388 23604 11394 23656
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 14737 23647 14795 23653
rect 14737 23613 14749 23647
rect 14783 23644 14795 23647
rect 15194 23644 15200 23656
rect 14783 23616 15200 23644
rect 14783 23613 14795 23616
rect 14737 23607 14795 23613
rect 15194 23604 15200 23616
rect 15252 23644 15258 23656
rect 15378 23644 15384 23656
rect 15252 23616 15384 23644
rect 15252 23604 15258 23616
rect 15378 23604 15384 23616
rect 15436 23604 15442 23656
rect 15470 23604 15476 23656
rect 15528 23644 15534 23656
rect 16132 23644 16160 23684
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 16945 23715 17003 23721
rect 16945 23681 16957 23715
rect 16991 23712 17003 23715
rect 17402 23712 17408 23724
rect 16991 23684 17408 23712
rect 16991 23681 17003 23684
rect 16945 23675 17003 23681
rect 17402 23672 17408 23684
rect 17460 23672 17466 23724
rect 23658 23672 23664 23724
rect 23716 23672 23722 23724
rect 15528 23616 16160 23644
rect 15528 23604 15534 23616
rect 17954 23604 17960 23656
rect 18012 23644 18018 23656
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 18012 23616 18061 23644
rect 18012 23604 18018 23616
rect 18049 23613 18061 23616
rect 18095 23613 18107 23647
rect 18325 23647 18383 23653
rect 18325 23644 18337 23647
rect 18049 23607 18107 23613
rect 18156 23616 18337 23644
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 18156 23576 18184 23616
rect 18325 23613 18337 23616
rect 18371 23613 18383 23647
rect 18325 23607 18383 23613
rect 20806 23604 20812 23656
rect 20864 23604 20870 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23613 20959 23647
rect 20901 23607 20959 23613
rect 20916 23576 20944 23607
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 2363 23548 18184 23576
rect 19812 23548 20944 23576
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 5166 23468 5172 23520
rect 5224 23508 5230 23520
rect 7926 23508 7932 23520
rect 5224 23480 7932 23508
rect 5224 23468 5230 23480
rect 7926 23468 7932 23480
rect 7984 23468 7990 23520
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 10962 23508 10968 23520
rect 10468 23480 10968 23508
rect 10468 23468 10474 23480
rect 10962 23468 10968 23480
rect 11020 23508 11026 23520
rect 11517 23511 11575 23517
rect 11517 23508 11529 23511
rect 11020 23480 11529 23508
rect 11020 23468 11026 23480
rect 11517 23477 11529 23480
rect 11563 23477 11575 23511
rect 11517 23471 11575 23477
rect 11793 23511 11851 23517
rect 11793 23477 11805 23511
rect 11839 23508 11851 23511
rect 12250 23508 12256 23520
rect 11839 23480 12256 23508
rect 11839 23477 11851 23480
rect 11793 23471 11851 23477
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 13814 23468 13820 23520
rect 13872 23468 13878 23520
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 15197 23511 15255 23517
rect 15197 23508 15209 23511
rect 14700 23480 15209 23508
rect 14700 23468 14706 23480
rect 15197 23477 15209 23480
rect 15243 23508 15255 23511
rect 15746 23508 15752 23520
rect 15243 23480 15752 23508
rect 15243 23477 15255 23480
rect 15197 23471 15255 23477
rect 15746 23468 15752 23480
rect 15804 23508 15810 23520
rect 17034 23508 17040 23520
rect 15804 23480 17040 23508
rect 15804 23468 15810 23480
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 17218 23468 17224 23520
rect 17276 23508 17282 23520
rect 17589 23511 17647 23517
rect 17589 23508 17601 23511
rect 17276 23480 17601 23508
rect 17276 23468 17282 23480
rect 17589 23477 17601 23480
rect 17635 23477 17647 23511
rect 17589 23471 17647 23477
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 19812 23517 19840 23548
rect 24946 23536 24952 23588
rect 25004 23576 25010 23588
rect 25148 23576 25176 23607
rect 25004 23548 25176 23576
rect 25004 23536 25010 23548
rect 19797 23511 19855 23517
rect 19797 23508 19809 23511
rect 19484 23480 19809 23508
rect 19484 23468 19490 23480
rect 19797 23477 19809 23480
rect 19843 23477 19855 23511
rect 19797 23471 19855 23477
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 21361 23511 21419 23517
rect 21361 23508 21373 23511
rect 20772 23480 21373 23508
rect 20772 23468 20778 23480
rect 21361 23477 21373 23480
rect 21407 23477 21419 23511
rect 21361 23471 21419 23477
rect 24026 23468 24032 23520
rect 24084 23468 24090 23520
rect 24581 23511 24639 23517
rect 24581 23477 24593 23511
rect 24627 23508 24639 23511
rect 25130 23508 25136 23520
rect 24627 23480 25136 23508
rect 24627 23477 24639 23480
rect 24581 23471 24639 23477
rect 25130 23468 25136 23480
rect 25188 23468 25194 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 3878 23264 3884 23316
rect 3936 23304 3942 23316
rect 4890 23304 4896 23316
rect 3936 23276 4896 23304
rect 3936 23264 3942 23276
rect 4890 23264 4896 23276
rect 4948 23264 4954 23316
rect 8386 23264 8392 23316
rect 8444 23304 8450 23316
rect 9309 23307 9367 23313
rect 9309 23304 9321 23307
rect 8444 23276 9321 23304
rect 8444 23264 8450 23276
rect 9309 23273 9321 23276
rect 9355 23273 9367 23307
rect 9309 23267 9367 23273
rect 11606 23264 11612 23316
rect 11664 23304 11670 23316
rect 11664 23276 12296 23304
rect 11664 23264 11670 23276
rect 11146 23236 11152 23248
rect 5276 23208 11152 23236
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 4614 23168 4620 23180
rect 3283 23140 4620 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 2222 23060 2228 23112
rect 2280 23060 2286 23112
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 5276 23100 5304 23208
rect 11146 23196 11152 23208
rect 11204 23196 11210 23248
rect 12268 23236 12296 23276
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 14461 23307 14519 23313
rect 14461 23304 14473 23307
rect 12492 23276 14473 23304
rect 12492 23264 12498 23276
rect 14461 23273 14473 23276
rect 14507 23273 14519 23307
rect 14461 23267 14519 23273
rect 15120 23276 16344 23304
rect 12618 23236 12624 23248
rect 12268 23208 12624 23236
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 13630 23196 13636 23248
rect 13688 23236 13694 23248
rect 15120 23236 15148 23276
rect 13688 23208 15148 23236
rect 13688 23196 13694 23208
rect 6549 23171 6607 23177
rect 6549 23137 6561 23171
rect 6595 23168 6607 23171
rect 7650 23168 7656 23180
rect 6595 23140 7656 23168
rect 6595 23137 6607 23140
rect 6549 23131 6607 23137
rect 7650 23128 7656 23140
rect 7708 23128 7714 23180
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23168 8263 23171
rect 9398 23168 9404 23180
rect 8251 23140 9404 23168
rect 8251 23137 8263 23140
rect 8205 23131 8263 23137
rect 9398 23128 9404 23140
rect 9456 23128 9462 23180
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 13906 23168 13912 23180
rect 13740 23140 13912 23168
rect 4295 23072 5304 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 5442 23060 5448 23112
rect 5500 23060 5506 23112
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 1578 22992 1584 23044
rect 1636 22992 1642 23044
rect 4982 22992 4988 23044
rect 5040 23032 5046 23044
rect 7208 23032 7236 23063
rect 9950 23060 9956 23112
rect 10008 23060 10014 23112
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 10192 23072 11713 23100
rect 10192 23060 10198 23072
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 11701 23063 11759 23069
rect 12250 23060 12256 23112
rect 12308 23100 12314 23112
rect 13740 23109 13768 23140
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15286 23128 15292 23180
rect 15344 23128 15350 23180
rect 16316 23168 16344 23276
rect 17034 23264 17040 23316
rect 17092 23304 17098 23316
rect 17678 23304 17684 23316
rect 17092 23276 17684 23304
rect 17092 23264 17098 23276
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 17770 23264 17776 23316
rect 17828 23264 17834 23316
rect 18322 23264 18328 23316
rect 18380 23264 18386 23316
rect 18598 23264 18604 23316
rect 18656 23264 18662 23316
rect 21542 23304 21548 23316
rect 19536 23276 21548 23304
rect 16482 23196 16488 23248
rect 16540 23236 16546 23248
rect 17494 23236 17500 23248
rect 16540 23208 17500 23236
rect 16540 23196 16546 23208
rect 17494 23196 17500 23208
rect 17552 23196 17558 23248
rect 17788 23236 17816 23264
rect 19536 23236 19564 23276
rect 21542 23264 21548 23276
rect 21600 23264 21606 23316
rect 22002 23264 22008 23316
rect 22060 23304 22066 23316
rect 23658 23304 23664 23316
rect 22060 23276 23664 23304
rect 22060 23264 22066 23276
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 21177 23239 21235 23245
rect 21177 23236 21189 23239
rect 17788 23208 19564 23236
rect 20732 23208 21189 23236
rect 17770 23168 17776 23180
rect 16316 23140 17776 23168
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 17920 23140 19717 23168
rect 17920 23128 17926 23140
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 19794 23128 19800 23180
rect 19852 23168 19858 23180
rect 20732 23168 20760 23208
rect 21177 23205 21189 23208
rect 21223 23205 21235 23239
rect 21177 23199 21235 23205
rect 19852 23140 20760 23168
rect 19852 23128 19858 23140
rect 20898 23128 20904 23180
rect 20956 23128 20962 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 22278 23168 22284 23180
rect 21683 23140 22284 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22278 23128 22284 23140
rect 22336 23168 22342 23180
rect 23290 23168 23296 23180
rect 22336 23140 23296 23168
rect 22336 23128 22342 23140
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23658 23128 23664 23180
rect 23716 23128 23722 23180
rect 24026 23128 24032 23180
rect 24084 23168 24090 23180
rect 25133 23171 25191 23177
rect 25133 23168 25145 23171
rect 24084 23140 25145 23168
rect 24084 23128 24090 23140
rect 25133 23137 25145 23140
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 13725 23103 13783 23109
rect 13725 23100 13737 23103
rect 12308 23072 13737 23100
rect 12308 23060 12314 23072
rect 13725 23069 13737 23072
rect 13771 23069 13783 23103
rect 13725 23063 13783 23069
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14274 23100 14280 23112
rect 13872 23072 14280 23100
rect 13872 23060 13878 23072
rect 14274 23060 14280 23072
rect 14332 23100 14338 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14332 23072 15025 23100
rect 14332 23060 14338 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 17126 23060 17132 23112
rect 17184 23100 17190 23112
rect 17494 23100 17500 23112
rect 17184 23072 17500 23100
rect 17184 23060 17190 23072
rect 17494 23060 17500 23072
rect 17552 23060 17558 23112
rect 17586 23060 17592 23112
rect 17644 23060 17650 23112
rect 17954 23060 17960 23112
rect 18012 23100 18018 23112
rect 19334 23100 19340 23112
rect 18012 23072 19340 23100
rect 18012 23060 18018 23072
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 20916 23100 20944 23128
rect 20838 23072 20944 23100
rect 19429 23063 19487 23069
rect 5040 23004 7236 23032
rect 9217 23035 9275 23041
rect 5040 22992 5046 23004
rect 9217 23001 9229 23035
rect 9263 23032 9275 23035
rect 9858 23032 9864 23044
rect 9263 23004 9864 23032
rect 9263 23001 9275 23004
rect 9217 22995 9275 23001
rect 9858 22992 9864 23004
rect 9916 22992 9922 23044
rect 11974 23032 11980 23044
rect 10244 23004 11980 23032
rect 1762 22924 1768 22976
rect 1820 22924 1826 22976
rect 2682 22924 2688 22976
rect 2740 22964 2746 22976
rect 3881 22967 3939 22973
rect 3881 22964 3893 22967
rect 2740 22936 3893 22964
rect 2740 22924 2746 22936
rect 3881 22933 3893 22936
rect 3927 22933 3939 22967
rect 3881 22927 3939 22933
rect 4893 22967 4951 22973
rect 4893 22933 4905 22967
rect 4939 22964 4951 22967
rect 7834 22964 7840 22976
rect 4939 22936 7840 22964
rect 4939 22933 4951 22936
rect 4893 22927 4951 22933
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 8938 22924 8944 22976
rect 8996 22964 9002 22976
rect 10244 22964 10272 23004
rect 11974 22992 11980 23004
rect 12032 22992 12038 23044
rect 12618 22992 12624 23044
rect 12676 22992 12682 23044
rect 14369 23035 14427 23041
rect 14369 23001 14381 23035
rect 14415 23032 14427 23035
rect 14826 23032 14832 23044
rect 14415 23004 14832 23032
rect 14415 23001 14427 23004
rect 14369 22995 14427 23001
rect 14826 22992 14832 23004
rect 14884 22992 14890 23044
rect 15746 22992 15752 23044
rect 15804 22992 15810 23044
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 17681 23035 17739 23041
rect 17681 23032 17693 23035
rect 17368 23004 17693 23032
rect 17368 22992 17374 23004
rect 17681 23001 17693 23004
rect 17727 23001 17739 23035
rect 17681 22995 17739 23001
rect 18322 22992 18328 23044
rect 18380 23032 18386 23044
rect 18509 23035 18567 23041
rect 18509 23032 18521 23035
rect 18380 23004 18521 23032
rect 18380 22992 18386 23004
rect 18509 23001 18521 23004
rect 18555 23001 18567 23035
rect 18690 23032 18696 23044
rect 18509 22995 18567 23001
rect 18616 23004 18696 23032
rect 8996 22936 10272 22964
rect 8996 22924 9002 22936
rect 10318 22924 10324 22976
rect 10376 22964 10382 22976
rect 12342 22964 12348 22976
rect 10376 22936 12348 22964
rect 10376 22924 10382 22936
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 13541 22967 13599 22973
rect 13541 22933 13553 22967
rect 13587 22964 13599 22967
rect 16666 22964 16672 22976
rect 13587 22936 16672 22964
rect 13587 22933 13599 22936
rect 13541 22927 13599 22933
rect 16666 22924 16672 22936
rect 16724 22924 16730 22976
rect 16758 22924 16764 22976
rect 16816 22924 16822 22976
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 17221 22967 17279 22973
rect 17221 22964 17233 22967
rect 17092 22936 17233 22964
rect 17092 22924 17098 22936
rect 17221 22933 17233 22936
rect 17267 22933 17279 22967
rect 17221 22927 17279 22933
rect 17586 22924 17592 22976
rect 17644 22964 17650 22976
rect 18616 22964 18644 23004
rect 18690 22992 18696 23004
rect 18748 23032 18754 23044
rect 19794 23032 19800 23044
rect 18748 23004 19800 23032
rect 18748 22992 18754 23004
rect 19794 22992 19800 23004
rect 19852 22992 19858 23044
rect 21913 23035 21971 23041
rect 21913 23032 21925 23035
rect 21008 23004 21925 23032
rect 17644 22936 18644 22964
rect 17644 22924 17650 22936
rect 18966 22924 18972 22976
rect 19024 22924 19030 22976
rect 19426 22924 19432 22976
rect 19484 22964 19490 22976
rect 21008 22964 21036 23004
rect 21913 23001 21925 23004
rect 21959 23001 21971 23035
rect 23676 23032 23704 23128
rect 24762 23032 24768 23044
rect 23138 23004 24768 23032
rect 21913 22995 21971 23001
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 24949 23035 25007 23041
rect 24949 23001 24961 23035
rect 24995 23032 25007 23035
rect 26786 23032 26792 23044
rect 24995 23004 26792 23032
rect 24995 23001 25007 23004
rect 24949 22995 25007 23001
rect 26786 22992 26792 23004
rect 26844 22992 26850 23044
rect 19484 22936 21036 22964
rect 19484 22924 19490 22936
rect 22738 22924 22744 22976
rect 22796 22964 22802 22976
rect 23385 22967 23443 22973
rect 23385 22964 23397 22967
rect 22796 22936 23397 22964
rect 22796 22924 22802 22936
rect 23385 22933 23397 22936
rect 23431 22933 23443 22967
rect 23385 22927 23443 22933
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 23845 22967 23903 22973
rect 23845 22964 23857 22967
rect 23624 22936 23857 22964
rect 23624 22924 23630 22936
rect 23845 22933 23857 22936
rect 23891 22933 23903 22967
rect 23845 22927 23903 22933
rect 23934 22924 23940 22976
rect 23992 22964 23998 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23992 22936 24593 22964
rect 23992 22924 23998 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 25038 22924 25044 22976
rect 25096 22924 25102 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 2222 22720 2228 22772
rect 2280 22760 2286 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 2280 22732 13093 22760
rect 2280 22720 2286 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13556 22732 15240 22760
rect 1762 22692 1768 22704
rect 1688 22664 1768 22692
rect 1688 22633 1716 22664
rect 1762 22652 1768 22664
rect 1820 22692 1826 22704
rect 3694 22692 3700 22704
rect 1820 22664 3700 22692
rect 1820 22652 1826 22664
rect 3694 22652 3700 22664
rect 3752 22652 3758 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 5350 22692 5356 22704
rect 4356 22664 5356 22692
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 4356 22624 4384 22664
rect 5350 22652 5356 22664
rect 5408 22652 5414 22704
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 5902 22652 5908 22704
rect 5960 22692 5966 22704
rect 5960 22664 7604 22692
rect 5960 22652 5966 22664
rect 3007 22596 4384 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 6638 22584 6644 22636
rect 6696 22584 6702 22636
rect 6914 22584 6920 22636
rect 6972 22624 6978 22636
rect 7282 22624 7288 22636
rect 6972 22596 7288 22624
rect 6972 22584 6978 22596
rect 7282 22584 7288 22596
rect 7340 22584 7346 22636
rect 7576 22633 7604 22664
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 11146 22652 11152 22704
rect 11204 22692 11210 22704
rect 13556 22692 13584 22732
rect 13814 22692 13820 22704
rect 11204 22664 13584 22692
rect 13648 22664 13820 22692
rect 11204 22652 11210 22664
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 10778 22584 10784 22636
rect 10836 22584 10842 22636
rect 11882 22624 11888 22636
rect 10888 22596 11888 22624
rect 2317 22559 2375 22565
rect 2317 22525 2329 22559
rect 2363 22556 2375 22559
rect 6730 22556 6736 22568
rect 2363 22528 6736 22556
rect 2363 22525 2375 22528
rect 2317 22519 2375 22525
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9677 22559 9735 22565
rect 9677 22556 9689 22559
rect 9401 22519 9459 22525
rect 9508 22528 9689 22556
rect 2746 22460 7696 22488
rect 1302 22380 1308 22432
rect 1360 22420 1366 22432
rect 2746 22420 2774 22460
rect 1360 22392 2774 22420
rect 1360 22380 1366 22392
rect 6730 22380 6736 22432
rect 6788 22380 6794 22432
rect 7668 22420 7696 22460
rect 7742 22448 7748 22500
rect 7800 22488 7806 22500
rect 9508 22488 9536 22528
rect 9677 22525 9689 22528
rect 9723 22525 9735 22559
rect 9677 22519 9735 22525
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 10888 22556 10916 22596
rect 11882 22584 11888 22596
rect 11940 22584 11946 22636
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12342 22624 12348 22636
rect 12207 22596 12348 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 9824 22528 10916 22556
rect 9824 22516 9830 22528
rect 11146 22516 11152 22568
rect 11204 22516 11210 22568
rect 11517 22491 11575 22497
rect 11517 22488 11529 22491
rect 7800 22460 9536 22488
rect 10704 22460 11529 22488
rect 7800 22448 7806 22460
rect 10704 22420 10732 22460
rect 11517 22457 11529 22460
rect 11563 22488 11575 22491
rect 12084 22488 12112 22587
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 13648 22633 13676 22664
rect 13814 22652 13820 22664
rect 13872 22652 13878 22704
rect 14550 22652 14556 22704
rect 14608 22652 14614 22704
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12492 22596 13001 22624
rect 12492 22584 12498 22596
rect 12989 22593 13001 22596
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22593 13691 22627
rect 15212 22624 15240 22732
rect 15378 22720 15384 22772
rect 15436 22720 15442 22772
rect 17862 22760 17868 22772
rect 16868 22732 17868 22760
rect 15930 22652 15936 22704
rect 15988 22692 15994 22704
rect 16298 22692 16304 22704
rect 15988 22664 16304 22692
rect 15988 22652 15994 22664
rect 16298 22652 16304 22664
rect 16356 22652 16362 22704
rect 16114 22624 16120 22636
rect 15212 22596 16120 22624
rect 13633 22587 13691 22593
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16868 22633 16896 22732
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18966 22760 18972 22772
rect 18012 22732 18972 22760
rect 18012 22720 18018 22732
rect 18966 22720 18972 22732
rect 19024 22720 19030 22772
rect 19518 22720 19524 22772
rect 19576 22760 19582 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 19576 22732 20269 22760
rect 19576 22720 19582 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 20257 22723 20315 22729
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20956 22732 21465 22760
rect 20956 22720 20962 22732
rect 21453 22729 21465 22732
rect 21499 22729 21511 22763
rect 21453 22723 21511 22729
rect 21542 22720 21548 22772
rect 21600 22760 21606 22772
rect 24302 22760 24308 22772
rect 21600 22732 24308 22760
rect 21600 22720 21606 22732
rect 24302 22720 24308 22732
rect 24360 22720 24366 22772
rect 17126 22652 17132 22704
rect 17184 22652 17190 22704
rect 17678 22652 17684 22704
rect 17736 22652 17742 22704
rect 19429 22695 19487 22701
rect 19429 22661 19441 22695
rect 19475 22692 19487 22695
rect 19886 22692 19892 22704
rect 19475 22664 19892 22692
rect 19475 22661 19487 22664
rect 19429 22655 19487 22661
rect 19886 22652 19892 22664
rect 19944 22652 19950 22704
rect 22278 22652 22284 22704
rect 22336 22692 22342 22704
rect 22373 22695 22431 22701
rect 22373 22692 22385 22695
rect 22336 22664 22385 22692
rect 22336 22652 22342 22664
rect 22373 22661 22385 22664
rect 22419 22661 22431 22695
rect 22373 22655 22431 22661
rect 23474 22652 23480 22704
rect 23532 22692 23538 22704
rect 23569 22695 23627 22701
rect 23569 22692 23581 22695
rect 23532 22664 23581 22692
rect 23532 22652 23538 22664
rect 23569 22661 23581 22664
rect 23615 22661 23627 22695
rect 23569 22655 23627 22661
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22624 19579 22627
rect 19702 22624 19708 22636
rect 19567 22596 19708 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 20625 22627 20683 22633
rect 20625 22593 20637 22627
rect 20671 22593 20683 22627
rect 24702 22596 24808 22624
rect 20625 22587 20683 22593
rect 12250 22516 12256 22568
rect 12308 22516 12314 22568
rect 13909 22559 13967 22565
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 13955 22528 14964 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 11563 22460 12112 22488
rect 14936 22488 14964 22528
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 16816 22528 19625 22556
rect 16816 22516 16822 22528
rect 19613 22525 19625 22528
rect 19659 22525 19671 22559
rect 20640 22556 20668 22587
rect 24780 22568 24808 22596
rect 19613 22519 19671 22525
rect 19720 22528 20668 22556
rect 15102 22488 15108 22500
rect 14936 22460 15108 22488
rect 11563 22457 11575 22460
rect 11517 22451 11575 22457
rect 15102 22448 15108 22460
rect 15160 22448 15166 22500
rect 15194 22448 15200 22500
rect 15252 22488 15258 22500
rect 16117 22491 16175 22497
rect 16117 22488 16129 22491
rect 15252 22460 16129 22488
rect 15252 22448 15258 22460
rect 16117 22457 16129 22460
rect 16163 22457 16175 22491
rect 16117 22451 16175 22457
rect 16316 22460 16988 22488
rect 7668 22392 10732 22420
rect 11698 22380 11704 22432
rect 11756 22380 11762 22432
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 16316 22420 16344 22460
rect 12032 22392 16344 22420
rect 12032 22380 12038 22392
rect 16390 22380 16396 22432
rect 16448 22380 16454 22432
rect 16960 22420 16988 22460
rect 18414 22448 18420 22500
rect 18472 22488 18478 22500
rect 19061 22491 19119 22497
rect 19061 22488 19073 22491
rect 18472 22460 19073 22488
rect 18472 22448 18478 22460
rect 19061 22457 19073 22460
rect 19107 22457 19119 22491
rect 19061 22451 19119 22457
rect 19242 22448 19248 22500
rect 19300 22488 19306 22500
rect 19720 22488 19748 22528
rect 20714 22516 20720 22568
rect 20772 22516 20778 22568
rect 20809 22559 20867 22565
rect 20809 22525 20821 22559
rect 20855 22525 20867 22559
rect 20809 22519 20867 22525
rect 19300 22460 19748 22488
rect 19300 22448 19306 22460
rect 20346 22448 20352 22500
rect 20404 22488 20410 22500
rect 20824 22488 20852 22519
rect 22462 22516 22468 22568
rect 22520 22516 22526 22568
rect 22557 22559 22615 22565
rect 22557 22525 22569 22559
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 20404 22460 20852 22488
rect 20404 22448 20410 22460
rect 22278 22448 22284 22500
rect 22336 22488 22342 22500
rect 22572 22488 22600 22519
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 22336 22460 22600 22488
rect 25041 22491 25099 22497
rect 22336 22448 22342 22460
rect 25041 22457 25053 22491
rect 25087 22488 25099 22491
rect 25406 22488 25412 22500
rect 25087 22460 25412 22488
rect 25087 22457 25099 22460
rect 25041 22451 25099 22457
rect 25406 22448 25412 22460
rect 25464 22448 25470 22500
rect 17586 22420 17592 22432
rect 16960 22392 17592 22420
rect 17586 22380 17592 22392
rect 17644 22380 17650 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18601 22423 18659 22429
rect 18601 22420 18613 22423
rect 17828 22392 18613 22420
rect 17828 22380 17834 22392
rect 18601 22389 18613 22392
rect 18647 22389 18659 22423
rect 18601 22383 18659 22389
rect 18966 22380 18972 22432
rect 19024 22420 19030 22432
rect 20714 22420 20720 22432
rect 19024 22392 20720 22420
rect 19024 22380 19030 22392
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 21358 22380 21364 22432
rect 21416 22380 21422 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22830 22420 22836 22432
rect 22051 22392 22836 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22830 22380 22836 22392
rect 22888 22380 22894 22432
rect 25314 22380 25320 22432
rect 25372 22380 25378 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 2498 22216 2504 22228
rect 2280 22188 2504 22216
rect 2280 22176 2286 22188
rect 2498 22176 2504 22188
rect 2556 22176 2562 22228
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 9582 22216 9588 22228
rect 4028 22188 9588 22216
rect 4028 22176 4034 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 11698 22216 11704 22228
rect 9732 22188 11704 22216
rect 9732 22176 9738 22188
rect 11698 22176 11704 22188
rect 11756 22176 11762 22228
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 14182 22216 14188 22228
rect 12768 22188 14188 22216
rect 12768 22176 12774 22188
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 14540 22219 14598 22225
rect 14540 22185 14552 22219
rect 14586 22216 14598 22219
rect 14918 22216 14924 22228
rect 14586 22188 14924 22216
rect 14586 22185 14598 22188
rect 14540 22179 14598 22185
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 15010 22176 15016 22228
rect 15068 22216 15074 22228
rect 15068 22188 16528 22216
rect 15068 22176 15074 22188
rect 1854 22108 1860 22160
rect 1912 22148 1918 22160
rect 10134 22148 10140 22160
rect 1912 22120 10140 22148
rect 1912 22108 1918 22120
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 14200 22120 14412 22148
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 1673 22083 1731 22089
rect 1673 22080 1685 22083
rect 1544 22052 1685 22080
rect 1544 22040 1550 22052
rect 1673 22049 1685 22052
rect 1719 22049 1731 22083
rect 1673 22043 1731 22049
rect 1688 21944 1716 22043
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 4264 22052 6040 22080
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2498 22012 2504 22024
rect 2271 21984 2504 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2498 21972 2504 21984
rect 2556 21972 2562 22024
rect 2590 21972 2596 22024
rect 2648 22012 2654 22024
rect 4264 22021 4292 22052
rect 4249 22015 4307 22021
rect 2648 21984 4108 22012
rect 2648 21972 2654 21984
rect 3970 21944 3976 21956
rect 1688 21916 3976 21944
rect 3970 21904 3976 21916
rect 4028 21904 4034 21956
rect 4080 21944 4108 21984
rect 4249 21981 4261 22015
rect 4295 21981 4307 22015
rect 4249 21975 4307 21981
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 21981 5411 22015
rect 5353 21975 5411 21981
rect 5368 21944 5396 21975
rect 4080 21916 5396 21944
rect 6012 21944 6040 22052
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 8404 22052 10057 22080
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 8404 21944 8432 22052
rect 10045 22049 10057 22052
rect 10091 22080 10103 22083
rect 10594 22080 10600 22092
rect 10091 22052 10600 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 10962 22040 10968 22092
rect 11020 22040 11026 22092
rect 11330 22040 11336 22092
rect 11388 22080 11394 22092
rect 14200 22080 14228 22120
rect 11388 22052 14228 22080
rect 11388 22040 11394 22052
rect 14274 22040 14280 22092
rect 14332 22040 14338 22092
rect 14384 22080 14412 22120
rect 16022 22108 16028 22160
rect 16080 22108 16086 22160
rect 15746 22080 15752 22092
rect 14384 22052 15752 22080
rect 15746 22040 15752 22052
rect 15804 22080 15810 22092
rect 16040 22080 16068 22108
rect 16500 22080 16528 22188
rect 17678 22176 17684 22228
rect 17736 22216 17742 22228
rect 18693 22219 18751 22225
rect 18693 22216 18705 22219
rect 17736 22188 18705 22216
rect 17736 22176 17742 22188
rect 18693 22185 18705 22188
rect 18739 22216 18751 22219
rect 19058 22216 19064 22228
rect 18739 22188 19064 22216
rect 18739 22185 18751 22188
rect 18693 22179 18751 22185
rect 19058 22176 19064 22188
rect 19116 22176 19122 22228
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20606 22219 20664 22225
rect 20606 22216 20618 22219
rect 20036 22188 20618 22216
rect 20036 22176 20042 22188
rect 20606 22185 20618 22188
rect 20652 22185 20664 22219
rect 20606 22179 20664 22185
rect 21910 22176 21916 22228
rect 21968 22216 21974 22228
rect 26878 22216 26884 22228
rect 21968 22188 26884 22216
rect 21968 22176 21974 22188
rect 26878 22176 26884 22188
rect 26936 22176 26942 22228
rect 23474 22148 23480 22160
rect 23216 22120 23480 22148
rect 16850 22080 16856 22092
rect 15804 22052 15976 22080
rect 16040 22052 16436 22080
rect 16500 22052 16856 22080
rect 15804 22040 15810 22052
rect 9030 21972 9036 22024
rect 9088 22012 9094 22024
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 9088 21984 10701 22012
rect 9088 21972 9094 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 13078 21972 13084 22024
rect 13136 21972 13142 22024
rect 15948 22012 15976 22052
rect 16408 22012 16436 22052
rect 16850 22040 16856 22052
rect 16908 22080 16914 22092
rect 17037 22083 17095 22089
rect 17037 22080 17049 22083
rect 16908 22052 17049 22080
rect 16908 22040 16914 22052
rect 17037 22049 17049 22052
rect 17083 22049 17095 22083
rect 17037 22043 17095 22049
rect 18230 22040 18236 22092
rect 18288 22040 18294 22092
rect 18690 22040 18696 22092
rect 18748 22080 18754 22092
rect 21266 22080 21272 22092
rect 18748 22052 21272 22080
rect 18748 22040 18754 22052
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 23216 22089 23244 22120
rect 23474 22108 23480 22120
rect 23532 22148 23538 22160
rect 24118 22148 24124 22160
rect 23532 22120 24124 22148
rect 23532 22108 23538 22120
rect 24118 22108 24124 22120
rect 24176 22108 24182 22160
rect 23201 22083 23259 22089
rect 23201 22049 23213 22083
rect 23247 22080 23259 22083
rect 23247 22052 23281 22080
rect 23247 22049 23259 22052
rect 23201 22043 23259 22049
rect 23750 22040 23756 22092
rect 23808 22080 23814 22092
rect 24029 22083 24087 22089
rect 24029 22080 24041 22083
rect 23808 22052 24041 22080
rect 23808 22040 23814 22052
rect 24029 22049 24041 22052
rect 24075 22049 24087 22083
rect 24029 22043 24087 22049
rect 25222 22040 25228 22092
rect 25280 22040 25286 22092
rect 16482 22012 16488 22024
rect 15948 21984 16344 22012
rect 16408 21984 16488 22012
rect 6012 21916 8432 21944
rect 8570 21904 8576 21956
rect 8628 21944 8634 21956
rect 9861 21947 9919 21953
rect 9861 21944 9873 21947
rect 8628 21916 9873 21944
rect 8628 21904 8634 21916
rect 9861 21913 9873 21916
rect 9907 21913 9919 21947
rect 9861 21907 9919 21913
rect 10870 21904 10876 21956
rect 10928 21944 10934 21956
rect 10928 21916 11454 21944
rect 10928 21904 10934 21916
rect 12342 21904 12348 21956
rect 12400 21944 12406 21956
rect 12400 21916 14412 21944
rect 12400 21904 12406 21916
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 3694 21876 3700 21888
rect 1627 21848 3700 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 3694 21836 3700 21848
rect 3752 21836 3758 21888
rect 3881 21879 3939 21885
rect 3881 21845 3893 21879
rect 3927 21876 3939 21879
rect 4246 21876 4252 21888
rect 3927 21848 4252 21876
rect 3927 21845 3939 21848
rect 3881 21839 3939 21845
rect 4246 21836 4252 21848
rect 4304 21836 4310 21888
rect 4893 21879 4951 21885
rect 4893 21845 4905 21879
rect 4939 21876 4951 21879
rect 5442 21876 5448 21888
rect 4939 21848 5448 21876
rect 4939 21845 4951 21848
rect 4893 21839 4951 21845
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 6454 21836 6460 21888
rect 6512 21876 6518 21888
rect 8938 21876 8944 21888
rect 6512 21848 8944 21876
rect 6512 21836 6518 21848
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 9217 21879 9275 21885
rect 9217 21845 9229 21879
rect 9263 21876 9275 21879
rect 9306 21876 9312 21888
rect 9263 21848 9312 21876
rect 9263 21845 9275 21848
rect 9217 21839 9275 21845
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 9493 21879 9551 21885
rect 9493 21876 9505 21879
rect 9456 21848 9505 21876
rect 9456 21836 9462 21848
rect 9493 21845 9505 21848
rect 9539 21845 9551 21879
rect 9493 21839 9551 21845
rect 9953 21879 10011 21885
rect 9953 21845 9965 21879
rect 9999 21876 10011 21879
rect 11790 21876 11796 21888
rect 9999 21848 11796 21876
rect 9999 21845 10011 21848
rect 9953 21839 10011 21845
rect 11790 21836 11796 21848
rect 11848 21836 11854 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 12250 21876 12256 21888
rect 12032 21848 12256 21876
rect 12032 21836 12038 21848
rect 12250 21836 12256 21848
rect 12308 21876 12314 21888
rect 12437 21879 12495 21885
rect 12437 21876 12449 21879
rect 12308 21848 12449 21876
rect 12308 21836 12314 21848
rect 12437 21845 12449 21848
rect 12483 21845 12495 21879
rect 12437 21839 12495 21845
rect 12526 21836 12532 21888
rect 12584 21876 12590 21888
rect 12713 21879 12771 21885
rect 12713 21876 12725 21879
rect 12584 21848 12725 21876
rect 12584 21836 12590 21848
rect 12713 21845 12725 21848
rect 12759 21845 12771 21879
rect 12713 21839 12771 21845
rect 13722 21836 13728 21888
rect 13780 21836 13786 21888
rect 14384 21876 14412 21916
rect 14550 21904 14556 21956
rect 14608 21944 14614 21956
rect 14608 21916 15042 21944
rect 14608 21904 14614 21916
rect 16022 21904 16028 21956
rect 16080 21944 16086 21956
rect 16206 21944 16212 21956
rect 16080 21916 16212 21944
rect 16080 21904 16086 21916
rect 16206 21904 16212 21916
rect 16264 21904 16270 21956
rect 16316 21944 16344 21984
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 18141 22015 18199 22021
rect 18141 22012 18153 22015
rect 16632 21984 18153 22012
rect 16632 21972 16638 21984
rect 18141 21981 18153 21984
rect 18187 22012 18199 22015
rect 18966 22012 18972 22024
rect 18187 21984 18972 22012
rect 18187 21981 18199 21984
rect 18141 21975 18199 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19518 21972 19524 22024
rect 19576 21972 19582 22024
rect 19610 21972 19616 22024
rect 19668 22012 19674 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19668 21984 20361 22012
rect 19668 21972 19674 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 21634 21972 21640 22024
rect 21692 22012 21698 22024
rect 22002 22012 22008 22024
rect 21692 21984 22008 22012
rect 21692 21972 21698 21984
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 23842 21972 23848 22024
rect 23900 21972 23906 22024
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 25590 22012 25596 22024
rect 24995 21984 25596 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 16945 21947 17003 21953
rect 16945 21944 16957 21947
rect 16316 21916 16957 21944
rect 16945 21913 16957 21916
rect 16991 21913 17003 21947
rect 16945 21907 17003 21913
rect 17494 21904 17500 21956
rect 17552 21944 17558 21956
rect 18877 21947 18935 21953
rect 18877 21944 18889 21947
rect 17552 21916 18889 21944
rect 17552 21904 17558 21916
rect 18877 21913 18889 21916
rect 18923 21913 18935 21947
rect 19981 21947 20039 21953
rect 19981 21944 19993 21947
rect 18877 21907 18935 21913
rect 19536 21916 19993 21944
rect 16485 21879 16543 21885
rect 16485 21876 16497 21879
rect 14384 21848 16497 21876
rect 16485 21845 16497 21848
rect 16531 21845 16543 21879
rect 16485 21839 16543 21845
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18049 21879 18107 21885
rect 18049 21876 18061 21879
rect 18012 21848 18061 21876
rect 18012 21836 18018 21848
rect 18049 21845 18061 21848
rect 18095 21845 18107 21879
rect 18049 21839 18107 21845
rect 19058 21836 19064 21888
rect 19116 21876 19122 21888
rect 19536 21876 19564 21916
rect 19981 21913 19993 21916
rect 20027 21944 20039 21947
rect 21082 21944 21088 21956
rect 20027 21916 21088 21944
rect 20027 21913 20039 21916
rect 19981 21907 20039 21913
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 23017 21947 23075 21953
rect 23017 21913 23029 21947
rect 23063 21944 23075 21947
rect 25774 21944 25780 21956
rect 23063 21916 25780 21944
rect 23063 21913 23075 21916
rect 23017 21907 23075 21913
rect 25774 21904 25780 21916
rect 25832 21904 25838 21956
rect 19116 21848 19564 21876
rect 19116 21836 19122 21848
rect 19610 21836 19616 21888
rect 19668 21836 19674 21888
rect 20714 21836 20720 21888
rect 20772 21876 20778 21888
rect 22002 21876 22008 21888
rect 20772 21848 22008 21876
rect 20772 21836 20778 21848
rect 22002 21836 22008 21848
rect 22060 21876 22066 21888
rect 22097 21879 22155 21885
rect 22097 21876 22109 21879
rect 22060 21848 22109 21876
rect 22060 21836 22066 21848
rect 22097 21845 22109 21848
rect 22143 21845 22155 21879
rect 22097 21839 22155 21845
rect 22462 21836 22468 21888
rect 22520 21876 22526 21888
rect 22557 21879 22615 21885
rect 22557 21876 22569 21879
rect 22520 21848 22569 21876
rect 22520 21836 22526 21848
rect 22557 21845 22569 21848
rect 22603 21845 22615 21879
rect 22557 21839 22615 21845
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 22925 21879 22983 21885
rect 22925 21876 22937 21879
rect 22704 21848 22937 21876
rect 22704 21836 22710 21848
rect 22925 21845 22937 21848
rect 22971 21845 22983 21879
rect 22925 21839 22983 21845
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23808 21848 24593 21876
rect 23808 21836 23814 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 26602 21876 26608 21888
rect 25087 21848 26608 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 2317 21675 2375 21681
rect 2317 21672 2329 21675
rect 1636 21644 2329 21672
rect 1636 21632 1642 21644
rect 2317 21641 2329 21644
rect 2363 21641 2375 21675
rect 2317 21635 2375 21641
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 4028 21644 11192 21672
rect 4028 21632 4034 21644
rect 1946 21564 1952 21616
rect 2004 21604 2010 21616
rect 2866 21604 2872 21616
rect 2004 21576 2872 21604
rect 2004 21564 2010 21576
rect 2866 21564 2872 21576
rect 2924 21564 2930 21616
rect 6730 21604 6736 21616
rect 2976 21576 6736 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 1762 21536 1768 21548
rect 1719 21508 1768 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 2976 21545 3004 21576
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 7834 21564 7840 21616
rect 7892 21604 7898 21616
rect 9309 21607 9367 21613
rect 9309 21604 9321 21607
rect 7892 21576 9321 21604
rect 7892 21564 7898 21576
rect 9309 21573 9321 21576
rect 9355 21573 9367 21607
rect 10778 21604 10784 21616
rect 10534 21576 10784 21604
rect 9309 21567 9367 21573
rect 10778 21564 10784 21576
rect 10836 21604 10842 21616
rect 11057 21607 11115 21613
rect 11057 21604 11069 21607
rect 10836 21576 11069 21604
rect 10836 21564 10842 21576
rect 11057 21573 11069 21576
rect 11103 21573 11115 21607
rect 11164 21604 11192 21644
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 11296 21644 11897 21672
rect 11296 21632 11302 21644
rect 11885 21641 11897 21644
rect 11931 21641 11943 21675
rect 11885 21635 11943 21641
rect 12161 21675 12219 21681
rect 12161 21641 12173 21675
rect 12207 21672 12219 21675
rect 12250 21672 12256 21684
rect 12207 21644 12256 21672
rect 12207 21641 12219 21644
rect 12161 21635 12219 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 12526 21632 12532 21684
rect 12584 21672 12590 21684
rect 13265 21675 13323 21681
rect 13265 21672 13277 21675
rect 12584 21644 13277 21672
rect 12584 21632 12590 21644
rect 13265 21641 13277 21644
rect 13311 21641 13323 21675
rect 14090 21672 14096 21684
rect 13265 21635 13323 21641
rect 13464 21644 14096 21672
rect 13464 21604 13492 21644
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 14182 21632 14188 21684
rect 14240 21632 14246 21684
rect 14277 21675 14335 21681
rect 14277 21641 14289 21675
rect 14323 21672 14335 21675
rect 17678 21672 17684 21684
rect 14323 21644 17684 21672
rect 14323 21641 14335 21644
rect 14277 21635 14335 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 18690 21672 18696 21684
rect 18064 21644 18696 21672
rect 11164 21576 13492 21604
rect 13541 21607 13599 21613
rect 11057 21567 11115 21573
rect 13541 21573 13553 21607
rect 13587 21604 13599 21607
rect 14458 21604 14464 21616
rect 13587 21576 14464 21604
rect 13587 21573 13599 21576
rect 13541 21567 13599 21573
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 3694 21496 3700 21548
rect 3752 21536 3758 21548
rect 4614 21536 4620 21548
rect 3752 21508 4620 21536
rect 3752 21496 3758 21508
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21536 4859 21539
rect 5258 21536 5264 21548
rect 4847 21508 5264 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 7098 21496 7104 21548
rect 7156 21536 7162 21548
rect 7193 21539 7251 21545
rect 7193 21536 7205 21539
rect 7156 21508 7205 21536
rect 7156 21496 7162 21508
rect 7193 21505 7205 21508
rect 7239 21505 7251 21539
rect 7193 21499 7251 21505
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 11072 21536 11100 21567
rect 14458 21564 14464 21576
rect 14516 21564 14522 21616
rect 15746 21564 15752 21616
rect 15804 21604 15810 21616
rect 16393 21607 16451 21613
rect 16393 21604 16405 21607
rect 15804 21576 16405 21604
rect 15804 21564 15810 21576
rect 16393 21573 16405 21576
rect 16439 21573 16451 21607
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 16393 21567 16451 21573
rect 16500 21576 17417 21604
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 11072 21508 11253 21536
rect 11241 21505 11253 21508
rect 11287 21536 11299 21539
rect 11514 21536 11520 21548
rect 11287 21508 11520 21536
rect 11287 21505 11299 21508
rect 11241 21499 11299 21505
rect 11514 21496 11520 21508
rect 11572 21536 11578 21548
rect 11701 21539 11759 21545
rect 11701 21536 11713 21539
rect 11572 21508 11713 21536
rect 11572 21496 11578 21508
rect 11701 21505 11713 21508
rect 11747 21536 11759 21539
rect 12526 21536 12532 21548
rect 11747 21508 12532 21536
rect 11747 21505 11759 21508
rect 11701 21499 11759 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 12621 21539 12679 21545
rect 12621 21505 12633 21539
rect 12667 21505 12679 21539
rect 12621 21499 12679 21505
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 6549 21471 6607 21477
rect 6549 21437 6561 21471
rect 6595 21437 6607 21471
rect 6549 21431 6607 21437
rect 2866 21360 2872 21412
rect 2924 21400 2930 21412
rect 6454 21400 6460 21412
rect 2924 21372 6460 21400
rect 2924 21360 2930 21372
rect 6454 21360 6460 21372
rect 6512 21360 6518 21412
rect 6564 21400 6592 21431
rect 7466 21428 7472 21480
rect 7524 21468 7530 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7524 21440 7665 21468
rect 7524 21428 7530 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 12158 21468 12164 21480
rect 7653 21431 7711 21437
rect 9140 21440 12164 21468
rect 9140 21400 9168 21440
rect 12158 21428 12164 21440
rect 12216 21428 12222 21480
rect 12250 21428 12256 21480
rect 12308 21468 12314 21480
rect 12636 21468 12664 21499
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 14918 21536 14924 21548
rect 14608 21508 14924 21536
rect 14608 21496 14614 21508
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21505 15439 21539
rect 16209 21539 16267 21545
rect 16209 21536 16221 21539
rect 15381 21499 15439 21505
rect 15580 21508 16221 21536
rect 12308 21440 12664 21468
rect 12713 21471 12771 21477
rect 12308 21428 12314 21440
rect 12713 21437 12725 21471
rect 12759 21437 12771 21471
rect 12713 21431 12771 21437
rect 6564 21372 9168 21400
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 10781 21403 10839 21409
rect 10781 21400 10793 21403
rect 10652 21372 10793 21400
rect 10652 21360 10658 21372
rect 10781 21369 10793 21372
rect 10827 21369 10839 21403
rect 10781 21363 10839 21369
rect 11609 21403 11667 21409
rect 11609 21369 11621 21403
rect 11655 21400 11667 21403
rect 12728 21400 12756 21431
rect 12802 21428 12808 21480
rect 12860 21428 12866 21480
rect 13078 21428 13084 21480
rect 13136 21468 13142 21480
rect 14461 21471 14519 21477
rect 14461 21468 14473 21471
rect 13136 21440 14473 21468
rect 13136 21428 13142 21440
rect 14461 21437 14473 21440
rect 14507 21468 14519 21471
rect 15286 21468 15292 21480
rect 14507 21440 15292 21468
rect 14507 21437 14519 21440
rect 14461 21431 14519 21437
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 15396 21412 15424 21499
rect 15580 21480 15608 21508
rect 16209 21505 16221 21508
rect 16255 21505 16267 21539
rect 16209 21499 16267 21505
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 16500 21536 16528 21576
rect 17405 21573 17417 21576
rect 17451 21604 17463 21607
rect 18064 21604 18092 21644
rect 18690 21632 18696 21644
rect 18748 21632 18754 21684
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21634 21672 21640 21684
rect 21140 21644 21640 21672
rect 21140 21632 21146 21644
rect 21634 21632 21640 21644
rect 21692 21632 21698 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22738 21672 22744 21684
rect 22244 21644 22744 21672
rect 22244 21632 22250 21644
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 24946 21632 24952 21684
rect 25004 21672 25010 21684
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 25004 21644 25145 21672
rect 25004 21632 25010 21644
rect 25133 21641 25145 21644
rect 25179 21641 25191 21675
rect 25133 21635 25191 21641
rect 25501 21675 25559 21681
rect 25501 21641 25513 21675
rect 25547 21672 25559 21675
rect 25774 21672 25780 21684
rect 25547 21644 25780 21672
rect 25547 21641 25559 21644
rect 25501 21635 25559 21641
rect 25774 21632 25780 21644
rect 25832 21632 25838 21684
rect 17451 21576 18092 21604
rect 18156 21576 22600 21604
rect 17451 21573 17463 21576
rect 17405 21567 17463 21573
rect 16356 21508 16528 21536
rect 16761 21539 16819 21545
rect 16356 21496 16362 21508
rect 16761 21505 16773 21539
rect 16807 21536 16819 21539
rect 17034 21536 17040 21548
rect 16807 21508 17040 21536
rect 16807 21505 16819 21508
rect 16761 21499 16819 21505
rect 17034 21496 17040 21508
rect 17092 21496 17098 21548
rect 18156 21536 18184 21576
rect 17420 21508 18184 21536
rect 18233 21539 18291 21545
rect 17420 21480 17448 21508
rect 18233 21505 18245 21539
rect 18279 21536 18291 21539
rect 19058 21536 19064 21548
rect 18279 21508 19064 21536
rect 18279 21505 18291 21508
rect 18233 21499 18291 21505
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 20806 21496 20812 21548
rect 20864 21496 20870 21548
rect 20990 21496 20996 21548
rect 21048 21536 21054 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 21048 21508 22385 21536
rect 21048 21496 21054 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 15562 21428 15568 21480
rect 15620 21428 15626 21480
rect 17310 21468 17316 21480
rect 15856 21440 17316 21468
rect 14182 21400 14188 21412
rect 11655 21372 12664 21400
rect 12728 21372 14188 21400
rect 11655 21369 11667 21372
rect 11609 21363 11667 21369
rect 4706 21292 4712 21344
rect 4764 21332 4770 21344
rect 6086 21332 6092 21344
rect 4764 21304 6092 21332
rect 4764 21292 4770 21304
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 9398 21332 9404 21344
rect 8536 21304 9404 21332
rect 8536 21292 8542 21304
rect 9398 21292 9404 21304
rect 9456 21292 9462 21344
rect 12250 21292 12256 21344
rect 12308 21292 12314 21344
rect 12636 21332 12664 21372
rect 14182 21360 14188 21372
rect 14240 21360 14246 21412
rect 15378 21360 15384 21412
rect 15436 21400 15442 21412
rect 15746 21400 15752 21412
rect 15436 21372 15752 21400
rect 15436 21360 15442 21372
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 13630 21332 13636 21344
rect 12636 21304 13636 21332
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 14366 21332 14372 21344
rect 13863 21304 14372 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 15013 21335 15071 21341
rect 15013 21301 15025 21335
rect 15059 21332 15071 21335
rect 15856 21332 15884 21440
rect 17310 21428 17316 21440
rect 17368 21428 17374 21480
rect 17402 21428 17408 21480
rect 17460 21428 17466 21480
rect 17494 21428 17500 21480
rect 17552 21428 17558 21480
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 16942 21360 16948 21412
rect 17000 21400 17006 21412
rect 17604 21400 17632 21431
rect 18414 21428 18420 21480
rect 18472 21468 18478 21480
rect 19610 21468 19616 21480
rect 18472 21440 19616 21468
rect 18472 21428 18478 21440
rect 19610 21428 19616 21440
rect 19668 21428 19674 21480
rect 19702 21428 19708 21480
rect 19760 21468 19766 21480
rect 19760 21440 20852 21468
rect 19760 21428 19766 21440
rect 17000 21372 17632 21400
rect 17000 21360 17006 21372
rect 18598 21360 18604 21412
rect 18656 21400 18662 21412
rect 20714 21400 20720 21412
rect 18656 21372 20720 21400
rect 18656 21360 18662 21372
rect 20714 21360 20720 21372
rect 20772 21360 20778 21412
rect 20824 21400 20852 21440
rect 20898 21428 20904 21480
rect 20956 21428 20962 21480
rect 21085 21471 21143 21477
rect 21085 21437 21097 21471
rect 21131 21468 21143 21471
rect 21358 21468 21364 21480
rect 21131 21440 21364 21468
rect 21131 21437 21143 21440
rect 21085 21431 21143 21437
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 22572 21477 22600 21576
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 24762 21496 24768 21548
rect 24820 21496 24826 21548
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22066 21440 22477 21468
rect 22066 21400 22094 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 22557 21431 22615 21437
rect 23216 21440 23673 21468
rect 20824 21372 22094 21400
rect 22738 21360 22744 21412
rect 22796 21400 22802 21412
rect 23216 21409 23244 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23201 21403 23259 21409
rect 23201 21400 23213 21403
rect 22796 21372 23213 21400
rect 22796 21360 22802 21372
rect 23201 21369 23213 21372
rect 23247 21369 23259 21403
rect 23201 21363 23259 21369
rect 15059 21304 15884 21332
rect 16117 21335 16175 21341
rect 15059 21301 15071 21304
rect 15013 21295 15071 21301
rect 16117 21301 16129 21335
rect 16163 21332 16175 21335
rect 16574 21332 16580 21344
rect 16163 21304 16580 21332
rect 16163 21301 16175 21304
rect 16117 21295 16175 21301
rect 16574 21292 16580 21304
rect 16632 21332 16638 21344
rect 16758 21332 16764 21344
rect 16632 21304 16764 21332
rect 16632 21292 16638 21304
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 17862 21332 17868 21344
rect 17083 21304 17868 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19521 21295 19579 21301
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 20036 21304 20453 21332
rect 20036 21292 20042 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 21542 21292 21548 21344
rect 21600 21292 21606 21344
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21968 21304 22017 21332
rect 21968 21292 21974 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22005 21295 22063 21301
rect 23109 21335 23167 21341
rect 23109 21301 23121 21335
rect 23155 21332 23167 21335
rect 24762 21332 24768 21344
rect 23155 21304 24768 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 24762 21292 24768 21304
rect 24820 21292 24826 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 4706 21128 4712 21140
rect 1820 21100 4712 21128
rect 1820 21088 1826 21100
rect 4706 21088 4712 21100
rect 4764 21088 4770 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 4816 21100 13645 21128
rect 4816 21060 4844 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 14182 21088 14188 21140
rect 14240 21128 14246 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 14240 21100 16681 21128
rect 14240 21088 14246 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 17586 21088 17592 21140
rect 17644 21128 17650 21140
rect 17865 21131 17923 21137
rect 17865 21128 17877 21131
rect 17644 21100 17877 21128
rect 17644 21088 17650 21100
rect 17865 21097 17877 21100
rect 17911 21097 17923 21131
rect 17865 21091 17923 21097
rect 18322 21088 18328 21140
rect 18380 21128 18386 21140
rect 20806 21128 20812 21140
rect 18380 21100 20812 21128
rect 18380 21088 18386 21100
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 22646 21128 22652 21140
rect 21744 21100 22652 21128
rect 2332 21032 4844 21060
rect 6457 21063 6515 21069
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 2332 20924 2360 21032
rect 6457 21029 6469 21063
rect 6503 21060 6515 21063
rect 6914 21060 6920 21072
rect 6503 21032 6920 21060
rect 6503 21029 6515 21032
rect 6457 21023 6515 21029
rect 6914 21020 6920 21032
rect 6972 21020 6978 21072
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 10226 21060 10232 21072
rect 9364 21032 10232 21060
rect 9364 21020 9370 21032
rect 10226 21020 10232 21032
rect 10284 21020 10290 21072
rect 12897 21063 12955 21069
rect 12897 21029 12909 21063
rect 12943 21060 12955 21063
rect 15010 21060 15016 21072
rect 12943 21032 15016 21060
rect 12943 21029 12955 21032
rect 12897 21023 12955 21029
rect 15010 21020 15016 21032
rect 15068 21020 15074 21072
rect 15473 21063 15531 21069
rect 15473 21029 15485 21063
rect 15519 21029 15531 21063
rect 16758 21060 16764 21072
rect 15473 21023 15531 21029
rect 15948 21032 16764 21060
rect 4890 20952 4896 21004
rect 4948 20952 4954 21004
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 6880 20964 7389 20992
rect 6880 20952 6886 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7377 20955 7435 20961
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 8846 20992 8852 21004
rect 8628 20964 8852 20992
rect 8628 20952 8634 20964
rect 8846 20952 8852 20964
rect 8904 20952 8910 21004
rect 9030 20952 9036 21004
rect 9088 20992 9094 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 9088 20964 11161 20992
rect 9088 20952 9094 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 15488 20992 15516 21023
rect 15948 21001 15976 21032
rect 16758 21020 16764 21032
rect 16816 21060 16822 21072
rect 17678 21060 17684 21072
rect 16816 21032 17684 21060
rect 16816 21020 16822 21032
rect 17678 21020 17684 21032
rect 17736 21020 17742 21072
rect 18414 21020 18420 21072
rect 18472 21060 18478 21072
rect 18472 21032 19564 21060
rect 18472 21020 18478 21032
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 11848 20964 15516 20992
rect 15580 20964 15945 20992
rect 11848 20952 11854 20964
rect 2271 20896 2360 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 2406 20884 2412 20936
rect 2464 20924 2470 20936
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2464 20896 2973 20924
rect 2464 20884 2470 20896
rect 2961 20893 2973 20896
rect 3007 20893 3019 20927
rect 2961 20887 3019 20893
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 1581 20859 1639 20865
rect 1581 20825 1593 20859
rect 1627 20856 1639 20859
rect 1946 20856 1952 20868
rect 1627 20828 1952 20856
rect 1627 20825 1639 20828
rect 1581 20819 1639 20825
rect 1946 20816 1952 20828
rect 2004 20816 2010 20868
rect 1394 20748 1400 20800
rect 1452 20788 1458 20800
rect 1673 20791 1731 20797
rect 1673 20788 1685 20791
rect 1452 20760 1685 20788
rect 1452 20748 1458 20760
rect 1673 20757 1685 20760
rect 1719 20788 1731 20791
rect 2682 20788 2688 20800
rect 1719 20760 2688 20788
rect 1719 20757 1731 20760
rect 1673 20751 1731 20757
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 4080 20788 4108 20887
rect 4246 20884 4252 20936
rect 4304 20924 4310 20936
rect 5813 20927 5871 20933
rect 5813 20924 5825 20927
rect 4304 20896 5825 20924
rect 4304 20884 4310 20896
rect 5813 20893 5825 20896
rect 5859 20893 5871 20927
rect 5813 20887 5871 20893
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7282 20924 7288 20936
rect 7147 20896 7288 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 5828 20856 5856 20887
rect 7282 20884 7288 20896
rect 7340 20884 7346 20936
rect 7558 20884 7564 20936
rect 7616 20924 7622 20936
rect 8386 20924 8392 20936
rect 7616 20896 8392 20924
rect 7616 20884 7622 20896
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 9122 20924 9128 20936
rect 8803 20896 9128 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 9398 20884 9404 20936
rect 9456 20884 9462 20936
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20924 10655 20927
rect 11054 20924 11060 20936
rect 10643 20896 11060 20924
rect 10643 20893 10655 20896
rect 10597 20887 10655 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 12952 20896 13553 20924
rect 12952 20884 12958 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14458 20924 14464 20936
rect 14323 20896 14464 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14458 20884 14464 20896
rect 14516 20884 14522 20936
rect 15580 20924 15608 20964
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 15933 20955 15991 20961
rect 16114 20952 16120 21004
rect 16172 20952 16178 21004
rect 16574 20952 16580 21004
rect 16632 20992 16638 21004
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 16632 20964 17233 20992
rect 16632 20952 16638 20964
rect 17221 20961 17233 20964
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 18322 20952 18328 21004
rect 18380 20952 18386 21004
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 19536 20992 19564 21032
rect 20714 21020 20720 21072
rect 20772 21060 20778 21072
rect 20772 21032 21312 21060
rect 20772 21020 20778 21032
rect 19702 20992 19708 21004
rect 19536 20964 19708 20992
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20346 20952 20352 21004
rect 20404 20992 20410 21004
rect 21177 20995 21235 21001
rect 21177 20992 21189 20995
rect 20404 20964 21189 20992
rect 20404 20952 20410 20964
rect 21177 20961 21189 20964
rect 21223 20961 21235 20995
rect 21284 20992 21312 21032
rect 21744 20992 21772 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 22833 21131 22891 21137
rect 22833 21097 22845 21131
rect 22879 21128 22891 21131
rect 22922 21128 22928 21140
rect 22879 21100 22928 21128
rect 22879 21097 22891 21100
rect 22833 21091 22891 21097
rect 22922 21088 22928 21100
rect 22980 21088 22986 21140
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 22060 21032 23428 21060
rect 22060 21020 22066 21032
rect 21284 20964 21772 20992
rect 21177 20955 21235 20961
rect 21910 20952 21916 21004
rect 21968 20992 21974 21004
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 21968 20964 22201 20992
rect 21968 20952 21974 20964
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 22830 20952 22836 21004
rect 22888 20992 22894 21004
rect 23400 21001 23428 21032
rect 23293 20995 23351 21001
rect 23293 20992 23305 20995
rect 22888 20964 23305 20992
rect 22888 20952 22894 20964
rect 23293 20961 23305 20964
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 24854 20952 24860 21004
rect 24912 20992 24918 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24912 20964 25053 20992
rect 24912 20952 24918 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20992 25283 20995
rect 25406 20992 25412 21004
rect 25271 20964 25412 20992
rect 25271 20961 25283 20964
rect 25225 20955 25283 20961
rect 25406 20952 25412 20964
rect 25464 20992 25470 21004
rect 26786 20992 26792 21004
rect 25464 20964 26792 20992
rect 25464 20952 25470 20964
rect 26786 20952 26792 20964
rect 26844 20952 26850 21004
rect 15396 20896 15608 20924
rect 8294 20856 8300 20868
rect 5828 20828 8300 20856
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 11425 20859 11483 20865
rect 11425 20856 11437 20859
rect 8628 20828 11437 20856
rect 8628 20816 8634 20828
rect 11425 20825 11437 20828
rect 11471 20825 11483 20859
rect 11425 20819 11483 20825
rect 11514 20816 11520 20868
rect 11572 20856 11578 20868
rect 11572 20828 11914 20856
rect 11572 20816 11578 20828
rect 14090 20816 14096 20868
rect 14148 20856 14154 20868
rect 15396 20856 15424 20896
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 18598 20924 18604 20936
rect 15712 20896 18604 20924
rect 15712 20884 15718 20896
rect 18598 20884 18604 20896
rect 18656 20884 18662 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 22097 20927 22155 20933
rect 22097 20924 22109 20927
rect 21140 20896 22109 20924
rect 21140 20884 21146 20896
rect 22097 20893 22109 20896
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 23201 20927 23259 20933
rect 23201 20924 23213 20927
rect 22612 20896 23213 20924
rect 22612 20884 22618 20896
rect 23201 20893 23213 20896
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 14148 20828 15424 20856
rect 14148 20816 14154 20828
rect 15470 20816 15476 20868
rect 15528 20856 15534 20868
rect 16206 20856 16212 20868
rect 15528 20828 16212 20856
rect 15528 20816 15534 20828
rect 16206 20816 16212 20828
rect 16264 20856 16270 20868
rect 18233 20859 18291 20865
rect 16264 20828 17172 20856
rect 16264 20816 16270 20828
rect 6454 20788 6460 20800
rect 4080 20760 6460 20788
rect 6454 20748 6460 20760
rect 6512 20748 6518 20800
rect 6638 20748 6644 20800
rect 6696 20788 6702 20800
rect 10413 20791 10471 20797
rect 10413 20788 10425 20791
rect 6696 20760 10425 20788
rect 6696 20748 6702 20760
rect 10413 20757 10425 20760
rect 10459 20757 10471 20791
rect 10413 20751 10471 20757
rect 10594 20748 10600 20800
rect 10652 20788 10658 20800
rect 14550 20788 14556 20800
rect 10652 20760 14556 20788
rect 10652 20748 10658 20760
rect 14550 20748 14556 20760
rect 14608 20748 14614 20800
rect 14918 20748 14924 20800
rect 14976 20748 14982 20800
rect 15562 20748 15568 20800
rect 15620 20788 15626 20800
rect 15841 20791 15899 20797
rect 15841 20788 15853 20791
rect 15620 20760 15853 20788
rect 15620 20748 15626 20760
rect 15841 20757 15853 20760
rect 15887 20757 15899 20791
rect 15841 20751 15899 20757
rect 17034 20748 17040 20800
rect 17092 20748 17098 20800
rect 17144 20797 17172 20828
rect 18233 20825 18245 20859
rect 18279 20856 18291 20859
rect 18279 20828 19656 20856
rect 18279 20825 18291 20828
rect 18233 20819 18291 20825
rect 17129 20791 17187 20797
rect 17129 20757 17141 20791
rect 17175 20788 17187 20791
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 17175 20760 18889 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 19628 20788 19656 20828
rect 19702 20816 19708 20868
rect 19760 20816 19766 20868
rect 20162 20816 20168 20868
rect 20220 20816 20226 20868
rect 21008 20828 22416 20856
rect 21008 20788 21036 20828
rect 19628 20760 21036 20788
rect 18877 20751 18935 20757
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 21637 20791 21695 20797
rect 21637 20788 21649 20791
rect 21324 20760 21649 20788
rect 21324 20748 21330 20760
rect 21637 20757 21649 20760
rect 21683 20757 21695 20791
rect 21637 20751 21695 20757
rect 22002 20748 22008 20800
rect 22060 20748 22066 20800
rect 22388 20788 22416 20828
rect 22462 20816 22468 20868
rect 22520 20856 22526 20868
rect 24949 20859 25007 20865
rect 24949 20856 24961 20859
rect 22520 20828 24961 20856
rect 22520 20816 22526 20828
rect 24949 20825 24961 20828
rect 24995 20825 25007 20859
rect 24949 20819 25007 20825
rect 23566 20788 23572 20800
rect 22388 20760 23572 20788
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 23934 20748 23940 20800
rect 23992 20748 23998 20800
rect 24026 20748 24032 20800
rect 24084 20748 24090 20800
rect 24578 20748 24584 20800
rect 24636 20748 24642 20800
rect 25406 20748 25412 20800
rect 25464 20788 25470 20800
rect 25590 20788 25596 20800
rect 25464 20760 25596 20788
rect 25464 20748 25470 20760
rect 25590 20748 25596 20760
rect 25648 20748 25654 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 5997 20587 6055 20593
rect 5997 20553 6009 20587
rect 6043 20584 6055 20587
rect 6914 20584 6920 20596
rect 6043 20556 6920 20584
rect 6043 20553 6055 20556
rect 5997 20547 6055 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7466 20544 7472 20596
rect 7524 20544 7530 20596
rect 12802 20584 12808 20596
rect 7852 20556 12808 20584
rect 7558 20516 7564 20528
rect 4908 20488 7564 20516
rect 1854 20408 1860 20460
rect 1912 20408 1918 20460
rect 4908 20457 4936 20488
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 4893 20451 4951 20457
rect 3099 20420 4844 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 1578 20340 1584 20392
rect 1636 20340 1642 20392
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 2832 20352 3341 20380
rect 2832 20340 2838 20352
rect 3329 20349 3341 20352
rect 3375 20349 3387 20383
rect 3329 20343 3387 20349
rect 4816 20312 4844 20420
rect 4893 20417 4905 20451
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 5994 20448 6000 20460
rect 5399 20420 6000 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 5994 20408 6000 20420
rect 6052 20408 6058 20460
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6457 20451 6515 20457
rect 6457 20448 6469 20451
rect 6144 20420 6469 20448
rect 6144 20408 6150 20420
rect 6457 20417 6469 20420
rect 6503 20417 6515 20451
rect 6457 20411 6515 20417
rect 6822 20408 6828 20460
rect 6880 20408 6886 20460
rect 6914 20408 6920 20460
rect 6972 20448 6978 20460
rect 7742 20448 7748 20460
rect 6972 20420 7748 20448
rect 6972 20408 6978 20420
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 7852 20448 7880 20556
rect 12802 20544 12808 20556
rect 12860 20584 12866 20596
rect 13354 20584 13360 20596
rect 12860 20556 13360 20584
rect 12860 20544 12866 20556
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14182 20544 14188 20596
rect 14240 20584 14246 20596
rect 16482 20584 16488 20596
rect 14240 20556 16488 20584
rect 14240 20544 14246 20556
rect 16482 20544 16488 20556
rect 16540 20584 16546 20596
rect 16540 20556 16988 20584
rect 16540 20544 16546 20556
rect 8570 20476 8576 20528
rect 8628 20476 8634 20528
rect 9582 20516 9588 20528
rect 8680 20488 9588 20516
rect 7917 20451 7975 20457
rect 7917 20448 7929 20451
rect 7852 20420 7929 20448
rect 7917 20417 7929 20420
rect 7963 20417 7975 20451
rect 7917 20411 7975 20417
rect 8110 20408 8116 20460
rect 8168 20448 8174 20460
rect 8680 20448 8708 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 11149 20519 11207 20525
rect 11149 20516 11161 20519
rect 10534 20488 11161 20516
rect 11149 20485 11161 20488
rect 11195 20516 11207 20519
rect 11333 20519 11391 20525
rect 11333 20516 11345 20519
rect 11195 20488 11345 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 11333 20485 11345 20488
rect 11379 20516 11391 20519
rect 11514 20516 11520 20528
rect 11379 20488 11520 20516
rect 11379 20485 11391 20488
rect 11333 20479 11391 20485
rect 11514 20476 11520 20488
rect 11572 20516 11578 20528
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 11572 20488 11713 20516
rect 11572 20476 11578 20488
rect 11701 20485 11713 20488
rect 11747 20485 11759 20519
rect 11701 20479 11759 20485
rect 12437 20519 12495 20525
rect 12437 20485 12449 20519
rect 12483 20516 12495 20519
rect 12618 20516 12624 20528
rect 12483 20488 12624 20516
rect 12483 20485 12495 20488
rect 12437 20479 12495 20485
rect 8168 20420 8708 20448
rect 8168 20408 8174 20420
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 11238 20448 11244 20460
rect 11112 20420 11244 20448
rect 11112 20408 11118 20420
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11716 20448 11744 20479
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 13814 20516 13820 20528
rect 13556 20488 13820 20516
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 11716 20420 13185 20448
rect 13173 20417 13185 20420
rect 13219 20448 13231 20451
rect 13446 20448 13452 20460
rect 13219 20420 13452 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13556 20457 13584 20488
rect 13814 20476 13820 20488
rect 13872 20516 13878 20528
rect 14200 20516 14228 20544
rect 13872 20488 14228 20516
rect 13872 20476 13878 20488
rect 16298 20476 16304 20528
rect 16356 20476 16362 20528
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 14950 20420 15240 20448
rect 13541 20411 13599 20417
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 5500 20352 9321 20380
rect 5500 20340 5506 20352
rect 9309 20349 9321 20352
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 12250 20380 12256 20392
rect 9456 20352 12256 20380
rect 9456 20340 9462 20352
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 8294 20312 8300 20324
rect 4816 20284 8300 20312
rect 8294 20272 8300 20284
rect 8352 20272 8358 20324
rect 10410 20272 10416 20324
rect 10468 20312 10474 20324
rect 11974 20312 11980 20324
rect 10468 20284 11980 20312
rect 10468 20272 10474 20284
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 12544 20312 12572 20343
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 15102 20380 15108 20392
rect 13863 20352 15108 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 12544 20284 13676 20312
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4709 20247 4767 20253
rect 4709 20244 4721 20247
rect 4028 20216 4721 20244
rect 4028 20204 4034 20216
rect 4709 20213 4721 20216
rect 4755 20213 4767 20247
rect 4709 20207 4767 20213
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 10781 20247 10839 20253
rect 10781 20244 10793 20247
rect 7984 20216 10793 20244
rect 7984 20204 7990 20216
rect 10781 20213 10793 20216
rect 10827 20244 10839 20247
rect 11054 20244 11060 20256
rect 10827 20216 11060 20244
rect 10827 20213 10839 20216
rect 10781 20207 10839 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11480 20216 11529 20244
rect 11480 20204 11486 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 11790 20204 11796 20256
rect 11848 20244 11854 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11848 20216 12081 20244
rect 11848 20204 11854 20216
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 13648 20244 13676 20284
rect 15010 20272 15016 20324
rect 15068 20312 15074 20324
rect 15212 20312 15240 20420
rect 16114 20408 16120 20460
rect 16172 20408 16178 20460
rect 16960 20457 16988 20556
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 20162 20584 20168 20596
rect 19904 20556 20168 20584
rect 17218 20476 17224 20528
rect 17276 20476 17282 20528
rect 19904 20516 19932 20556
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 22002 20584 22008 20596
rect 21600 20556 22008 20584
rect 21600 20544 21606 20556
rect 22002 20544 22008 20556
rect 22060 20584 22066 20596
rect 23109 20587 23167 20593
rect 23109 20584 23121 20587
rect 22060 20556 23121 20584
rect 22060 20544 22066 20556
rect 23109 20553 23121 20556
rect 23155 20553 23167 20587
rect 23109 20547 23167 20553
rect 18892 20488 20010 20516
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 15286 20340 15292 20392
rect 15344 20340 15350 20392
rect 18340 20380 18368 20434
rect 18892 20380 18920 20488
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22465 20519 22523 20525
rect 22465 20516 22477 20519
rect 22152 20488 22477 20516
rect 22152 20476 22158 20488
rect 22465 20485 22477 20488
rect 22511 20485 22523 20519
rect 22465 20479 22523 20485
rect 24762 20476 24768 20528
rect 24820 20476 24826 20528
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 22370 20448 22376 20460
rect 21508 20420 22376 20448
rect 21508 20408 21514 20420
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22557 20451 22615 20457
rect 22557 20417 22569 20451
rect 22603 20448 22615 20451
rect 22830 20448 22836 20460
rect 22603 20420 22836 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 22830 20408 22836 20420
rect 22888 20408 22894 20460
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 16408 20352 18920 20380
rect 16408 20324 16436 20352
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 20254 20380 20260 20392
rect 19567 20352 20260 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 20806 20340 20812 20392
rect 20864 20380 20870 20392
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20864 20352 21281 20380
rect 20864 20340 20870 20352
rect 21269 20349 21281 20352
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20380 23811 20383
rect 24210 20380 24216 20392
rect 23799 20352 24216 20380
rect 23799 20349 23811 20352
rect 23753 20343 23811 20349
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 15068 20284 15577 20312
rect 15068 20272 15074 20284
rect 15565 20281 15577 20284
rect 15611 20312 15623 20315
rect 16390 20312 16396 20324
rect 15611 20284 16396 20312
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 22278 20312 22284 20324
rect 21008 20284 22284 20312
rect 15470 20244 15476 20256
rect 13648 20216 15476 20244
rect 12069 20207 12127 20213
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 19702 20204 19708 20256
rect 19760 20244 19766 20256
rect 21008 20253 21036 20284
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 22664 20312 22692 20343
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 22612 20284 22692 20312
rect 22612 20272 22618 20284
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 19760 20216 21005 20244
rect 19760 20204 19766 20216
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 20993 20207 21051 20213
rect 21542 20204 21548 20256
rect 21600 20204 21606 20256
rect 22097 20247 22155 20253
rect 22097 20213 22109 20247
rect 22143 20244 22155 20247
rect 23842 20244 23848 20256
rect 22143 20216 23848 20244
rect 22143 20213 22155 20216
rect 22097 20207 22155 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 25225 20247 25283 20253
rect 25225 20213 25237 20247
rect 25271 20244 25283 20247
rect 25682 20244 25688 20256
rect 25271 20216 25688 20244
rect 25271 20213 25283 20216
rect 25225 20207 25283 20213
rect 25682 20204 25688 20216
rect 25740 20204 25746 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 1486 20000 1492 20052
rect 1544 20040 1550 20052
rect 1581 20043 1639 20049
rect 1581 20040 1593 20043
rect 1544 20012 1593 20040
rect 1544 20000 1550 20012
rect 1581 20009 1593 20012
rect 1627 20040 1639 20043
rect 4154 20040 4160 20052
rect 1627 20012 4160 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 7469 20043 7527 20049
rect 7469 20009 7481 20043
rect 7515 20040 7527 20043
rect 7650 20040 7656 20052
rect 7515 20012 7656 20040
rect 7515 20009 7527 20012
rect 7469 20003 7527 20009
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8938 20040 8944 20052
rect 8128 20012 8944 20040
rect 5994 19932 6000 19984
rect 6052 19972 6058 19984
rect 8018 19972 8024 19984
rect 6052 19944 8024 19972
rect 6052 19932 6058 19944
rect 8018 19932 8024 19944
rect 8076 19932 8082 19984
rect 2314 19864 2320 19916
rect 2372 19904 2378 19916
rect 2501 19907 2559 19913
rect 2501 19904 2513 19907
rect 2372 19876 2513 19904
rect 2372 19864 2378 19876
rect 2501 19873 2513 19876
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 6362 19904 6368 19916
rect 4019 19876 6368 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 8128 19904 8156 20012
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 9766 20000 9772 20052
rect 9824 20040 9830 20052
rect 10594 20040 10600 20052
rect 9824 20012 10600 20040
rect 9824 20000 9830 20012
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 10888 20012 14933 20040
rect 9306 19932 9312 19984
rect 9364 19972 9370 19984
rect 10778 19972 10784 19984
rect 9364 19944 10784 19972
rect 9364 19932 9370 19944
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 6840 19876 8156 19904
rect 2130 19796 2136 19848
rect 2188 19796 2194 19848
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 4798 19836 4804 19848
rect 4663 19808 4804 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 6840 19845 6868 19876
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 10410 19904 10416 19916
rect 9640 19876 10416 19904
rect 9640 19864 9646 19876
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 10888 19913 10916 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15470 20000 15476 20052
rect 15528 20040 15534 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 15528 20012 17693 20040
rect 15528 20000 15534 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 20441 20043 20499 20049
rect 20441 20040 20453 20043
rect 20220 20012 20453 20040
rect 20220 20000 20226 20012
rect 20441 20009 20453 20012
rect 20487 20009 20499 20043
rect 20441 20003 20499 20009
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 20588 20012 20913 20040
rect 20588 20000 20594 20012
rect 20901 20009 20913 20012
rect 20947 20040 20959 20043
rect 21342 20043 21400 20049
rect 21342 20040 21354 20043
rect 20947 20012 21354 20040
rect 20947 20009 20959 20012
rect 20901 20003 20959 20009
rect 21342 20009 21354 20012
rect 21388 20009 21400 20043
rect 21342 20003 21400 20009
rect 21450 20000 21456 20052
rect 21508 20040 21514 20052
rect 21910 20040 21916 20052
rect 21508 20012 21916 20040
rect 21508 20000 21514 20012
rect 21910 20000 21916 20012
rect 21968 20040 21974 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 21968 20012 22845 20040
rect 21968 20000 21974 20012
rect 22833 20009 22845 20012
rect 22879 20009 22891 20043
rect 22833 20003 22891 20009
rect 24581 20043 24639 20049
rect 24581 20009 24593 20043
rect 24627 20040 24639 20043
rect 25038 20040 25044 20052
rect 24627 20012 25044 20040
rect 24627 20009 24639 20012
rect 24581 20003 24639 20009
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 25590 20000 25596 20052
rect 25648 20040 25654 20052
rect 26050 20040 26056 20052
rect 25648 20012 26056 20040
rect 25648 20000 25654 20012
rect 26050 20000 26056 20012
rect 26108 20000 26114 20052
rect 12912 19944 15516 19972
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 5460 19808 6837 19836
rect 3418 19728 3424 19780
rect 3476 19768 3482 19780
rect 3786 19768 3792 19780
rect 3476 19740 3792 19768
rect 3476 19728 3482 19740
rect 3786 19728 3792 19740
rect 3844 19728 3850 19780
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1673 19703 1731 19709
rect 1673 19700 1685 19703
rect 1452 19672 1685 19700
rect 1452 19660 1458 19672
rect 1673 19669 1685 19672
rect 1719 19669 1731 19703
rect 1673 19663 1731 19669
rect 1946 19660 1952 19712
rect 2004 19700 2010 19712
rect 5460 19700 5488 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 7926 19796 7932 19848
rect 7984 19796 7990 19848
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 9309 19839 9367 19845
rect 8076 19808 8892 19836
rect 8076 19796 8082 19808
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 5994 19768 6000 19780
rect 5776 19740 6000 19768
rect 5776 19728 5782 19740
rect 5994 19728 6000 19740
rect 6052 19728 6058 19780
rect 6546 19728 6552 19780
rect 6604 19728 6610 19780
rect 7006 19728 7012 19780
rect 7064 19768 7070 19780
rect 7282 19768 7288 19780
rect 7064 19740 7288 19768
rect 7064 19728 7070 19740
rect 7282 19728 7288 19740
rect 7340 19728 7346 19780
rect 8864 19768 8892 19808
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9766 19836 9772 19848
rect 9355 19808 9772 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 10980 19836 11008 19867
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 12912 19904 12940 19944
rect 11112 19876 12940 19904
rect 11112 19864 11118 19876
rect 13354 19864 13360 19916
rect 13412 19864 13418 19916
rect 15488 19913 15516 19944
rect 15746 19932 15752 19984
rect 15804 19972 15810 19984
rect 17037 19975 17095 19981
rect 17037 19972 17049 19975
rect 15804 19944 17049 19972
rect 15804 19932 15810 19944
rect 17037 19941 17049 19944
rect 17083 19972 17095 19975
rect 17313 19975 17371 19981
rect 17313 19972 17325 19975
rect 17083 19944 17325 19972
rect 17083 19941 17095 19944
rect 17037 19935 17095 19941
rect 17313 19941 17325 19944
rect 17359 19972 17371 19975
rect 17586 19972 17592 19984
rect 17359 19944 17592 19972
rect 17359 19941 17371 19944
rect 17313 19935 17371 19941
rect 17586 19932 17592 19944
rect 17644 19972 17650 19984
rect 18138 19972 18144 19984
rect 17644 19944 18144 19972
rect 17644 19932 17650 19944
rect 18138 19932 18144 19944
rect 18196 19972 18202 19984
rect 18414 19972 18420 19984
rect 18196 19944 18420 19972
rect 18196 19932 18202 19944
rect 18414 19932 18420 19944
rect 18472 19932 18478 19984
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 15473 19867 15531 19873
rect 15580 19876 18245 19904
rect 10376 19808 11008 19836
rect 10376 19796 10382 19808
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 13909 19839 13967 19845
rect 13909 19836 13921 19839
rect 13464 19808 13921 19836
rect 13464 19780 13492 19808
rect 13909 19805 13921 19808
rect 13955 19836 13967 19839
rect 13998 19836 14004 19848
rect 13955 19808 14004 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 15580 19836 15608 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 18233 19867 18291 19873
rect 18340 19876 19993 19904
rect 14240 19808 15608 19836
rect 14240 19796 14246 19808
rect 16022 19796 16028 19848
rect 16080 19836 16086 19848
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 16080 19808 16129 19836
rect 16080 19796 16086 19808
rect 16117 19805 16129 19808
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16298 19796 16304 19848
rect 16356 19836 16362 19848
rect 18340 19836 18368 19876
rect 19981 19873 19993 19876
rect 20027 19904 20039 19907
rect 20806 19904 20812 19916
rect 20027 19876 20812 19904
rect 20027 19873 20039 19876
rect 19981 19867 20039 19873
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23290 19904 23296 19916
rect 21131 19876 23296 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23658 19864 23664 19916
rect 23716 19904 23722 19916
rect 23753 19907 23811 19913
rect 23753 19904 23765 19907
rect 23716 19876 23765 19904
rect 23716 19864 23722 19876
rect 23753 19873 23765 19876
rect 23799 19873 23811 19907
rect 23753 19867 23811 19873
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19904 23995 19907
rect 24486 19904 24492 19916
rect 23983 19876 24492 19904
rect 23983 19873 23995 19876
rect 23937 19867 23995 19873
rect 24486 19864 24492 19876
rect 24544 19864 24550 19916
rect 24854 19864 24860 19916
rect 24912 19904 24918 19916
rect 25133 19907 25191 19913
rect 25133 19904 25145 19907
rect 24912 19876 25145 19904
rect 24912 19864 24918 19876
rect 25133 19873 25145 19876
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 16356 19808 18368 19836
rect 16356 19796 16362 19808
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 18472 19808 19901 19836
rect 18472 19796 18478 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 24946 19836 24952 19848
rect 19889 19799 19947 19805
rect 19996 19808 21128 19836
rect 22494 19808 24952 19836
rect 9582 19768 9588 19780
rect 8864 19740 9588 19768
rect 9582 19728 9588 19740
rect 9640 19728 9646 19780
rect 9953 19771 10011 19777
rect 9953 19737 9965 19771
rect 9999 19768 10011 19771
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 9999 19740 11897 19768
rect 9999 19737 10011 19740
rect 9953 19731 10011 19737
rect 11885 19737 11897 19740
rect 11931 19737 11943 19771
rect 13446 19768 13452 19780
rect 13110 19740 13452 19768
rect 11885 19731 11943 19737
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 13538 19728 13544 19780
rect 13596 19768 13602 19780
rect 19702 19768 19708 19780
rect 13596 19740 19708 19768
rect 13596 19728 13602 19740
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 2004 19672 5488 19700
rect 2004 19660 2010 19672
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 5810 19700 5816 19712
rect 5592 19672 5816 19700
rect 5592 19660 5598 19672
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 5905 19703 5963 19709
rect 5905 19669 5917 19703
rect 5951 19700 5963 19703
rect 8386 19700 8392 19712
rect 5951 19672 8392 19700
rect 5951 19669 5963 19672
rect 5905 19663 5963 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 8570 19660 8576 19712
rect 8628 19660 8634 19712
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 10413 19703 10471 19709
rect 10413 19700 10425 19703
rect 9824 19672 10425 19700
rect 9824 19660 9830 19672
rect 10413 19669 10425 19672
rect 10459 19669 10471 19703
rect 10413 19663 10471 19669
rect 10594 19660 10600 19712
rect 10652 19700 10658 19712
rect 10781 19703 10839 19709
rect 10781 19700 10793 19703
rect 10652 19672 10793 19700
rect 10652 19660 10658 19672
rect 10781 19669 10793 19672
rect 10827 19669 10839 19703
rect 10781 19663 10839 19669
rect 10870 19660 10876 19712
rect 10928 19700 10934 19712
rect 13170 19700 13176 19712
rect 10928 19672 13176 19700
rect 10928 19660 10934 19672
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13630 19660 13636 19712
rect 13688 19660 13694 19712
rect 14274 19660 14280 19712
rect 14332 19660 14338 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 15160 19672 15301 19700
rect 15160 19660 15166 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 15289 19663 15347 19669
rect 15378 19660 15384 19712
rect 15436 19660 15442 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 16298 19700 16304 19712
rect 15528 19672 16304 19700
rect 15528 19660 15534 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16758 19660 16764 19712
rect 16816 19660 16822 19712
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 17460 19672 17509 19700
rect 17460 19660 17466 19672
rect 17497 19669 17509 19672
rect 17543 19700 17555 19703
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 17543 19672 18061 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18049 19663 18107 19669
rect 18138 19660 18144 19712
rect 18196 19660 18202 19712
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 18693 19703 18751 19709
rect 18693 19700 18705 19703
rect 18564 19672 18705 19700
rect 18564 19660 18570 19672
rect 18693 19669 18705 19672
rect 18739 19669 18751 19703
rect 18693 19663 18751 19669
rect 18874 19660 18880 19712
rect 18932 19700 18938 19712
rect 18969 19703 19027 19709
rect 18969 19700 18981 19703
rect 18932 19672 18981 19700
rect 18932 19660 18938 19672
rect 18969 19669 18981 19672
rect 19015 19669 19027 19703
rect 18969 19663 19027 19669
rect 19426 19660 19432 19712
rect 19484 19660 19490 19712
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 19996 19700 20024 19808
rect 21100 19768 21128 19808
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 21450 19768 21456 19780
rect 21100 19740 21456 19768
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 22738 19728 22744 19780
rect 22796 19768 22802 19780
rect 23661 19771 23719 19777
rect 23661 19768 23673 19771
rect 22796 19740 23673 19768
rect 22796 19728 22802 19740
rect 23661 19737 23673 19740
rect 23707 19768 23719 19771
rect 25406 19768 25412 19780
rect 23707 19740 25412 19768
rect 23707 19737 23719 19740
rect 23661 19731 23719 19737
rect 19843 19672 20024 19700
rect 20717 19703 20775 19709
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20717 19669 20729 19703
rect 20763 19700 20775 19703
rect 20806 19700 20812 19712
rect 20763 19672 20812 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 20806 19660 20812 19672
rect 20864 19660 20870 19712
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21634 19700 21640 19712
rect 21324 19672 21640 19700
rect 21324 19660 21330 19672
rect 21634 19660 21640 19672
rect 21692 19660 21698 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22756 19700 22784 19728
rect 22428 19672 22784 19700
rect 23293 19703 23351 19709
rect 22428 19660 22434 19672
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23566 19700 23572 19712
rect 23339 19672 23572 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23566 19660 23572 19672
rect 23624 19660 23630 19712
rect 24964 19709 24992 19740
rect 25406 19728 25412 19740
rect 25464 19728 25470 19780
rect 24949 19703 25007 19709
rect 24949 19669 24961 19703
rect 24995 19669 25007 19703
rect 24949 19663 25007 19669
rect 25038 19660 25044 19712
rect 25096 19660 25102 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 1486 19456 1492 19508
rect 1544 19456 1550 19508
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4525 19499 4583 19505
rect 4525 19496 4537 19499
rect 4212 19468 4537 19496
rect 4212 19456 4218 19468
rect 4525 19465 4537 19468
rect 4571 19465 4583 19499
rect 9674 19496 9680 19508
rect 4525 19459 4583 19465
rect 4724 19468 9680 19496
rect 4338 19428 4344 19440
rect 1964 19400 4344 19428
rect 1964 19369 1992 19400
rect 4338 19388 4344 19400
rect 4396 19388 4402 19440
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19360 4123 19363
rect 4246 19360 4252 19372
rect 4111 19332 4252 19360
rect 4111 19329 4123 19332
rect 4065 19323 4123 19329
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 4724 19369 4752 19468
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 13814 19496 13820 19508
rect 11664 19468 13820 19496
rect 11664 19456 11670 19468
rect 7466 19388 7472 19440
rect 7524 19388 7530 19440
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 8628 19400 9321 19428
rect 8628 19388 8634 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 10870 19428 10876 19440
rect 10534 19400 10876 19428
rect 9309 19391 9367 19397
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 4798 19320 4804 19372
rect 4856 19320 4862 19372
rect 5810 19320 5816 19372
rect 5868 19360 5874 19372
rect 5997 19363 6055 19369
rect 5997 19360 6009 19363
rect 5868 19332 6009 19360
rect 5868 19320 5874 19332
rect 5997 19329 6009 19332
rect 6043 19329 6055 19363
rect 5997 19323 6055 19329
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 7892 19332 7941 19360
rect 7892 19320 7898 19332
rect 7929 19329 7941 19332
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 12636 19360 12664 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14461 19499 14519 19505
rect 14461 19465 14473 19499
rect 14507 19496 14519 19499
rect 14550 19496 14556 19508
rect 14507 19468 14556 19496
rect 14507 19465 14519 19468
rect 14461 19459 14519 19465
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14792 19468 14933 19496
rect 14792 19456 14798 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 19426 19496 19432 19508
rect 15335 19468 19432 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19659 19468 20453 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 21266 19456 21272 19508
rect 21324 19496 21330 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21324 19468 22017 19496
rect 21324 19456 21330 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22373 19499 22431 19505
rect 22373 19496 22385 19499
rect 22152 19468 22385 19496
rect 22152 19456 22158 19468
rect 22373 19465 22385 19468
rect 22419 19465 22431 19499
rect 22373 19459 22431 19465
rect 22462 19456 22468 19508
rect 22520 19496 22526 19508
rect 23934 19496 23940 19508
rect 22520 19468 23940 19496
rect 22520 19456 22526 19468
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 25041 19499 25099 19505
rect 25041 19465 25053 19499
rect 25087 19496 25099 19499
rect 25222 19496 25228 19508
rect 25087 19468 25228 19496
rect 25087 19465 25099 19468
rect 25041 19459 25099 19465
rect 25222 19456 25228 19468
rect 25280 19496 25286 19508
rect 26510 19496 26516 19508
rect 25280 19468 26516 19496
rect 25280 19456 25286 19468
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 13446 19388 13452 19440
rect 13504 19388 13510 19440
rect 14274 19388 14280 19440
rect 14332 19428 14338 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14332 19400 15393 19428
rect 14332 19388 14338 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 15381 19391 15439 19397
rect 16390 19388 16396 19440
rect 16448 19428 16454 19440
rect 20809 19431 20867 19437
rect 16448 19400 17802 19428
rect 16448 19388 16454 19400
rect 20809 19397 20821 19431
rect 20855 19428 20867 19431
rect 20898 19428 20904 19440
rect 20855 19400 20904 19428
rect 20855 19397 20867 19400
rect 20809 19391 20867 19397
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 24946 19428 24952 19440
rect 24794 19400 24952 19428
rect 24946 19388 24952 19400
rect 25004 19388 25010 19440
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 12636 19332 12725 19360
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 16117 19363 16175 19369
rect 16117 19360 16129 19363
rect 14056 19332 14228 19360
rect 14384 19334 16129 19360
rect 14056 19320 14062 19332
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1728 19264 2237 19292
rect 1728 19252 1734 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 3605 19295 3663 19301
rect 3605 19261 3617 19295
rect 3651 19292 3663 19295
rect 3878 19292 3884 19304
rect 3651 19264 3884 19292
rect 3651 19261 3663 19264
rect 3605 19255 3663 19261
rect 3878 19252 3884 19264
rect 3936 19292 3942 19304
rect 4816 19292 4844 19320
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 3936 19264 4844 19292
rect 5092 19264 5365 19292
rect 3936 19252 3942 19264
rect 5092 19168 5120 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 6917 19295 6975 19301
rect 6917 19261 6929 19295
rect 6963 19292 6975 19295
rect 9398 19292 9404 19304
rect 6963 19264 9404 19292
rect 6963 19261 6975 19264
rect 6917 19255 6975 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 10686 19252 10692 19304
rect 10744 19292 10750 19304
rect 11606 19292 11612 19304
rect 10744 19264 11612 19292
rect 10744 19252 10750 19264
rect 11606 19252 11612 19264
rect 11664 19252 11670 19304
rect 11698 19252 11704 19304
rect 11756 19292 11762 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11756 19264 12265 19292
rect 11756 19252 11762 19264
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 13722 19292 13728 19304
rect 13035 19264 13728 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 8573 19227 8631 19233
rect 8573 19193 8585 19227
rect 8619 19224 8631 19227
rect 8662 19224 8668 19236
rect 8619 19196 8668 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 10962 19184 10968 19236
rect 11020 19224 11026 19236
rect 11020 19196 11468 19224
rect 11020 19184 11026 19196
rect 5074 19116 5080 19168
rect 5132 19116 5138 19168
rect 6549 19159 6607 19165
rect 6549 19125 6561 19159
rect 6595 19156 6607 19159
rect 6822 19156 6828 19168
rect 6595 19128 6828 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 10042 19156 10048 19168
rect 7892 19128 10048 19156
rect 7892 19116 7898 19128
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10468 19128 10793 19156
rect 10468 19116 10474 19128
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 10781 19119 10839 19125
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11057 19159 11115 19165
rect 11057 19156 11069 19159
rect 10928 19128 11069 19156
rect 10928 19116 10934 19128
rect 11057 19125 11069 19128
rect 11103 19125 11115 19159
rect 11057 19119 11115 19125
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11440 19156 11468 19196
rect 13998 19184 14004 19236
rect 14056 19224 14062 19236
rect 14200 19224 14228 19332
rect 14056 19196 14228 19224
rect 14292 19332 16129 19334
rect 14292 19306 14412 19332
rect 16117 19329 16129 19332
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16540 19332 17049 19360
rect 16540 19320 16546 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 17037 19323 17095 19329
rect 18524 19332 19717 19360
rect 14056 19184 14062 19196
rect 13170 19156 13176 19168
rect 11440 19128 13176 19156
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14292 19156 14320 19306
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 17310 19252 17316 19304
rect 17368 19252 17374 19304
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18524 19292 18552 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 22646 19360 22652 19372
rect 19705 19323 19763 19329
rect 20916 19332 22652 19360
rect 17920 19264 18552 19292
rect 18785 19295 18843 19301
rect 17920 19252 17926 19264
rect 18785 19261 18797 19295
rect 18831 19292 18843 19295
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 18831 19264 19901 19292
rect 18831 19261 18843 19264
rect 18785 19255 18843 19261
rect 19889 19261 19901 19264
rect 19935 19292 19947 19295
rect 20162 19292 20168 19304
rect 19935 19264 20168 19292
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 20916 19301 20944 19332
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 24964 19360 24992 19388
rect 25222 19360 25228 19372
rect 24964 19332 25228 19360
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 26234 19360 26240 19372
rect 26108 19332 26240 19360
rect 26108 19320 26114 19332
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 20901 19295 20959 19301
rect 20901 19292 20913 19295
rect 20772 19264 20913 19292
rect 20772 19252 20778 19264
rect 20901 19261 20913 19264
rect 20947 19261 20959 19295
rect 20901 19255 20959 19261
rect 21085 19295 21143 19301
rect 21085 19261 21097 19295
rect 21131 19292 21143 19295
rect 21174 19292 21180 19304
rect 21131 19264 21180 19292
rect 21131 19261 21143 19264
rect 21085 19255 21143 19261
rect 15010 19184 15016 19236
rect 15068 19224 15074 19236
rect 15746 19224 15752 19236
rect 15068 19196 15752 19224
rect 15068 19184 15074 19196
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 16390 19184 16396 19236
rect 16448 19224 16454 19236
rect 17034 19224 17040 19236
rect 16448 19196 17040 19224
rect 16448 19184 16454 19196
rect 17034 19184 17040 19196
rect 17092 19184 17098 19236
rect 21100 19224 21128 19255
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 22278 19252 22284 19304
rect 22336 19292 22342 19304
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22336 19264 22569 19292
rect 22336 19252 22342 19264
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 23658 19292 23664 19304
rect 23615 19264 23664 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 25409 19295 25467 19301
rect 25409 19261 25421 19295
rect 25455 19292 25467 19295
rect 25498 19292 25504 19304
rect 25455 19264 25504 19292
rect 25455 19261 25467 19264
rect 25409 19255 25467 19261
rect 19168 19196 21128 19224
rect 13412 19128 14320 19156
rect 13412 19116 13418 19128
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 14918 19156 14924 19168
rect 14792 19128 14924 19156
rect 14792 19116 14798 19128
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 16206 19156 16212 19168
rect 15436 19128 16212 19156
rect 15436 19116 15442 19128
rect 16206 19116 16212 19128
rect 16264 19156 16270 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16264 19128 16681 19156
rect 16264 19116 16270 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 19168 19156 19196 19196
rect 21542 19184 21548 19236
rect 21600 19224 21606 19236
rect 21726 19224 21732 19236
rect 21600 19196 21732 19224
rect 21600 19184 21606 19196
rect 21726 19184 21732 19196
rect 21784 19224 21790 19236
rect 21784 19196 23428 19224
rect 21784 19184 21790 19196
rect 17000 19128 19196 19156
rect 19245 19159 19303 19165
rect 17000 19116 17006 19128
rect 19245 19125 19257 19159
rect 19291 19156 19303 19159
rect 19334 19156 19340 19168
rect 19291 19128 19340 19156
rect 19291 19125 19303 19128
rect 19245 19119 19303 19125
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 19484 19128 21465 19156
rect 19484 19116 19490 19128
rect 21453 19125 21465 19128
rect 21499 19156 21511 19159
rect 22094 19156 22100 19168
rect 21499 19128 22100 19156
rect 21499 19125 21511 19128
rect 21453 19119 21511 19125
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 22554 19116 22560 19168
rect 22612 19156 22618 19168
rect 22738 19156 22744 19168
rect 22612 19128 22744 19156
rect 22612 19116 22618 19128
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 23400 19156 23428 19196
rect 25424 19156 25452 19255
rect 25498 19252 25504 19264
rect 25556 19252 25562 19304
rect 23400 19128 25452 19156
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 2590 18912 2596 18964
rect 2648 18912 2654 18964
rect 4614 18912 4620 18964
rect 4672 18952 4678 18964
rect 5442 18952 5448 18964
rect 4672 18924 5448 18952
rect 4672 18912 4678 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 7469 18955 7527 18961
rect 7469 18921 7481 18955
rect 7515 18952 7527 18955
rect 8754 18952 8760 18964
rect 7515 18924 8760 18952
rect 7515 18921 7527 18924
rect 7469 18915 7527 18921
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10226 18952 10232 18964
rect 9824 18924 10232 18952
rect 9824 18912 9830 18924
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 11606 18912 11612 18964
rect 11664 18952 11670 18964
rect 13630 18952 13636 18964
rect 11664 18924 13636 18952
rect 11664 18912 11670 18924
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 23382 18952 23388 18964
rect 14608 18924 23388 18952
rect 14608 18912 14614 18924
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 25314 18912 25320 18964
rect 25372 18952 25378 18964
rect 26050 18952 26056 18964
rect 25372 18924 26056 18952
rect 25372 18912 25378 18924
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 1673 18887 1731 18893
rect 1673 18853 1685 18887
rect 1719 18884 1731 18887
rect 2774 18884 2780 18896
rect 1719 18856 2780 18884
rect 1719 18853 1731 18856
rect 1673 18847 1731 18853
rect 2774 18844 2780 18856
rect 2832 18884 2838 18896
rect 3786 18884 3792 18896
rect 2832 18856 3792 18884
rect 2832 18844 2838 18856
rect 3786 18844 3792 18856
rect 3844 18844 3850 18896
rect 12989 18887 13047 18893
rect 12989 18884 13001 18887
rect 8772 18856 13001 18884
rect 8772 18828 8800 18856
rect 12989 18853 13001 18856
rect 13035 18853 13047 18887
rect 15378 18884 15384 18896
rect 12989 18847 13047 18853
rect 13464 18856 15384 18884
rect 3237 18819 3295 18825
rect 3237 18785 3249 18819
rect 3283 18816 3295 18819
rect 3326 18816 3332 18828
rect 3283 18788 3332 18816
rect 3283 18785 3295 18788
rect 3237 18779 3295 18785
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 3970 18776 3976 18828
rect 4028 18776 4034 18828
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18816 4307 18819
rect 5166 18816 5172 18828
rect 4295 18788 5172 18816
rect 4295 18785 4307 18788
rect 4249 18779 4307 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18816 5871 18819
rect 6546 18816 6552 18828
rect 5859 18788 6552 18816
rect 5859 18785 5871 18788
rect 5813 18779 5871 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 8754 18776 8760 18828
rect 8812 18776 8818 18828
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10042 18816 10048 18828
rect 9907 18788 10048 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 11940 18788 12449 18816
rect 11940 18776 11946 18788
rect 12437 18785 12449 18788
rect 12483 18816 12495 18819
rect 13464 18816 13492 18856
rect 12483 18788 13492 18816
rect 13633 18819 13691 18825
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 13633 18785 13645 18819
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 2130 18708 2136 18760
rect 2188 18708 2194 18760
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 6086 18748 6092 18760
rect 2823 18720 6092 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 7929 18751 7987 18757
rect 6880 18720 7880 18748
rect 6880 18708 6886 18720
rect 7558 18680 7564 18692
rect 1964 18652 7564 18680
rect 1486 18572 1492 18624
rect 1544 18572 1550 18624
rect 1964 18621 1992 18652
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 7852 18680 7880 18720
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 10318 18748 10324 18760
rect 7975 18720 10324 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 10413 18751 10471 18757
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11330 18748 11336 18760
rect 10459 18720 11336 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 13648 18692 13676 18779
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14274 18816 14280 18828
rect 13872 18788 14280 18816
rect 13872 18776 13878 18788
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14752 18825 14780 18856
rect 15378 18844 15384 18856
rect 15436 18844 15442 18896
rect 15470 18844 15476 18896
rect 15528 18844 15534 18896
rect 17218 18844 17224 18896
rect 17276 18844 17282 18896
rect 19426 18884 19432 18896
rect 18892 18856 19432 18884
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18785 14795 18819
rect 14737 18779 14795 18785
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18816 14979 18819
rect 15488 18816 15516 18844
rect 14967 18788 15516 18816
rect 15749 18819 15807 18825
rect 14967 18785 14979 18788
rect 14921 18779 14979 18785
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 16758 18816 16764 18828
rect 15795 18788 16764 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 17586 18776 17592 18828
rect 17644 18816 17650 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 17644 18788 18613 18816
rect 17644 18776 17650 18788
rect 18601 18785 18613 18788
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 13924 18720 14504 18748
rect 11054 18680 11060 18692
rect 7852 18652 11060 18680
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 13262 18680 13268 18692
rect 11624 18652 13268 18680
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18581 2007 18615
rect 1949 18575 2007 18581
rect 3050 18572 3056 18624
rect 3108 18612 3114 18624
rect 3602 18612 3608 18624
rect 3108 18584 3608 18612
rect 3108 18572 3114 18584
rect 3602 18572 3608 18584
rect 3660 18572 3666 18624
rect 5166 18572 5172 18624
rect 5224 18572 5230 18624
rect 6362 18572 6368 18624
rect 6420 18572 6426 18624
rect 6822 18572 6828 18624
rect 6880 18612 6886 18624
rect 7742 18612 7748 18624
rect 6880 18584 7748 18612
rect 6880 18572 6886 18584
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 8570 18572 8576 18624
rect 8628 18572 8634 18624
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 8720 18584 9229 18612
rect 8720 18572 8726 18584
rect 9217 18581 9229 18584
rect 9263 18581 9275 18615
rect 9217 18575 9275 18581
rect 9582 18572 9588 18624
rect 9640 18572 9646 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 11624 18612 11652 18652
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 13446 18640 13452 18692
rect 13504 18640 13510 18692
rect 13630 18640 13636 18692
rect 13688 18640 13694 18692
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 13924 18680 13952 18720
rect 13780 18652 13952 18680
rect 13780 18640 13786 18652
rect 9723 18584 11652 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 12713 18615 12771 18621
rect 12713 18581 12725 18615
rect 12759 18612 12771 18615
rect 12894 18612 12900 18624
rect 12759 18584 12900 18612
rect 12759 18581 12771 18584
rect 12713 18575 12771 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14476 18612 14504 18720
rect 15010 18708 15016 18760
rect 15068 18748 15074 18760
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 15068 18720 15485 18748
rect 15068 18708 15074 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17092 18720 17693 18748
rect 17092 18708 17098 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 17920 18720 18429 18748
rect 17920 18708 17926 18720
rect 18417 18717 18429 18720
rect 18463 18748 18475 18751
rect 18892 18748 18920 18856
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 19610 18844 19616 18896
rect 19668 18884 19674 18896
rect 19705 18887 19763 18893
rect 19705 18884 19717 18887
rect 19668 18856 19717 18884
rect 19668 18844 19674 18856
rect 19705 18853 19717 18856
rect 19751 18853 19763 18887
rect 19705 18847 19763 18853
rect 22557 18887 22615 18893
rect 22557 18853 22569 18887
rect 22603 18884 22615 18887
rect 24581 18887 24639 18893
rect 22603 18856 24532 18884
rect 22603 18853 22615 18856
rect 22557 18847 22615 18853
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19392 18788 22094 18816
rect 19392 18776 19398 18788
rect 18463 18720 18920 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 19300 18720 20361 18748
rect 19300 18708 19306 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 21726 18708 21732 18760
rect 21784 18708 21790 18760
rect 22066 18748 22094 18788
rect 22738 18776 22744 18828
rect 22796 18816 22802 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22796 18788 23121 18816
rect 22796 18776 22802 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23845 18751 23903 18757
rect 23845 18748 23857 18751
rect 22066 18720 23857 18748
rect 23845 18717 23857 18720
rect 23891 18717 23903 18751
rect 24504 18748 24532 18856
rect 24581 18853 24593 18887
rect 24627 18884 24639 18887
rect 25498 18884 25504 18896
rect 24627 18856 25504 18884
rect 24627 18853 24639 18856
rect 24581 18847 24639 18853
rect 25498 18844 25504 18856
rect 25556 18844 25562 18896
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18816 25283 18819
rect 25682 18816 25688 18828
rect 25271 18788 25688 18816
rect 25271 18785 25283 18788
rect 25225 18779 25283 18785
rect 25682 18776 25688 18788
rect 25740 18776 25746 18828
rect 24504 18720 25360 18748
rect 23845 18711 23903 18717
rect 16206 18640 16212 18692
rect 16264 18640 16270 18692
rect 17770 18640 17776 18692
rect 17828 18680 17834 18692
rect 18509 18683 18567 18689
rect 17828 18652 18460 18680
rect 17828 18640 17834 18652
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 14476 18584 14657 18612
rect 14645 18581 14657 18584
rect 14691 18612 14703 18615
rect 15746 18612 15752 18624
rect 14691 18584 15752 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 15746 18572 15752 18584
rect 15804 18612 15810 18624
rect 17034 18612 17040 18624
rect 15804 18584 17040 18612
rect 15804 18572 15810 18584
rect 17034 18572 17040 18584
rect 17092 18612 17098 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17092 18584 17509 18612
rect 17092 18572 17098 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 18049 18615 18107 18621
rect 18049 18581 18061 18615
rect 18095 18612 18107 18615
rect 18322 18612 18328 18624
rect 18095 18584 18328 18612
rect 18095 18581 18107 18584
rect 18049 18575 18107 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18432 18612 18460 18652
rect 18509 18649 18521 18683
rect 18555 18680 18567 18683
rect 19150 18680 19156 18692
rect 18555 18652 19156 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 19150 18640 19156 18652
rect 19208 18640 19214 18692
rect 19426 18640 19432 18692
rect 19484 18680 19490 18692
rect 19521 18683 19579 18689
rect 19521 18680 19533 18683
rect 19484 18652 19533 18680
rect 19484 18640 19490 18652
rect 19521 18649 19533 18652
rect 19567 18649 19579 18683
rect 19521 18643 19579 18649
rect 20622 18640 20628 18692
rect 20680 18640 20686 18692
rect 23014 18640 23020 18692
rect 23072 18680 23078 18692
rect 24026 18680 24032 18692
rect 23072 18652 24032 18680
rect 23072 18640 23078 18652
rect 24026 18640 24032 18652
rect 24084 18640 24090 18692
rect 25041 18683 25099 18689
rect 25041 18649 25053 18683
rect 25087 18680 25099 18683
rect 25130 18680 25136 18692
rect 25087 18652 25136 18680
rect 25087 18649 25099 18652
rect 25041 18643 25099 18649
rect 25130 18640 25136 18652
rect 25188 18640 25194 18692
rect 25332 18624 25360 18720
rect 20073 18615 20131 18621
rect 20073 18612 20085 18615
rect 18432 18584 20085 18612
rect 20073 18581 20085 18584
rect 20119 18612 20131 18615
rect 20530 18612 20536 18624
rect 20119 18584 20536 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 22097 18615 22155 18621
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22370 18612 22376 18624
rect 22143 18584 22376 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22646 18572 22652 18624
rect 22704 18612 22710 18624
rect 22925 18615 22983 18621
rect 22925 18612 22937 18615
rect 22704 18584 22937 18612
rect 22704 18572 22710 18584
rect 22925 18581 22937 18584
rect 22971 18612 22983 18615
rect 23382 18612 23388 18624
rect 22971 18584 23388 18612
rect 22971 18581 22983 18584
rect 22925 18575 22983 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23716 18584 23949 18612
rect 23716 18572 23722 18584
rect 23937 18581 23949 18584
rect 23983 18581 23995 18615
rect 23937 18575 23995 18581
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 25314 18572 25320 18624
rect 25372 18572 25378 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 8662 18408 8668 18420
rect 3620 18380 8668 18408
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 2777 18275 2835 18281
rect 2777 18272 2789 18275
rect 1627 18244 2789 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2777 18241 2789 18244
rect 2823 18272 2835 18275
rect 3050 18272 3056 18284
rect 2823 18244 3056 18272
rect 2823 18241 2835 18244
rect 2777 18235 2835 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3620 18281 3648 18380
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 9364 18380 10701 18408
rect 9364 18368 9370 18380
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 10689 18371 10747 18377
rect 5626 18340 5632 18352
rect 4724 18312 5632 18340
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 4338 18272 4344 18284
rect 4295 18244 4344 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 4338 18232 4344 18244
rect 4396 18232 4402 18284
rect 4724 18281 4752 18312
rect 5626 18300 5632 18312
rect 5684 18340 5690 18352
rect 5813 18343 5871 18349
rect 5813 18340 5825 18343
rect 5684 18312 5825 18340
rect 5684 18300 5690 18312
rect 5813 18309 5825 18312
rect 5859 18309 5871 18343
rect 5813 18303 5871 18309
rect 6178 18300 6184 18352
rect 6236 18300 6242 18352
rect 8294 18340 8300 18352
rect 6380 18312 8300 18340
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18272 5043 18275
rect 6380 18272 6408 18312
rect 8294 18300 8300 18312
rect 8352 18300 8358 18352
rect 8570 18300 8576 18352
rect 8628 18340 8634 18352
rect 9217 18343 9275 18349
rect 9217 18340 9229 18343
rect 8628 18312 9229 18340
rect 8628 18300 8634 18312
rect 9217 18309 9229 18312
rect 9263 18309 9275 18343
rect 10704 18340 10732 18371
rect 10870 18368 10876 18420
rect 10928 18408 10934 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10928 18380 11069 18408
rect 10928 18368 10934 18380
rect 11057 18377 11069 18380
rect 11103 18408 11115 18411
rect 11241 18411 11299 18417
rect 11241 18408 11253 18411
rect 11103 18380 11253 18408
rect 11103 18377 11115 18380
rect 11057 18371 11115 18377
rect 11241 18377 11253 18380
rect 11287 18377 11299 18411
rect 11241 18371 11299 18377
rect 11330 18368 11336 18420
rect 11388 18408 11394 18420
rect 13538 18408 13544 18420
rect 11388 18380 13544 18408
rect 11388 18368 11394 18380
rect 13004 18349 13032 18380
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 13998 18408 14004 18420
rect 13872 18380 14004 18408
rect 13872 18368 13878 18380
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 14274 18368 14280 18420
rect 14332 18408 14338 18420
rect 14918 18408 14924 18420
rect 14332 18380 14924 18408
rect 14332 18368 14338 18380
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 15120 18380 15209 18408
rect 12989 18343 13047 18349
rect 10704 18312 12296 18340
rect 9217 18303 9275 18309
rect 5031 18244 6408 18272
rect 6457 18275 6515 18281
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 6457 18241 6469 18275
rect 6503 18272 6515 18275
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6503 18244 6745 18272
rect 6503 18241 6515 18244
rect 6457 18235 6515 18241
rect 6733 18241 6745 18244
rect 6779 18272 6791 18275
rect 7374 18272 7380 18284
rect 6779 18244 7380 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7837 18275 7895 18281
rect 7837 18241 7849 18275
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 1854 18164 1860 18216
rect 1912 18164 1918 18216
rect 2961 18207 3019 18213
rect 2961 18173 2973 18207
rect 3007 18204 3019 18207
rect 7650 18204 7656 18216
rect 3007 18176 7656 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7852 18204 7880 18235
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 10870 18272 10876 18284
rect 10350 18244 10876 18272
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 12158 18232 12164 18284
rect 12216 18232 12222 18284
rect 12268 18272 12296 18312
rect 12989 18309 13001 18343
rect 13035 18309 13047 18343
rect 12989 18303 13047 18309
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 15120 18340 15148 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15378 18408 15384 18420
rect 15344 18380 15384 18408
rect 15344 18368 15350 18380
rect 15378 18368 15384 18380
rect 15436 18408 15442 18420
rect 15436 18380 15700 18408
rect 15436 18368 15442 18380
rect 15672 18349 15700 18380
rect 17310 18368 17316 18420
rect 17368 18408 17374 18420
rect 17368 18380 23244 18408
rect 17368 18368 17374 18380
rect 15657 18343 15715 18349
rect 13320 18312 15148 18340
rect 15396 18312 15608 18340
rect 13320 18300 13326 18312
rect 15396 18284 15424 18312
rect 13538 18272 13544 18284
rect 12268 18244 13544 18272
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 15378 18232 15384 18284
rect 15436 18232 15442 18284
rect 15580 18281 15608 18312
rect 15657 18309 15669 18343
rect 15703 18309 15715 18343
rect 15657 18303 15715 18309
rect 16209 18343 16267 18349
rect 16209 18309 16221 18343
rect 16255 18340 16267 18343
rect 16574 18340 16580 18352
rect 16255 18312 16580 18340
rect 16255 18309 16267 18312
rect 16209 18303 16267 18309
rect 16574 18300 16580 18312
rect 16632 18340 16638 18352
rect 18417 18343 18475 18349
rect 16632 18312 17908 18340
rect 16632 18300 16638 18312
rect 15565 18275 15623 18281
rect 15565 18241 15577 18275
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17770 18272 17776 18284
rect 17359 18244 17776 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 9950 18204 9956 18216
rect 7852 18176 9956 18204
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 12066 18204 12072 18216
rect 10468 18176 12072 18204
rect 10468 18164 10474 18176
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 3145 18139 3203 18145
rect 3145 18105 3157 18139
rect 3191 18136 3203 18139
rect 4065 18139 4123 18145
rect 3191 18108 4016 18136
rect 3191 18105 3203 18108
rect 3145 18099 3203 18105
rect 3418 18028 3424 18080
rect 3476 18028 3482 18080
rect 3988 18068 4016 18108
rect 4065 18105 4077 18139
rect 4111 18136 4123 18139
rect 8202 18136 8208 18148
rect 4111 18108 8208 18136
rect 4111 18105 4123 18108
rect 4065 18099 4123 18105
rect 8202 18096 8208 18108
rect 8260 18096 8266 18148
rect 12268 18136 12296 18167
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 12710 18204 12716 18216
rect 12492 18176 12716 18204
rect 12492 18164 12498 18176
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13354 18204 13360 18216
rect 12952 18176 13360 18204
rect 12952 18164 12958 18176
rect 13354 18164 13360 18176
rect 13412 18204 13418 18216
rect 13412 18176 15332 18204
rect 13412 18164 13418 18176
rect 15010 18136 15016 18148
rect 12268 18108 15016 18136
rect 15010 18096 15016 18108
rect 15068 18096 15074 18148
rect 15304 18136 15332 18176
rect 15470 18164 15476 18216
rect 15528 18164 15534 18216
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 17497 18167 17555 18173
rect 15488 18136 15516 18164
rect 15304 18108 15516 18136
rect 4890 18068 4896 18080
rect 3988 18040 4896 18068
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6638 18068 6644 18080
rect 6328 18040 6644 18068
rect 6328 18028 6334 18040
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7377 18071 7435 18077
rect 7377 18037 7389 18071
rect 7423 18068 7435 18071
rect 7650 18068 7656 18080
rect 7423 18040 7656 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 8481 18071 8539 18077
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 9950 18068 9956 18080
rect 8527 18040 9956 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11388 18040 11805 18068
rect 11388 18028 11394 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 15102 18068 15108 18080
rect 12768 18040 15108 18068
rect 12768 18028 12774 18040
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15764 18068 15792 18167
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 17512 18136 17540 18167
rect 16356 18108 17540 18136
rect 17880 18136 17908 18312
rect 18417 18309 18429 18343
rect 18463 18340 18475 18343
rect 20809 18343 20867 18349
rect 20809 18340 20821 18343
rect 18463 18312 20821 18340
rect 18463 18309 18475 18312
rect 18417 18303 18475 18309
rect 20809 18309 20821 18312
rect 20855 18340 20867 18343
rect 21453 18343 21511 18349
rect 21453 18340 21465 18343
rect 20855 18312 21465 18340
rect 20855 18309 20867 18312
rect 20809 18303 20867 18309
rect 21453 18309 21465 18312
rect 21499 18340 21511 18343
rect 21542 18340 21548 18352
rect 21499 18312 21548 18340
rect 21499 18309 21511 18312
rect 21453 18303 21511 18309
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 22002 18300 22008 18352
rect 22060 18300 22066 18352
rect 23216 18340 23244 18380
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 25317 18411 25375 18417
rect 25317 18408 25329 18411
rect 23440 18380 25329 18408
rect 23440 18368 23446 18380
rect 25317 18377 25329 18380
rect 25363 18408 25375 18411
rect 25406 18408 25412 18420
rect 25363 18380 25412 18408
rect 25363 18377 25375 18380
rect 25317 18371 25375 18377
rect 25406 18368 25412 18380
rect 25464 18408 25470 18420
rect 25774 18408 25780 18420
rect 25464 18380 25780 18408
rect 25464 18368 25470 18380
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 24857 18343 24915 18349
rect 24857 18340 24869 18343
rect 23216 18312 24869 18340
rect 24857 18309 24869 18312
rect 24903 18309 24915 18343
rect 24857 18303 24915 18309
rect 25222 18300 25228 18352
rect 25280 18300 25286 18352
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 18748 18244 19625 18272
rect 18748 18232 18754 18244
rect 19613 18241 19625 18244
rect 19659 18272 19671 18275
rect 20714 18272 20720 18284
rect 19659 18244 20720 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21174 18232 21180 18284
rect 21232 18272 21238 18284
rect 24213 18275 24271 18281
rect 24213 18272 24225 18275
rect 21232 18244 24225 18272
rect 21232 18232 21238 18244
rect 24213 18241 24225 18244
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 18506 18164 18512 18216
rect 18564 18164 18570 18216
rect 18598 18164 18604 18216
rect 18656 18164 18662 18216
rect 18874 18164 18880 18216
rect 18932 18204 18938 18216
rect 19705 18207 19763 18213
rect 19705 18204 19717 18207
rect 18932 18176 19717 18204
rect 18932 18164 18938 18176
rect 19705 18173 19717 18176
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 19886 18164 19892 18216
rect 19944 18164 19950 18216
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21085 18207 21143 18213
rect 21085 18173 21097 18207
rect 21131 18204 21143 18207
rect 24026 18204 24032 18216
rect 21131 18176 24032 18204
rect 21131 18173 21143 18176
rect 21085 18167 21143 18173
rect 19058 18136 19064 18148
rect 17880 18108 19064 18136
rect 16356 18096 16362 18108
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 20806 18136 20812 18148
rect 19392 18108 20812 18136
rect 19392 18096 19398 18108
rect 20806 18096 20812 18108
rect 20864 18136 20870 18148
rect 20916 18136 20944 18167
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 20864 18108 20944 18136
rect 20864 18096 20870 18108
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 26694 18136 26700 18148
rect 21968 18108 26700 18136
rect 21968 18096 21974 18108
rect 26694 18096 26700 18108
rect 26752 18096 26758 18148
rect 15528 18040 15792 18068
rect 15528 18028 15534 18040
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16264 18040 16405 18068
rect 16264 18028 16270 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16393 18031 16451 18037
rect 16758 18028 16764 18080
rect 16816 18068 16822 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16816 18040 16865 18068
rect 16816 18028 16822 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 17494 18028 17500 18080
rect 17552 18068 17558 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17552 18040 18061 18068
rect 17552 18028 17558 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 19245 18071 19303 18077
rect 19245 18037 19257 18071
rect 19291 18068 19303 18071
rect 19794 18068 19800 18080
rect 19291 18040 19800 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 21082 18068 21088 18080
rect 20487 18040 21088 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 22554 18068 22560 18080
rect 22244 18040 22560 18068
rect 22244 18028 22250 18040
rect 22554 18028 22560 18040
rect 22612 18068 22618 18080
rect 23290 18068 23296 18080
rect 22612 18040 23296 18068
rect 22612 18028 22618 18040
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 6914 17864 6920 17876
rect 1872 17836 6920 17864
rect 1872 17737 1900 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 12618 17864 12624 17876
rect 8864 17836 12624 17864
rect 3237 17799 3295 17805
rect 3237 17765 3249 17799
rect 3283 17796 3295 17799
rect 5902 17796 5908 17808
rect 3283 17768 5908 17796
rect 3283 17765 3295 17768
rect 3237 17759 3295 17765
rect 5902 17756 5908 17768
rect 5960 17756 5966 17808
rect 5997 17799 6055 17805
rect 5997 17765 6009 17799
rect 6043 17796 6055 17799
rect 8662 17796 8668 17808
rect 6043 17768 8668 17796
rect 6043 17765 6055 17768
rect 5997 17759 6055 17765
rect 8662 17756 8668 17768
rect 8720 17756 8726 17808
rect 1857 17731 1915 17737
rect 1857 17697 1869 17731
rect 1903 17697 1915 17731
rect 4154 17728 4160 17740
rect 1857 17691 1915 17697
rect 2746 17700 4160 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 2746 17660 2774 17700
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 4430 17688 4436 17740
rect 4488 17728 4494 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4488 17700 4813 17728
rect 4488 17688 4494 17700
rect 4801 17697 4813 17700
rect 4847 17697 4859 17731
rect 6730 17728 6736 17740
rect 4801 17691 4859 17697
rect 5644 17700 6736 17728
rect 1627 17632 2774 17660
rect 3421 17663 3479 17669
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3881 17663 3939 17669
rect 3881 17660 3893 17663
rect 3467 17632 3893 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3881 17629 3893 17632
rect 3927 17660 3939 17663
rect 3970 17660 3976 17672
rect 3927 17632 3976 17660
rect 3927 17629 3939 17632
rect 3881 17623 3939 17629
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 4525 17663 4583 17669
rect 4525 17629 4537 17663
rect 4571 17660 4583 17663
rect 5644 17660 5672 17700
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 8864 17728 8892 17836
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 13504 17836 17141 17864
rect 13504 17824 13510 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 23382 17864 23388 17876
rect 17129 17827 17187 17833
rect 17236 17836 23388 17864
rect 11514 17756 11520 17808
rect 11572 17756 11578 17808
rect 11606 17756 11612 17808
rect 11664 17796 11670 17808
rect 13725 17799 13783 17805
rect 11664 17768 12112 17796
rect 11664 17756 11670 17768
rect 7944 17700 8892 17728
rect 9769 17731 9827 17737
rect 4571 17632 5672 17660
rect 5721 17663 5779 17669
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 5721 17629 5733 17663
rect 5767 17660 5779 17663
rect 6178 17660 6184 17672
rect 5767 17632 6184 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6825 17663 6883 17669
rect 6825 17660 6837 17663
rect 6328 17632 6837 17660
rect 6328 17620 6334 17632
rect 6825 17629 6837 17632
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 7466 17620 7472 17672
rect 7524 17620 7530 17672
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 7834 17660 7840 17672
rect 7708 17632 7840 17660
rect 7708 17620 7714 17632
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 7944 17669 7972 17700
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 11698 17728 11704 17740
rect 9815 17700 11704 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9784 17660 9812 17691
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11756 17700 11989 17728
rect 11756 17688 11762 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 12084 17728 12112 17768
rect 13725 17765 13737 17799
rect 13771 17796 13783 17799
rect 14458 17796 14464 17808
rect 13771 17768 14464 17796
rect 13771 17765 13783 17768
rect 13725 17759 13783 17765
rect 14458 17756 14464 17768
rect 14516 17796 14522 17808
rect 14516 17768 15056 17796
rect 14516 17756 14522 17768
rect 14185 17731 14243 17737
rect 12084 17700 13492 17728
rect 11977 17691 12035 17697
rect 8996 17632 9812 17660
rect 13464 17660 13492 17700
rect 14185 17697 14197 17731
rect 14231 17728 14243 17731
rect 14274 17728 14280 17740
rect 14231 17700 14280 17728
rect 14231 17697 14243 17700
rect 14185 17691 14243 17697
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 14918 17688 14924 17740
rect 14976 17688 14982 17740
rect 15028 17728 15056 17768
rect 16298 17756 16304 17808
rect 16356 17756 16362 17808
rect 16482 17756 16488 17808
rect 16540 17796 16546 17808
rect 17236 17796 17264 17836
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 16540 17768 17264 17796
rect 16540 17756 16546 17768
rect 17310 17756 17316 17808
rect 17368 17796 17374 17808
rect 18601 17799 18659 17805
rect 18601 17796 18613 17799
rect 17368 17768 18613 17796
rect 17368 17756 17374 17768
rect 18601 17765 18613 17768
rect 18647 17765 18659 17799
rect 18601 17759 18659 17765
rect 22465 17799 22523 17805
rect 22465 17765 22477 17799
rect 22511 17765 22523 17799
rect 22465 17759 22523 17765
rect 16316 17728 16344 17756
rect 15028 17700 16344 17728
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16632 17700 17693 17728
rect 16632 17688 16638 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 19242 17728 19248 17740
rect 18380 17700 19248 17728
rect 18380 17688 18386 17700
rect 19242 17688 19248 17700
rect 19300 17688 19306 17740
rect 20070 17688 20076 17740
rect 20128 17688 20134 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 22186 17728 22192 17740
rect 20763 17700 22192 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 22480 17672 22508 17759
rect 22922 17756 22928 17808
rect 22980 17796 22986 17808
rect 23109 17799 23167 17805
rect 23109 17796 23121 17799
rect 22980 17768 23121 17796
rect 22980 17756 22986 17768
rect 23109 17765 23121 17768
rect 23155 17765 23167 17799
rect 23109 17759 23167 17765
rect 23124 17728 23152 17759
rect 23474 17756 23480 17808
rect 23532 17796 23538 17808
rect 23532 17768 23888 17796
rect 23532 17756 23538 17768
rect 23124 17700 23704 17728
rect 14550 17660 14556 17672
rect 13464 17632 14556 17660
rect 8996 17620 9002 17632
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 16666 17620 16672 17672
rect 16724 17660 16730 17672
rect 17497 17663 17555 17669
rect 17497 17660 17509 17663
rect 16724 17632 17509 17660
rect 16724 17620 16730 17632
rect 17497 17629 17509 17632
rect 17543 17629 17555 17663
rect 17497 17623 17555 17629
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 17828 17632 19901 17660
rect 17828 17620 17834 17632
rect 19889 17629 19901 17632
rect 19935 17660 19947 17663
rect 20622 17660 20628 17672
rect 19935 17632 20628 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 23474 17660 23480 17672
rect 22879 17632 23480 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 23676 17669 23704 17700
rect 23750 17688 23756 17740
rect 23808 17688 23814 17740
rect 23860 17737 23888 17768
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17697 23903 17731
rect 23845 17691 23903 17697
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 2869 17595 2927 17601
rect 2869 17592 2881 17595
rect 1544 17564 2881 17592
rect 1544 17552 1550 17564
rect 2869 17561 2881 17564
rect 2915 17592 2927 17595
rect 5442 17592 5448 17604
rect 2915 17564 5448 17592
rect 2915 17561 2927 17564
rect 2869 17555 2927 17561
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 8478 17592 8484 17604
rect 6656 17564 8484 17592
rect 2774 17484 2780 17536
rect 2832 17484 2838 17536
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 3973 17527 4031 17533
rect 3973 17524 3985 17527
rect 3936 17496 3985 17524
rect 3936 17484 3942 17496
rect 3973 17493 3985 17496
rect 4019 17524 4031 17527
rect 4154 17524 4160 17536
rect 4019 17496 4160 17524
rect 4019 17493 4031 17496
rect 3973 17487 4031 17493
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 5626 17524 5632 17536
rect 4304 17496 5632 17524
rect 4304 17484 4310 17496
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 6656 17533 6684 17564
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 8573 17595 8631 17601
rect 8573 17561 8585 17595
rect 8619 17592 8631 17595
rect 8619 17564 9904 17592
rect 8619 17561 8631 17564
rect 8573 17555 8631 17561
rect 6641 17527 6699 17533
rect 6641 17493 6653 17527
rect 6687 17493 6699 17527
rect 6641 17487 6699 17493
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17524 7343 17527
rect 7834 17524 7840 17536
rect 7331 17496 7840 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 7834 17484 7840 17496
rect 7892 17484 7898 17536
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17524 9183 17527
rect 9582 17524 9588 17536
rect 9171 17496 9588 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9876 17524 9904 17564
rect 9950 17552 9956 17604
rect 10008 17592 10014 17604
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 10008 17564 10057 17592
rect 10008 17552 10014 17564
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 10778 17552 10784 17604
rect 10836 17552 10842 17604
rect 12253 17595 12311 17601
rect 12253 17592 12265 17595
rect 11348 17564 12265 17592
rect 11348 17524 11376 17564
rect 12253 17561 12265 17564
rect 12299 17561 12311 17595
rect 12253 17555 12311 17561
rect 12986 17552 12992 17604
rect 13044 17552 13050 17604
rect 15194 17552 15200 17604
rect 15252 17552 15258 17604
rect 15304 17564 15686 17592
rect 9876 17496 11376 17524
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 12526 17524 12532 17536
rect 11480 17496 12532 17524
rect 11480 17484 11486 17496
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 14734 17524 14740 17536
rect 14056 17496 14740 17524
rect 14056 17484 14062 17496
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 15010 17484 15016 17536
rect 15068 17524 15074 17536
rect 15304 17524 15332 17564
rect 15068 17496 15332 17524
rect 15580 17524 15608 17564
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 18417 17595 18475 17601
rect 18417 17592 18429 17595
rect 16540 17564 18429 17592
rect 16540 17552 16546 17564
rect 18417 17561 18429 17564
rect 18463 17561 18475 17595
rect 18417 17555 18475 17561
rect 18966 17552 18972 17604
rect 19024 17592 19030 17604
rect 19797 17595 19855 17601
rect 19797 17592 19809 17595
rect 19024 17564 19809 17592
rect 19024 17552 19030 17564
rect 19797 17561 19809 17564
rect 19843 17561 19855 17595
rect 19797 17555 19855 17561
rect 16206 17524 16212 17536
rect 15580 17496 16212 17524
rect 15068 17484 15074 17496
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16669 17527 16727 17533
rect 16669 17493 16681 17527
rect 16715 17524 16727 17527
rect 16942 17524 16948 17536
rect 16715 17496 16948 17524
rect 16715 17493 16727 17496
rect 16669 17487 16727 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 17034 17484 17040 17536
rect 17092 17524 17098 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 17092 17496 17601 17524
rect 17092 17484 17098 17496
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 17589 17487 17647 17493
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 18877 17527 18935 17533
rect 18877 17524 18889 17527
rect 17736 17496 18889 17524
rect 17736 17484 17742 17496
rect 18877 17493 18889 17496
rect 18923 17493 18935 17527
rect 18877 17487 18935 17493
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19610 17524 19616 17536
rect 19475 17496 19616 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 19812 17524 19840 17555
rect 20990 17552 20996 17604
rect 21048 17552 21054 17604
rect 21726 17552 21732 17604
rect 21784 17552 21790 17604
rect 22922 17552 22928 17604
rect 22980 17592 22986 17604
rect 25225 17595 25283 17601
rect 25225 17592 25237 17595
rect 22980 17564 25237 17592
rect 22980 17552 22986 17564
rect 25225 17561 25237 17564
rect 25271 17561 25283 17595
rect 25225 17555 25283 17561
rect 22646 17524 22652 17536
rect 19812 17496 22652 17524
rect 22646 17484 22652 17496
rect 22704 17524 22710 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22704 17496 23029 17524
rect 22704 17484 22710 17496
rect 23017 17493 23029 17496
rect 23063 17524 23075 17527
rect 23198 17524 23204 17536
rect 23063 17496 23204 17524
rect 23063 17493 23075 17496
rect 23017 17487 23075 17493
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23290 17484 23296 17536
rect 23348 17484 23354 17536
rect 23474 17484 23480 17536
rect 23532 17524 23538 17536
rect 24210 17524 24216 17536
rect 23532 17496 24216 17524
rect 23532 17484 23538 17496
rect 24210 17484 24216 17496
rect 24268 17484 24274 17536
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 2130 17320 2136 17332
rect 1719 17292 2136 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 3467 17323 3525 17329
rect 3467 17289 3479 17323
rect 3513 17320 3525 17323
rect 7006 17320 7012 17332
rect 3513 17292 7012 17320
rect 3513 17289 3525 17292
rect 3467 17283 3525 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7190 17320 7196 17332
rect 7116 17292 7196 17320
rect 1489 17255 1547 17261
rect 1489 17221 1501 17255
rect 1535 17252 1547 17255
rect 1762 17252 1768 17264
rect 1535 17224 1768 17252
rect 1535 17221 1547 17224
rect 1489 17215 1547 17221
rect 1762 17212 1768 17224
rect 1820 17212 1826 17264
rect 4246 17212 4252 17264
rect 4304 17252 4310 17264
rect 6914 17252 6920 17264
rect 4304 17224 6920 17252
rect 4304 17212 4310 17224
rect 6914 17212 6920 17224
rect 6972 17212 6978 17264
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 2096 17156 2237 17184
rect 2096 17144 2102 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17184 3295 17187
rect 4614 17184 4620 17196
rect 3283 17156 4620 17184
rect 3283 17153 3295 17156
rect 3237 17147 3295 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4982 17184 4988 17196
rect 4847 17156 4988 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 7116 17184 7144 17292
rect 7190 17280 7196 17292
rect 7248 17320 7254 17332
rect 7653 17323 7711 17329
rect 7653 17320 7665 17323
rect 7248 17292 7665 17320
rect 7248 17280 7254 17292
rect 7653 17289 7665 17292
rect 7699 17289 7711 17323
rect 7653 17283 7711 17289
rect 8757 17323 8815 17329
rect 8757 17289 8769 17323
rect 8803 17320 8815 17323
rect 8803 17292 12020 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 10778 17212 10784 17264
rect 10836 17252 10842 17264
rect 11422 17252 11428 17264
rect 10836 17224 11428 17252
rect 10836 17212 10842 17224
rect 11422 17212 11428 17224
rect 11480 17212 11486 17264
rect 11992 17261 12020 17292
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 13449 17323 13507 17329
rect 13449 17320 13461 17323
rect 12676 17292 13461 17320
rect 12676 17280 12682 17292
rect 13449 17289 13461 17292
rect 13495 17289 13507 17323
rect 13449 17283 13507 17289
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 14090 17320 14096 17332
rect 13780 17292 14096 17320
rect 13780 17280 13786 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 15013 17323 15071 17329
rect 15013 17289 15025 17323
rect 15059 17320 15071 17323
rect 15194 17320 15200 17332
rect 15059 17292 15200 17320
rect 15059 17289 15071 17292
rect 15013 17283 15071 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 15470 17280 15476 17332
rect 15528 17280 15534 17332
rect 15838 17280 15844 17332
rect 15896 17280 15902 17332
rect 17218 17280 17224 17332
rect 17276 17320 17282 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 17276 17292 21189 17320
rect 17276 17280 17282 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 24578 17320 24584 17332
rect 21177 17283 21235 17289
rect 21284 17292 24584 17320
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17221 12035 17255
rect 11977 17215 12035 17221
rect 13538 17212 13544 17264
rect 13596 17252 13602 17264
rect 15488 17252 15516 17280
rect 13596 17224 15516 17252
rect 13596 17212 13602 17224
rect 20162 17212 20168 17264
rect 20220 17252 20226 17264
rect 21284 17252 21312 17292
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 25406 17280 25412 17332
rect 25464 17280 25470 17332
rect 20220 17224 21312 17252
rect 21545 17255 21603 17261
rect 20220 17212 20226 17224
rect 21545 17221 21557 17255
rect 21591 17252 21603 17255
rect 21726 17252 21732 17264
rect 21591 17224 21732 17252
rect 21591 17221 21603 17224
rect 21545 17215 21603 17221
rect 21726 17212 21732 17224
rect 21784 17252 21790 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21784 17224 22017 17252
rect 21784 17212 21790 17224
rect 22005 17221 22017 17224
rect 22051 17252 22063 17255
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 22051 17224 22201 17252
rect 22051 17221 22063 17224
rect 22005 17215 22063 17221
rect 22189 17221 22201 17224
rect 22235 17221 22247 17255
rect 22189 17215 22247 17221
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 22922 17252 22928 17264
rect 22520 17224 22928 17252
rect 22520 17212 22526 17224
rect 22922 17212 22928 17224
rect 22980 17212 22986 17264
rect 24210 17252 24216 17264
rect 24058 17224 24216 17252
rect 24210 17212 24216 17224
rect 24268 17252 24274 17264
rect 25222 17252 25228 17264
rect 24268 17224 25228 17252
rect 24268 17212 24274 17224
rect 25222 17212 25228 17224
rect 25280 17212 25286 17264
rect 6595 17156 7144 17184
rect 8113 17187 8171 17193
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8159 17156 8892 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 1946 17076 1952 17128
rect 2004 17076 2010 17128
rect 4522 17076 4528 17128
rect 4580 17076 4586 17128
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 8294 17116 8300 17128
rect 6871 17088 8300 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 5828 17048 5856 17079
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 7282 17048 7288 17060
rect 5828 17020 7288 17048
rect 7282 17008 7288 17020
rect 7340 17008 7346 17060
rect 3878 16940 3884 16992
rect 3936 16980 3942 16992
rect 5994 16980 6000 16992
rect 3936 16952 6000 16980
rect 3936 16940 3942 16952
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 8864 16980 8892 17156
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8996 17156 9229 17184
rect 8996 17144 9002 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 10870 17184 10876 17196
rect 10626 17156 10876 17184
rect 9217 17147 9275 17153
rect 10870 17144 10876 17156
rect 10928 17184 10934 17196
rect 11241 17187 11299 17193
rect 11241 17184 11253 17187
rect 10928 17156 11253 17184
rect 10928 17144 10934 17156
rect 11241 17153 11253 17156
rect 11287 17153 11299 17187
rect 11241 17147 11299 17153
rect 9490 17076 9496 17128
rect 9548 17076 9554 17128
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10100 17088 10977 17116
rect 10100 17076 10106 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 11256 17116 11284 17147
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 12710 17116 12716 17128
rect 11256 17088 12716 17116
rect 10965 17079 11023 17085
rect 12710 17076 12716 17088
rect 12768 17116 12774 17128
rect 12986 17116 12992 17128
rect 12768 17088 12992 17116
rect 12768 17076 12774 17088
rect 12986 17076 12992 17088
rect 13044 17116 13050 17128
rect 13096 17116 13124 17170
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 13688 17156 14381 17184
rect 13688 17144 13694 17156
rect 14369 17153 14381 17156
rect 14415 17184 14427 17187
rect 14642 17184 14648 17196
rect 14415 17156 14648 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 17678 17184 17684 17196
rect 17359 17156 17684 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 19628 17156 19734 17184
rect 13814 17116 13820 17128
rect 13044 17088 13820 17116
rect 13044 17076 13050 17088
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 14148 17088 15945 17116
rect 14148 17076 14154 17088
rect 15933 17085 15945 17088
rect 15979 17085 15991 17119
rect 15933 17079 15991 17085
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 11514 17048 11520 17060
rect 10520 17020 11520 17048
rect 10520 16980 10548 17020
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 16040 17048 16068 17079
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 16264 17088 17417 17116
rect 16264 17076 16270 17088
rect 17405 17085 17417 17088
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 13596 17020 16068 17048
rect 13596 17008 13602 17020
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 17770 17048 17776 17060
rect 16356 17020 17776 17048
rect 16356 17008 16362 17020
rect 17770 17008 17776 17020
rect 17828 17008 17834 17060
rect 8864 16952 10548 16980
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 13354 16980 13360 16992
rect 11112 16952 13360 16980
rect 11112 16940 11118 16952
rect 13354 16940 13360 16952
rect 13412 16940 13418 16992
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 14148 16952 15485 16980
rect 14148 16940 14154 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 17862 16940 17868 16992
rect 17920 16940 17926 16992
rect 18588 16983 18646 16989
rect 18588 16949 18600 16983
rect 18634 16980 18646 16983
rect 18966 16980 18972 16992
rect 18634 16952 18972 16980
rect 18634 16949 18646 16952
rect 18588 16943 18646 16949
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 19628 16980 19656 17156
rect 20254 17144 20260 17196
rect 20312 17184 20318 17196
rect 20533 17187 20591 17193
rect 20533 17184 20545 17187
rect 20312 17156 20545 17184
rect 20312 17144 20318 17156
rect 20533 17153 20545 17156
rect 20579 17153 20591 17187
rect 20533 17147 20591 17153
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 20680 17156 21833 17184
rect 20680 17144 20686 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 24857 17187 24915 17193
rect 24857 17153 24869 17187
rect 24903 17184 24915 17187
rect 25406 17184 25412 17196
rect 24903 17156 25412 17184
rect 24903 17153 24915 17156
rect 24857 17147 24915 17153
rect 25406 17144 25412 17156
rect 25464 17184 25470 17196
rect 26050 17184 26056 17196
rect 25464 17156 26056 17184
rect 25464 17144 25470 17156
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17116 20131 17119
rect 21450 17116 21456 17128
rect 20119 17088 21456 17116
rect 20119 17085 20131 17088
rect 20073 17079 20131 17085
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 22462 17076 22468 17128
rect 22520 17116 22526 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 22520 17088 22845 17116
rect 22520 17076 22526 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 22922 17076 22928 17128
rect 22980 17116 22986 17128
rect 24394 17116 24400 17128
rect 22980 17088 24400 17116
rect 22980 17076 22986 17088
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 22554 17048 22560 17060
rect 19760 17020 22560 17048
rect 19760 17008 19766 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 26694 17048 26700 17060
rect 25087 17020 26700 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 26694 17008 26700 17020
rect 26752 17008 26758 17060
rect 20806 16980 20812 16992
rect 19300 16952 20812 16980
rect 19300 16940 19306 16952
rect 20806 16940 20812 16952
rect 20864 16980 20870 16992
rect 21726 16980 21732 16992
rect 20864 16952 21732 16980
rect 20864 16940 20870 16952
rect 21726 16940 21732 16952
rect 21784 16940 21790 16992
rect 22646 16940 22652 16992
rect 22704 16980 22710 16992
rect 23382 16980 23388 16992
rect 22704 16952 23388 16980
rect 22704 16940 22710 16952
rect 23382 16940 23388 16952
rect 23440 16980 23446 16992
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 23440 16952 24317 16980
rect 23440 16940 23446 16952
rect 24305 16949 24317 16952
rect 24351 16949 24363 16983
rect 24305 16943 24363 16949
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 6914 16776 6920 16788
rect 2608 16748 2820 16776
rect 2608 16649 2636 16748
rect 2593 16643 2651 16649
rect 2593 16609 2605 16643
rect 2639 16609 2651 16643
rect 2593 16603 2651 16609
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2133 16575 2191 16581
rect 2133 16572 2145 16575
rect 1719 16544 2145 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2133 16541 2145 16544
rect 2179 16572 2191 16575
rect 2222 16572 2228 16584
rect 2179 16544 2228 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2792 16572 2820 16748
rect 2884 16748 6920 16776
rect 2884 16649 2912 16748
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 7524 16748 7573 16776
rect 7524 16736 7530 16748
rect 7561 16745 7573 16748
rect 7607 16745 7619 16779
rect 7561 16739 7619 16745
rect 9033 16779 9091 16785
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9122 16776 9128 16788
rect 9079 16748 9128 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9401 16779 9459 16785
rect 9401 16745 9413 16779
rect 9447 16776 9459 16779
rect 9674 16776 9680 16788
rect 9447 16748 9680 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 11146 16776 11152 16788
rect 10100 16748 11152 16776
rect 10100 16736 10106 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 14090 16776 14096 16788
rect 11348 16748 14096 16776
rect 3878 16708 3884 16720
rect 2976 16680 3884 16708
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16609 2927 16643
rect 2869 16603 2927 16609
rect 2976 16572 3004 16680
rect 3878 16668 3884 16680
rect 3936 16668 3942 16720
rect 4154 16668 4160 16720
rect 4212 16668 4218 16720
rect 6454 16708 6460 16720
rect 5184 16680 6460 16708
rect 3050 16600 3056 16652
rect 3108 16640 3114 16652
rect 5184 16649 5212 16680
rect 6454 16668 6460 16680
rect 6512 16668 6518 16720
rect 9214 16668 9220 16720
rect 9272 16708 9278 16720
rect 10778 16708 10784 16720
rect 9272 16680 10784 16708
rect 9272 16668 9278 16680
rect 10778 16668 10784 16680
rect 10836 16668 10842 16720
rect 3973 16643 4031 16649
rect 3973 16640 3985 16643
rect 3108 16612 3985 16640
rect 3108 16600 3114 16612
rect 3973 16609 3985 16612
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 5408 16612 5457 16640
rect 5408 16600 5414 16612
rect 5445 16609 5457 16612
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 5960 16612 6500 16640
rect 5960 16600 5966 16612
rect 2792 16544 3004 16572
rect 4706 16532 4712 16584
rect 4764 16532 4770 16584
rect 6472 16581 6500 16612
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6604 16612 6745 16640
rect 6604 16600 6610 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 6733 16603 6791 16609
rect 8220 16612 8585 16640
rect 8220 16581 8248 16612
rect 8573 16609 8585 16612
rect 8619 16640 8631 16643
rect 9398 16640 9404 16652
rect 8619 16612 9404 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 10594 16640 10600 16652
rect 9508 16612 10600 16640
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 9508 16572 9536 16612
rect 10594 16600 10600 16612
rect 10652 16640 10658 16652
rect 11054 16640 11060 16652
rect 10652 16612 11060 16640
rect 10652 16600 10658 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11348 16640 11376 16748
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 19150 16776 19156 16788
rect 17920 16748 19156 16776
rect 17920 16736 17926 16748
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 19444 16748 22094 16776
rect 15654 16668 15660 16720
rect 15712 16708 15718 16720
rect 16758 16708 16764 16720
rect 15712 16680 16764 16708
rect 15712 16668 15718 16680
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 11287 16612 11376 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11422 16600 11428 16652
rect 11480 16600 11486 16652
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 13998 16640 14004 16652
rect 12299 16612 14004 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14918 16640 14924 16652
rect 14323 16612 14924 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 19150 16640 19156 16652
rect 17451 16612 19156 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19444 16649 19472 16748
rect 21637 16711 21695 16717
rect 21637 16677 21649 16711
rect 21683 16677 21695 16711
rect 21637 16671 21695 16677
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 19702 16600 19708 16652
rect 19760 16600 19766 16652
rect 8803 16544 9536 16572
rect 9677 16575 9735 16581
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 9723 16544 11560 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 5442 16464 5448 16516
rect 5500 16504 5506 16516
rect 5500 16476 5948 16504
rect 5500 16464 5506 16476
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16436 2007 16439
rect 2038 16436 2044 16448
rect 1995 16408 2044 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 5718 16436 5724 16448
rect 4571 16408 5724 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5920 16436 5948 16476
rect 5994 16464 6000 16516
rect 6052 16504 6058 16516
rect 6052 16476 10824 16504
rect 6052 16464 6058 16476
rect 7558 16436 7564 16448
rect 5920 16408 7564 16436
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 8021 16439 8079 16445
rect 8021 16405 8033 16439
rect 8067 16436 8079 16439
rect 8662 16436 8668 16448
rect 8067 16408 8668 16436
rect 8067 16405 8079 16408
rect 8021 16399 8079 16405
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 9125 16439 9183 16445
rect 9125 16436 9137 16439
rect 8996 16408 9137 16436
rect 8996 16396 9002 16408
rect 9125 16405 9137 16408
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9766 16436 9772 16448
rect 9456 16408 9772 16436
rect 9456 16396 9462 16408
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 10318 16396 10324 16448
rect 10376 16396 10382 16448
rect 10796 16445 10824 16476
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 10870 16396 10876 16448
rect 10928 16436 10934 16448
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 10928 16408 11161 16436
rect 10928 16396 10934 16408
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11532 16436 11560 16544
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16572 16727 16575
rect 16758 16572 16764 16584
rect 16715 16544 16764 16572
rect 16715 16541 16727 16544
rect 16669 16535 16727 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17126 16532 17132 16584
rect 17184 16532 17190 16584
rect 18966 16532 18972 16584
rect 19024 16572 19030 16584
rect 19242 16572 19248 16584
rect 19024 16544 19248 16572
rect 19024 16532 19030 16544
rect 19242 16532 19248 16544
rect 19300 16532 19306 16584
rect 20806 16532 20812 16584
rect 20864 16532 20870 16584
rect 21652 16572 21680 16671
rect 22066 16640 22094 16748
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 23106 16776 23112 16788
rect 22336 16748 23112 16776
rect 22336 16736 22342 16748
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 22278 16640 22284 16652
rect 22066 16612 22284 16640
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 25130 16640 25136 16652
rect 22603 16612 25136 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 26142 16600 26148 16652
rect 26200 16600 26206 16652
rect 21008 16544 21680 16572
rect 21821 16575 21879 16581
rect 12710 16464 12716 16516
rect 12768 16464 12774 16516
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 14516 16476 14565 16504
rect 14516 16464 14522 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 14553 16467 14611 16473
rect 15010 16464 15016 16516
rect 15068 16464 15074 16516
rect 17310 16464 17316 16516
rect 17368 16504 17374 16516
rect 17862 16504 17868 16516
rect 17368 16476 17868 16504
rect 17368 16464 17374 16476
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 19426 16504 19432 16516
rect 18708 16476 19432 16504
rect 12342 16436 12348 16448
rect 11532 16408 12348 16436
rect 11149 16399 11207 16405
rect 12342 16396 12348 16408
rect 12400 16436 12406 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12400 16408 13737 16436
rect 12400 16396 12406 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 16206 16436 16212 16448
rect 14056 16408 16212 16436
rect 14056 16396 14062 16408
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16485 16439 16543 16445
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 18708 16436 18736 16476
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 16531 16408 18736 16436
rect 18877 16439 18935 16445
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 18877 16405 18889 16439
rect 18923 16436 18935 16439
rect 20346 16436 20352 16448
rect 18923 16408 20352 16436
rect 18923 16405 18935 16408
rect 18877 16399 18935 16405
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 21008 16436 21036 16544
rect 21821 16541 21833 16575
rect 21867 16572 21879 16575
rect 24210 16572 24216 16584
rect 21867 16544 22324 16572
rect 23690 16544 24216 16572
rect 21867 16541 21879 16544
rect 21821 16535 21879 16541
rect 22296 16504 22324 16544
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 22646 16504 22652 16516
rect 21468 16476 22094 16504
rect 22296 16476 22652 16504
rect 20496 16408 21036 16436
rect 21177 16439 21235 16445
rect 20496 16396 20502 16408
rect 21177 16405 21189 16439
rect 21223 16436 21235 16439
rect 21358 16436 21364 16448
rect 21223 16408 21364 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21358 16396 21364 16408
rect 21416 16436 21422 16448
rect 21468 16436 21496 16476
rect 21416 16408 21496 16436
rect 22066 16436 22094 16476
rect 22646 16464 22652 16476
rect 22704 16464 22710 16516
rect 24596 16504 24624 16535
rect 23860 16476 24624 16504
rect 23860 16436 23888 16476
rect 22066 16408 23888 16436
rect 21416 16396 21422 16408
rect 24026 16396 24032 16448
rect 24084 16396 24090 16448
rect 25222 16396 25228 16448
rect 25280 16396 25286 16448
rect 25774 16396 25780 16448
rect 25832 16436 25838 16448
rect 25958 16436 25964 16448
rect 25832 16408 25964 16436
rect 25832 16396 25838 16408
rect 25958 16396 25964 16408
rect 26016 16396 26022 16448
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 26050 16328 26056 16380
rect 26108 16368 26114 16380
rect 26160 16368 26188 16600
rect 26108 16340 26188 16368
rect 26108 16328 26114 16340
rect 1104 16272 25852 16294
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 9122 16232 9128 16244
rect 5859 16204 9128 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 9122 16192 9128 16204
rect 9180 16192 9186 16244
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 9953 16235 10011 16241
rect 9953 16232 9965 16235
rect 9548 16204 9965 16232
rect 9548 16192 9554 16204
rect 9953 16201 9965 16204
rect 9999 16201 10011 16235
rect 10870 16232 10876 16244
rect 9953 16195 10011 16201
rect 10060 16204 10876 16232
rect 2961 16167 3019 16173
rect 2961 16133 2973 16167
rect 3007 16164 3019 16167
rect 3510 16164 3516 16176
rect 3007 16136 3516 16164
rect 3007 16133 3019 16136
rect 2961 16127 3019 16133
rect 3510 16124 3516 16136
rect 3568 16124 3574 16176
rect 6638 16164 6644 16176
rect 4540 16136 6644 16164
rect 1854 16056 1860 16108
rect 1912 16056 1918 16108
rect 3237 16099 3295 16105
rect 3237 16065 3249 16099
rect 3283 16096 3295 16099
rect 3418 16096 3424 16108
rect 3283 16068 3424 16096
rect 3283 16065 3295 16068
rect 3237 16059 3295 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 4540 16105 4568 16136
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 10060 16164 10088 16204
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 11296 16204 13921 16232
rect 11296 16192 11302 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 14415 16204 19349 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 19337 16201 19349 16204
rect 19383 16201 19395 16235
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 19337 16195 19395 16201
rect 19444 16204 21005 16232
rect 6748 16136 10088 16164
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 5350 16096 5356 16108
rect 4847 16068 5356 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6362 16096 6368 16108
rect 6043 16068 6368 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 6362 16056 6368 16068
rect 6420 16096 6426 16108
rect 6457 16099 6515 16105
rect 6457 16096 6469 16099
rect 6420 16068 6469 16096
rect 6420 16056 6426 16068
rect 6457 16065 6469 16068
rect 6503 16065 6515 16099
rect 6457 16059 6515 16065
rect 6546 16056 6552 16108
rect 6604 16096 6610 16108
rect 6748 16096 6776 16136
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 11977 16167 12035 16173
rect 11977 16164 11989 16167
rect 10376 16136 11989 16164
rect 10376 16124 10382 16136
rect 11977 16133 11989 16136
rect 12023 16133 12035 16167
rect 11977 16127 12035 16133
rect 12710 16124 12716 16176
rect 12768 16124 12774 16176
rect 15197 16167 15255 16173
rect 15197 16133 15209 16167
rect 15243 16164 15255 16167
rect 15286 16164 15292 16176
rect 15243 16136 15292 16164
rect 15243 16133 15255 16136
rect 15197 16127 15255 16133
rect 15286 16124 15292 16136
rect 15344 16164 15350 16176
rect 15933 16167 15991 16173
rect 15933 16164 15945 16167
rect 15344 16136 15945 16164
rect 15344 16124 15350 16136
rect 15933 16133 15945 16136
rect 15979 16133 15991 16167
rect 15933 16127 15991 16133
rect 16390 16124 16396 16176
rect 16448 16164 16454 16176
rect 16448 16136 19104 16164
rect 16448 16124 16454 16136
rect 6604 16068 6776 16096
rect 6604 16056 6610 16068
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 7248 16068 7297 16096
rect 7248 16056 7254 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 8297 16099 8355 16105
rect 8297 16096 8309 16099
rect 7616 16068 8309 16096
rect 7616 16056 7622 16068
rect 8297 16065 8309 16068
rect 8343 16065 8355 16099
rect 8297 16059 8355 16065
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9030 16096 9036 16108
rect 8895 16068 9036 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 2777 16031 2835 16037
rect 2777 16028 2789 16031
rect 1627 16000 2789 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 2777 15997 2789 16000
rect 2823 16028 2835 16031
rect 3326 16028 3332 16040
rect 2823 16000 3332 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 15997 3571 16031
rect 7009 16031 7067 16037
rect 7009 16028 7021 16031
rect 3513 15991 3571 15997
rect 4908 16000 7021 16028
rect 3528 15892 3556 15991
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 4908 15960 4936 16000
rect 7009 15997 7021 16000
rect 7055 15997 7067 16031
rect 8312 16028 8340 16059
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9306 16056 9312 16108
rect 9364 16056 9370 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 9640 16068 10793 16096
rect 9640 16056 9646 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 10686 16028 10692 16040
rect 8312 16000 10692 16028
rect 7009 15991 7067 15997
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 4212 15932 4936 15960
rect 4212 15920 4218 15932
rect 6638 15920 6644 15972
rect 6696 15960 6702 15972
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 6696 15932 10425 15960
rect 6696 15920 6702 15932
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 7098 15892 7104 15904
rect 3528 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 8113 15895 8171 15901
rect 8113 15892 8125 15895
rect 7248 15864 8125 15892
rect 7248 15852 7254 15864
rect 8113 15861 8125 15864
rect 8159 15861 8171 15895
rect 8113 15855 8171 15861
rect 8662 15852 8668 15904
rect 8720 15852 8726 15904
rect 10888 15892 10916 15991
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11974 15988 11980 16040
rect 12032 16028 12038 16040
rect 14292 16028 14320 16059
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 18966 16096 18972 16108
rect 17175 16068 18972 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18966 16056 18972 16068
rect 19024 16056 19030 16108
rect 19076 16096 19104 16136
rect 19444 16096 19472 16204
rect 20993 16201 21005 16204
rect 21039 16201 21051 16235
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 20993 16195 21051 16201
rect 21100 16204 21680 16232
rect 21100 16164 21128 16204
rect 19076 16068 19472 16096
rect 19536 16136 21128 16164
rect 21545 16167 21603 16173
rect 12032 16000 14320 16028
rect 12032 15988 12038 16000
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 16022 15988 16028 16040
rect 16080 15988 16086 16040
rect 18877 16031 18935 16037
rect 18877 15997 18889 16031
rect 18923 16028 18935 16031
rect 19058 16028 19064 16040
rect 18923 16000 19064 16028
rect 18923 15997 18935 16000
rect 18877 15991 18935 15997
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19536 16028 19564 16136
rect 21545 16133 21557 16167
rect 21591 16133 21603 16167
rect 21545 16127 21603 16133
rect 19610 16056 19616 16108
rect 19668 16096 19674 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19668 16068 19717 16096
rect 19668 16056 19674 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 19843 16068 20300 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 19300 16000 19564 16028
rect 19981 16031 20039 16037
rect 19300 15988 19306 16000
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 20162 16028 20168 16040
rect 20027 16000 20168 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 20272 16028 20300 16068
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20772 16068 20913 16096
rect 20772 16056 20778 16068
rect 20901 16065 20913 16068
rect 20947 16065 20959 16099
rect 21560 16096 21588 16127
rect 20901 16059 20959 16065
rect 21008 16068 21588 16096
rect 21652 16096 21680 16204
rect 22066 16204 23213 16232
rect 21726 16124 21732 16176
rect 21784 16164 21790 16176
rect 22066 16164 22094 16204
rect 23201 16201 23213 16204
rect 23247 16232 23259 16235
rect 23753 16235 23811 16241
rect 23753 16232 23765 16235
rect 23247 16204 23765 16232
rect 23247 16201 23259 16204
rect 23201 16195 23259 16201
rect 23753 16201 23765 16204
rect 23799 16201 23811 16235
rect 23753 16195 23811 16201
rect 23842 16192 23848 16244
rect 23900 16192 23906 16244
rect 25222 16164 25228 16176
rect 21784 16136 22094 16164
rect 22296 16136 25228 16164
rect 21784 16124 21790 16136
rect 22296 16096 22324 16136
rect 25222 16124 25228 16136
rect 25280 16124 25286 16176
rect 21652 16068 22324 16096
rect 22373 16099 22431 16105
rect 20530 16028 20536 16040
rect 20272 16000 20536 16028
rect 20530 15988 20536 16000
rect 20588 16028 20594 16040
rect 21008 16028 21036 16068
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22419 16068 23029 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 20588 16000 21036 16028
rect 20588 15988 20594 16000
rect 21174 15988 21180 16040
rect 21232 15988 21238 16040
rect 22094 16028 22100 16040
rect 21284 16000 22100 16028
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 13372 15932 15485 15960
rect 13372 15892 13400 15932
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 15473 15923 15531 15929
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 21284 15960 21312 16000
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22388 16028 22416 16059
rect 23106 16056 23112 16108
rect 23164 16096 23170 16108
rect 23474 16096 23480 16108
rect 23164 16068 23480 16096
rect 23164 16056 23170 16068
rect 23474 16056 23480 16068
rect 23532 16096 23538 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 23532 16068 24593 16096
rect 23532 16056 23538 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 22244 16000 22416 16028
rect 22465 16031 22523 16037
rect 22244 15988 22250 16000
rect 22465 15997 22477 16031
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22557 16031 22615 16037
rect 22557 15997 22569 16031
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 16816 15932 21312 15960
rect 16816 15920 16822 15932
rect 21634 15920 21640 15972
rect 21692 15960 21698 15972
rect 22480 15960 22508 15991
rect 21692 15932 22508 15960
rect 21692 15920 21698 15932
rect 10888 15864 13400 15892
rect 13449 15895 13507 15901
rect 13449 15861 13461 15895
rect 13495 15892 13507 15895
rect 13538 15892 13544 15904
rect 13495 15864 13544 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14550 15892 14556 15904
rect 14240 15864 14556 15892
rect 14240 15852 14246 15864
rect 14550 15852 14556 15864
rect 14608 15852 14614 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16264 15864 16681 15892
rect 16264 15852 16270 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 20530 15852 20536 15904
rect 20588 15852 20594 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 20680 15864 22017 15892
rect 20680 15852 20686 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 22572 15892 22600 15991
rect 24026 15988 24032 16040
rect 24084 15988 24090 16040
rect 22646 15920 22652 15972
rect 22704 15960 22710 15972
rect 25225 15963 25283 15969
rect 25225 15960 25237 15963
rect 22704 15932 25237 15960
rect 22704 15920 22710 15932
rect 25225 15929 25237 15932
rect 25271 15929 25283 15963
rect 25225 15923 25283 15929
rect 22428 15864 22600 15892
rect 22428 15852 22434 15864
rect 23382 15852 23388 15904
rect 23440 15852 23446 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 4706 15688 4712 15700
rect 1995 15660 4712 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 5813 15691 5871 15697
rect 5813 15657 5825 15691
rect 5859 15688 5871 15691
rect 6086 15688 6092 15700
rect 5859 15660 6092 15688
rect 5859 15657 5871 15660
rect 5813 15651 5871 15657
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 6454 15648 6460 15700
rect 6512 15648 6518 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 6880 15660 7113 15688
rect 6880 15648 6886 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 12618 15688 12624 15700
rect 8720 15660 12624 15688
rect 8720 15648 8726 15660
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 16850 15688 16856 15700
rect 13188 15660 16856 15688
rect 10502 15620 10508 15632
rect 8404 15592 10508 15620
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 2869 15555 2927 15561
rect 2869 15552 2881 15555
rect 2832 15524 2881 15552
rect 2832 15512 2838 15524
rect 2869 15521 2881 15524
rect 2915 15521 2927 15555
rect 2869 15515 2927 15521
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 8202 15552 8208 15564
rect 4847 15524 8208 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8404 15561 8432 15592
rect 10502 15580 10508 15592
rect 10560 15580 10566 15632
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 12066 15552 12072 15564
rect 10827 15524 12072 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13188 15561 13216 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 19150 15648 19156 15700
rect 19208 15688 19214 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 19208 15660 23673 15688
rect 19208 15648 19214 15660
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 23750 15648 23756 15700
rect 23808 15688 23814 15700
rect 24210 15688 24216 15700
rect 23808 15660 24216 15688
rect 23808 15648 23814 15660
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 16669 15623 16727 15629
rect 16669 15589 16681 15623
rect 16715 15620 16727 15623
rect 16758 15620 16764 15632
rect 16715 15592 16764 15620
rect 16715 15589 16727 15592
rect 16669 15583 16727 15589
rect 16758 15580 16764 15592
rect 16816 15580 16822 15632
rect 20530 15580 20536 15632
rect 20588 15620 20594 15632
rect 20588 15592 22968 15620
rect 20588 15580 20594 15592
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13354 15512 13360 15564
rect 13412 15512 13418 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 16850 15552 16856 15564
rect 14332 15524 16856 15552
rect 14332 15512 14338 15524
rect 16850 15512 16856 15524
rect 16908 15552 16914 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16908 15524 16957 15552
rect 16908 15512 16914 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 18693 15555 18751 15561
rect 18693 15521 18705 15555
rect 18739 15521 18751 15555
rect 18693 15515 18751 15521
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 4430 15484 4436 15496
rect 2639 15456 4436 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 2148 15416 2176 15447
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 5534 15484 5540 15496
rect 4571 15456 5540 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5994 15444 6000 15496
rect 6052 15444 6058 15496
rect 6638 15444 6644 15496
rect 6696 15444 6702 15496
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7248 15456 7297 15484
rect 7248 15444 7254 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7285 15447 7343 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8754 15484 8760 15496
rect 7975 15456 8760 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 9953 15487 10011 15493
rect 9953 15484 9965 15487
rect 9732 15456 9965 15484
rect 9732 15444 9738 15456
rect 9953 15453 9965 15456
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 12342 15484 12348 15496
rect 11914 15456 12348 15484
rect 10505 15447 10563 15453
rect 10226 15416 10232 15428
rect 2148 15388 10232 15416
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 10520 15416 10548 15447
rect 12342 15444 12348 15456
rect 12400 15484 12406 15496
rect 12710 15484 12716 15496
rect 12400 15456 12716 15484
rect 12400 15444 12406 15456
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13906 15484 13912 15496
rect 13127 15456 13912 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 18708 15484 18736 15515
rect 19978 15512 19984 15564
rect 20036 15512 20042 15564
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15552 20223 15555
rect 20254 15552 20260 15564
rect 20211 15524 20260 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 21177 15555 21235 15561
rect 21177 15521 21189 15555
rect 21223 15552 21235 15555
rect 21266 15552 21272 15564
rect 21223 15524 21272 15552
rect 21223 15521 21235 15524
rect 21177 15515 21235 15521
rect 21266 15512 21272 15524
rect 21324 15512 21330 15564
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 22940 15552 22968 15592
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 23474 15620 23480 15632
rect 23072 15592 23480 15620
rect 23072 15580 23078 15592
rect 23474 15580 23480 15592
rect 23532 15580 23538 15632
rect 25774 15552 25780 15564
rect 21508 15524 22094 15552
rect 22940 15524 25780 15552
rect 21508 15512 21514 15524
rect 19886 15484 19892 15496
rect 18708 15456 19892 15484
rect 19886 15444 19892 15456
rect 19944 15484 19950 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 19944 15456 21925 15484
rect 19944 15444 19950 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 22066 15484 22094 15524
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22066 15456 23029 15484
rect 21913 15447 21971 15453
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 24026 15444 24032 15496
rect 24084 15484 24090 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24084 15456 24593 15484
rect 24084 15444 24090 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 10870 15416 10876 15428
rect 10520 15388 10876 15416
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 12728 15416 12756 15444
rect 12728 15388 12940 15416
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 4430 15348 4436 15360
rect 3927 15320 4436 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 7745 15351 7803 15357
rect 7745 15348 7757 15351
rect 7248 15320 7757 15348
rect 7248 15308 7254 15320
rect 7745 15317 7757 15320
rect 7791 15317 7803 15351
rect 7745 15311 7803 15317
rect 9122 15308 9128 15360
rect 9180 15308 9186 15360
rect 9766 15308 9772 15360
rect 9824 15308 9830 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 11422 15348 11428 15360
rect 10560 15320 11428 15348
rect 10560 15308 10566 15320
rect 11422 15308 11428 15320
rect 11480 15348 11486 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 11480 15320 12265 15348
rect 11480 15308 11486 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 12710 15308 12716 15360
rect 12768 15308 12774 15360
rect 12912 15348 12940 15388
rect 14550 15376 14556 15428
rect 14608 15376 14614 15428
rect 15010 15376 15016 15428
rect 15068 15376 15074 15428
rect 17218 15376 17224 15428
rect 17276 15416 17282 15428
rect 21085 15419 21143 15425
rect 17276 15388 17710 15416
rect 17276 15376 17282 15388
rect 13630 15348 13636 15360
rect 12912 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15348 13694 15360
rect 13725 15351 13783 15357
rect 13725 15348 13737 15351
rect 13688 15320 13737 15348
rect 13688 15308 13694 15320
rect 13725 15317 13737 15320
rect 13771 15317 13783 15351
rect 13725 15311 13783 15317
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 16025 15351 16083 15357
rect 16025 15348 16037 15351
rect 14700 15320 16037 15348
rect 14700 15308 14706 15320
rect 16025 15317 16037 15320
rect 16071 15317 16083 15351
rect 16025 15311 16083 15317
rect 16206 15308 16212 15360
rect 16264 15348 16270 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16264 15320 16313 15348
rect 16264 15308 16270 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 17604 15348 17632 15388
rect 21085 15385 21097 15419
rect 21131 15416 21143 15419
rect 21266 15416 21272 15428
rect 21131 15388 21272 15416
rect 21131 15385 21143 15388
rect 21085 15379 21143 15385
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 21818 15376 21824 15428
rect 21876 15416 21882 15428
rect 23290 15416 23296 15428
rect 21876 15388 23296 15416
rect 21876 15376 21882 15388
rect 23290 15376 23296 15388
rect 23348 15376 23354 15428
rect 23474 15376 23480 15428
rect 23532 15416 23538 15428
rect 23937 15419 23995 15425
rect 23937 15416 23949 15419
rect 23532 15388 23949 15416
rect 23532 15376 23538 15388
rect 23937 15385 23949 15388
rect 23983 15385 23995 15419
rect 23937 15379 23995 15385
rect 18969 15351 19027 15357
rect 18969 15348 18981 15351
rect 17604 15320 18981 15348
rect 16301 15311 16359 15317
rect 18969 15317 18981 15320
rect 19015 15317 19027 15351
rect 18969 15311 19027 15317
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 19521 15351 19579 15357
rect 19521 15348 19533 15351
rect 19208 15320 19533 15348
rect 19208 15308 19214 15320
rect 19521 15317 19533 15320
rect 19567 15317 19579 15351
rect 19521 15311 19579 15317
rect 19886 15308 19892 15360
rect 19944 15308 19950 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 21542 15348 21548 15360
rect 20763 15320 21548 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 21542 15308 21548 15320
rect 21600 15308 21606 15360
rect 22554 15308 22560 15360
rect 22612 15308 22618 15360
rect 23750 15308 23756 15360
rect 23808 15348 23814 15360
rect 24026 15348 24032 15360
rect 23808 15320 24032 15348
rect 23808 15308 23814 15320
rect 24026 15308 24032 15320
rect 24084 15308 24090 15360
rect 24302 15308 24308 15360
rect 24360 15348 24366 15360
rect 25225 15351 25283 15357
rect 25225 15348 25237 15351
rect 24360 15320 25237 15348
rect 24360 15308 24366 15320
rect 25225 15317 25237 15320
rect 25271 15317 25283 15351
rect 25225 15311 25283 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 1360 15116 1777 15144
rect 1360 15104 1366 15116
rect 1765 15113 1777 15116
rect 1811 15144 1823 15147
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1811 15116 1961 15144
rect 1811 15113 1823 15116
rect 1765 15107 1823 15113
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2096 15116 2605 15144
rect 2096 15104 2102 15116
rect 2593 15113 2605 15116
rect 2639 15113 2651 15147
rect 2593 15107 2651 15113
rect 3786 15104 3792 15156
rect 3844 15104 3850 15156
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 4580 15116 5825 15144
rect 4580 15104 4586 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 8570 15144 8576 15156
rect 5813 15107 5871 15113
rect 6012 15116 8576 15144
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3804 15008 3832 15104
rect 5534 15036 5540 15088
rect 5592 15036 5598 15088
rect 6012 15017 6040 15116
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 9214 15104 9220 15156
rect 9272 15104 9278 15156
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 9950 15144 9956 15156
rect 9907 15116 9956 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11882 15144 11888 15156
rect 11112 15116 11888 15144
rect 11112 15104 11118 15116
rect 11882 15104 11888 15116
rect 11940 15144 11946 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 11940 15116 13461 15144
rect 11940 15104 11946 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13630 15104 13636 15156
rect 13688 15144 13694 15156
rect 13725 15147 13783 15153
rect 13725 15144 13737 15147
rect 13688 15116 13737 15144
rect 13688 15104 13694 15116
rect 13725 15113 13737 15116
rect 13771 15144 13783 15147
rect 13814 15144 13820 15156
rect 13771 15116 13820 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 14608 15116 16313 15144
rect 14608 15104 14614 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 16301 15107 16359 15113
rect 17144 15116 18920 15144
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 7892 15048 10272 15076
rect 7892 15036 7898 15048
rect 3467 14980 3832 15008
rect 5997 15011 6055 15017
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 5997 14977 6009 15011
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 8481 15011 8539 15017
rect 6871 14980 8432 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3752 14912 4077 14940
rect 3752 14900 3758 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 4338 14900 4344 14952
rect 4396 14900 4402 14952
rect 6546 14900 6552 14952
rect 6604 14900 6610 14952
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8294 14940 8300 14952
rect 7975 14912 8300 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8404 14940 8432 14980
rect 8481 14977 8493 15011
rect 8527 15008 8539 15011
rect 8754 15008 8760 15020
rect 8527 14980 8760 15008
rect 8527 14977 8539 14980
rect 8481 14971 8539 14977
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 9272 14980 9413 15008
rect 9272 14968 9278 14980
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10045 15011 10103 15017
rect 10045 15008 10057 15011
rect 9916 14980 10057 15008
rect 9916 14968 9922 14980
rect 10045 14977 10057 14980
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10134 14940 10140 14952
rect 8404 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 10244 14940 10272 15048
rect 10318 15036 10324 15088
rect 10376 15076 10382 15088
rect 11606 15076 11612 15088
rect 10376 15048 11612 15076
rect 10376 15036 10382 15048
rect 11606 15036 11612 15048
rect 11664 15036 11670 15088
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 12250 15076 12256 15088
rect 12023 15048 12256 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 12618 15036 12624 15088
rect 12676 15036 12682 15088
rect 15010 15036 15016 15088
rect 15068 15076 15074 15088
rect 15289 15079 15347 15085
rect 15289 15076 15301 15079
rect 15068 15048 15301 15076
rect 15068 15036 15074 15048
rect 15289 15045 15301 15048
rect 15335 15076 15347 15079
rect 16206 15076 16212 15088
rect 15335 15048 16212 15076
rect 15335 15045 15347 15048
rect 15289 15039 15347 15045
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 17144 15085 17172 15116
rect 17129 15079 17187 15085
rect 17129 15045 17141 15079
rect 17175 15045 17187 15079
rect 17129 15039 17187 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 18892 15076 18920 15116
rect 18966 15104 18972 15156
rect 19024 15104 19030 15156
rect 22554 15144 22560 15156
rect 19628 15116 22560 15144
rect 19628 15076 19656 15116
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 23014 15144 23020 15156
rect 22664 15116 23020 15144
rect 17276 15048 17618 15076
rect 18892 15048 19656 15076
rect 21637 15079 21695 15085
rect 17276 15036 17282 15048
rect 21637 15045 21649 15079
rect 21683 15076 21695 15079
rect 22002 15076 22008 15088
rect 21683 15048 22008 15076
rect 21683 15045 21695 15048
rect 21637 15039 21695 15045
rect 22002 15036 22008 15048
rect 22060 15036 22066 15088
rect 22094 15036 22100 15088
rect 22152 15036 22158 15088
rect 22664 15076 22692 15116
rect 23014 15104 23020 15116
rect 23072 15104 23078 15156
rect 23290 15104 23296 15156
rect 23348 15144 23354 15156
rect 23348 15116 25176 15144
rect 23348 15104 23354 15116
rect 22204 15048 22692 15076
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 11698 15008 11704 15020
rect 10928 14980 11704 15008
rect 10928 14968 10934 14980
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 16574 15008 16580 15020
rect 15703 14980 16580 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16816 14980 16865 15008
rect 16816 14968 16822 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 20714 14968 20720 15020
rect 20772 14968 20778 15020
rect 17862 14940 17868 14952
rect 10244 14912 11376 14940
rect 3237 14875 3295 14881
rect 3237 14841 3249 14875
rect 3283 14872 3295 14875
rect 6730 14872 6736 14884
rect 3283 14844 6736 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 11348 14872 11376 14912
rect 11808 14912 15516 14940
rect 11808 14872 11836 14912
rect 7616 14844 11284 14872
rect 11348 14844 11836 14872
rect 7616 14832 7622 14844
rect 7837 14807 7895 14813
rect 7837 14773 7849 14807
rect 7883 14804 7895 14807
rect 8294 14804 8300 14816
rect 7883 14776 8300 14804
rect 7883 14773 7895 14776
rect 7837 14767 7895 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 8570 14764 8576 14816
rect 8628 14764 8634 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 11020 14776 11161 14804
rect 11020 14764 11026 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11256 14804 11284 14844
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 15378 14872 15384 14884
rect 13688 14844 15384 14872
rect 13688 14832 13694 14844
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 15488 14872 15516 14912
rect 16960 14912 17868 14940
rect 16960 14872 16988 14912
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 19334 14940 19340 14952
rect 18156 14912 19340 14940
rect 15488 14844 16988 14872
rect 13722 14804 13728 14816
rect 11256 14776 13728 14804
rect 11149 14767 11207 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14829 14807 14887 14813
rect 14829 14804 14841 14807
rect 14608 14776 14841 14804
rect 14608 14764 14614 14776
rect 14829 14773 14841 14776
rect 14875 14773 14887 14807
rect 14829 14767 14887 14773
rect 15194 14764 15200 14816
rect 15252 14764 15258 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 17126 14804 17132 14816
rect 16816 14776 17132 14804
rect 16816 14764 16822 14776
rect 17126 14764 17132 14776
rect 17184 14804 17190 14816
rect 18156 14804 18184 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 21085 14943 21143 14949
rect 19659 14912 21036 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 18601 14875 18659 14881
rect 18601 14841 18613 14875
rect 18647 14872 18659 14875
rect 19242 14872 19248 14884
rect 18647 14844 19248 14872
rect 18647 14841 18659 14844
rect 18601 14835 18659 14841
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 21008 14872 21036 14912
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 22204 14940 22232 15048
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 25148 15085 25176 15116
rect 25133 15079 25191 15085
rect 25133 15045 25145 15079
rect 25179 15045 25191 15079
rect 25133 15039 25191 15045
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22336 14980 22845 15008
rect 22336 14968 22342 14980
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 21131 14912 22232 14940
rect 23109 14943 23167 14949
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 23109 14909 23121 14943
rect 23155 14940 23167 14943
rect 24302 14940 24308 14952
rect 23155 14912 24308 14940
rect 23155 14909 23167 14912
rect 23109 14903 23167 14909
rect 24302 14900 24308 14912
rect 24360 14900 24366 14952
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 24544 14912 24593 14940
rect 24544 14900 24550 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 22830 14872 22836 14884
rect 21008 14844 22836 14872
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 17184 14776 18184 14804
rect 17184 14764 17190 14776
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 18932 14776 21373 14804
rect 18932 14764 18938 14776
rect 21361 14773 21373 14776
rect 21407 14804 21419 14807
rect 21818 14804 21824 14816
rect 21407 14776 21824 14804
rect 21407 14773 21419 14776
rect 21361 14767 21419 14773
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 23750 14804 23756 14816
rect 22235 14776 23756 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 23750 14764 23756 14776
rect 23808 14764 23814 14816
rect 25222 14764 25228 14816
rect 25280 14764 25286 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2832 14572 2881 14600
rect 2832 14560 2838 14572
rect 2869 14569 2881 14572
rect 2915 14569 2927 14603
rect 2869 14563 2927 14569
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 4246 14600 4252 14612
rect 4203 14572 4252 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4614 14560 4620 14612
rect 4672 14600 4678 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 4672 14572 4721 14600
rect 4672 14560 4678 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 4709 14563 4767 14569
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 6454 14600 6460 14612
rect 4856 14572 6460 14600
rect 4856 14560 4862 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 6604 14572 9321 14600
rect 6604 14560 6610 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 10796 14572 12020 14600
rect 3237 14535 3295 14541
rect 3237 14501 3249 14535
rect 3283 14532 3295 14535
rect 5626 14532 5632 14544
rect 3283 14504 5632 14532
rect 3283 14501 3295 14504
rect 3237 14495 3295 14501
rect 5626 14492 5632 14504
rect 5684 14492 5690 14544
rect 7742 14532 7748 14544
rect 6012 14504 7748 14532
rect 2314 14356 2320 14408
rect 2372 14356 2378 14408
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2823 14368 3433 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 3421 14365 3433 14368
rect 3467 14396 3479 14399
rect 3510 14396 3516 14408
rect 3467 14368 3516 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 4890 14356 4896 14408
rect 4948 14356 4954 14408
rect 5534 14356 5540 14408
rect 5592 14356 5598 14408
rect 6012 14405 6040 14504
rect 7742 14492 7748 14504
rect 7800 14492 7806 14544
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 8386 14532 8392 14544
rect 7892 14504 8392 14532
rect 7892 14492 7898 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 10045 14535 10103 14541
rect 10045 14501 10057 14535
rect 10091 14532 10103 14535
rect 10410 14532 10416 14544
rect 10091 14504 10416 14532
rect 10091 14501 10103 14504
rect 10045 14495 10103 14501
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 9950 14464 9956 14476
rect 6144 14436 9956 14464
rect 6144 14424 6150 14436
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10796 14464 10824 14572
rect 11992 14532 12020 14572
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 12124 14572 13553 14600
rect 12124 14560 12130 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 16022 14600 16028 14612
rect 13541 14563 13599 14569
rect 13740 14572 16028 14600
rect 12437 14535 12495 14541
rect 11992 14504 12112 14532
rect 10152 14436 10824 14464
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6270 14356 6276 14408
rect 6328 14356 6334 14408
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 7834 14396 7840 14408
rect 7515 14368 7840 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 7834 14356 7840 14368
rect 7892 14356 7898 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 8846 14396 8852 14408
rect 8435 14368 8852 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 10152 14396 10180 14436
rect 10962 14424 10968 14476
rect 11020 14424 11026 14476
rect 12084 14464 12112 14504
rect 12437 14501 12449 14535
rect 12483 14532 12495 14535
rect 12618 14532 12624 14544
rect 12483 14504 12624 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 12618 14492 12624 14504
rect 12676 14532 12682 14544
rect 13740 14532 13768 14572
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 16758 14600 16764 14612
rect 16592 14572 16764 14600
rect 12676 14504 13768 14532
rect 12676 14492 12682 14504
rect 13814 14492 13820 14544
rect 13872 14492 13878 14544
rect 14090 14464 14096 14476
rect 12084 14436 14096 14464
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16592 14464 16620 14572
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14600 18291 14603
rect 18598 14600 18604 14612
rect 18279 14572 18604 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 19518 14600 19524 14612
rect 18739 14572 19524 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 20533 14603 20591 14609
rect 20533 14569 20545 14603
rect 20579 14600 20591 14603
rect 20714 14600 20720 14612
rect 20579 14572 20720 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 22830 14560 22836 14612
rect 22888 14600 22894 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 22888 14572 25237 14600
rect 22888 14560 22894 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 25225 14563 25283 14569
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 19300 14504 20024 14532
rect 19300 14492 19306 14504
rect 16540 14436 16620 14464
rect 16761 14467 16819 14473
rect 16540 14424 16546 14436
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 17770 14464 17776 14476
rect 16807 14436 17776 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 19996 14473 20024 14504
rect 20346 14492 20352 14544
rect 20404 14532 20410 14544
rect 23382 14532 23388 14544
rect 20404 14504 23388 14532
rect 20404 14492 20410 14504
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 26142 14532 26148 14544
rect 23492 14504 26148 14532
rect 19889 14467 19947 14473
rect 19889 14464 19901 14467
rect 19852 14436 19901 14464
rect 19852 14424 19858 14436
rect 19889 14433 19901 14436
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 23492 14464 23520 14504
rect 26142 14492 26148 14504
rect 26200 14492 26206 14544
rect 20312 14436 23520 14464
rect 20312 14424 20318 14436
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23624 14436 23765 14464
rect 23624 14424 23630 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24486 14464 24492 14476
rect 23983 14436 24492 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 9539 14368 10180 14396
rect 10229 14399 10287 14405
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10318 14396 10324 14408
rect 10275 14368 10324 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 9674 14328 9680 14340
rect 2148 14300 9680 14328
rect 2148 14269 2176 14300
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 10704 14328 10732 14359
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12342 14396 12348 14408
rect 12124 14368 12348 14396
rect 12124 14356 12130 14368
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14396 12955 14399
rect 13538 14396 13544 14408
rect 12943 14368 13544 14396
rect 12943 14365 12955 14368
rect 12897 14359 12955 14365
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 19058 14356 19064 14408
rect 19116 14396 19122 14408
rect 20806 14396 20812 14408
rect 19116 14368 20812 14396
rect 19116 14356 19122 14368
rect 20806 14356 20812 14368
rect 20864 14396 20870 14408
rect 22002 14396 22008 14408
rect 20864 14368 22008 14396
rect 20864 14356 20870 14368
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 22112 14368 24593 14396
rect 10870 14328 10876 14340
rect 10704 14300 10876 14328
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 12268 14300 14964 14328
rect 2133 14263 2191 14269
rect 2133 14229 2145 14263
rect 2179 14229 2191 14263
rect 2133 14223 2191 14229
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 5258 14260 5264 14272
rect 3476 14232 5264 14260
rect 3476 14220 3482 14232
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5353 14263 5411 14269
rect 5353 14229 5365 14263
rect 5399 14260 5411 14263
rect 5442 14260 5448 14272
rect 5399 14232 5448 14260
rect 5399 14229 5411 14232
rect 5353 14223 5411 14229
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 7929 14263 7987 14269
rect 7929 14260 7941 14263
rect 7800 14232 7941 14260
rect 7800 14220 7806 14232
rect 7929 14229 7941 14232
rect 7975 14229 7987 14263
rect 7929 14223 7987 14229
rect 9033 14263 9091 14269
rect 9033 14229 9045 14263
rect 9079 14260 9091 14263
rect 9858 14260 9864 14272
rect 9079 14232 9864 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 12268 14260 12296 14300
rect 11204 14232 12296 14260
rect 11204 14220 11210 14232
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14550 14260 14556 14272
rect 13872 14232 14556 14260
rect 13872 14220 13878 14232
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 14936 14260 14964 14300
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 15856 14300 17172 14328
rect 15856 14260 15884 14300
rect 14936 14232 15884 14260
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16574 14260 16580 14272
rect 16071 14232 16580 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 17144 14260 17172 14300
rect 17218 14288 17224 14340
rect 17276 14288 17282 14340
rect 21358 14328 21364 14340
rect 18064 14300 21364 14328
rect 18064 14260 18092 14300
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 21634 14288 21640 14340
rect 21692 14328 21698 14340
rect 22112 14328 22140 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 21692 14300 22140 14328
rect 22925 14331 22983 14337
rect 21692 14288 21698 14300
rect 22925 14297 22937 14331
rect 22971 14328 22983 14331
rect 24026 14328 24032 14340
rect 22971 14300 24032 14328
rect 22971 14297 22983 14300
rect 22925 14291 22983 14297
rect 24026 14288 24032 14300
rect 24084 14328 24090 14340
rect 24210 14328 24216 14340
rect 24084 14300 24216 14328
rect 24084 14288 24090 14300
rect 24210 14288 24216 14300
rect 24268 14288 24274 14340
rect 17144 14232 18092 14260
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19392 14232 19441 14260
rect 19392 14220 19398 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 19794 14220 19800 14272
rect 19852 14220 19858 14272
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 22888 14232 23305 14260
rect 22888 14220 22894 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 23566 14220 23572 14272
rect 23624 14260 23630 14272
rect 23661 14263 23719 14269
rect 23661 14260 23673 14263
rect 23624 14232 23673 14260
rect 23624 14220 23630 14232
rect 23661 14229 23673 14232
rect 23707 14229 23719 14263
rect 23661 14223 23719 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 2148 13988 2176 14019
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2372 14028 2605 14056
rect 2372 14016 2378 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 4062 14056 4068 14068
rect 3283 14028 4068 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4798 14056 4804 14068
rect 4571 14028 4804 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 5184 13988 5212 14019
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 5592 14028 5641 14056
rect 5592 14016 5598 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6086 14056 6092 14068
rect 5951 14028 6092 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 7285 14059 7343 14065
rect 7285 14056 7297 14059
rect 6880 14028 7297 14056
rect 6880 14016 6886 14028
rect 7285 14025 7297 14028
rect 7331 14025 7343 14059
rect 7285 14019 7343 14025
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8536 14028 8769 14056
rect 8536 14016 8542 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 8757 14019 8815 14025
rect 9214 14016 9220 14068
rect 9272 14016 9278 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 10226 14056 10232 14068
rect 9447 14028 10232 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11011 14028 12204 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 7006 13988 7012 14000
rect 2148 13960 5120 13988
rect 5184 13960 7012 13988
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 2314 13920 2320 13932
rect 1903 13892 2320 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3418 13920 3424 13932
rect 3007 13892 3424 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13920 4123 13923
rect 4111 13892 5028 13920
rect 4111 13889 4123 13892
rect 4065 13883 4123 13889
rect 4154 13852 4160 13864
rect 3896 13824 4160 13852
rect 3896 13793 3924 13824
rect 4154 13812 4160 13824
rect 4212 13812 4218 13864
rect 3881 13787 3939 13793
rect 3881 13753 3893 13787
rect 3927 13753 3939 13787
rect 5000 13784 5028 13892
rect 5092 13852 5120 13960
rect 7006 13948 7012 13960
rect 7064 13948 7070 14000
rect 7650 13988 7656 14000
rect 7392 13960 7656 13988
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 6086 13920 6092 13932
rect 5399 13892 6092 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7098 13920 7104 13932
rect 6779 13892 7104 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7098 13880 7104 13892
rect 7156 13920 7162 13932
rect 7392 13920 7420 13960
rect 7650 13948 7656 13960
rect 7708 13948 7714 14000
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 10134 13988 10140 14000
rect 7984 13960 10140 13988
rect 7984 13948 7990 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10321 13991 10379 13997
rect 10321 13957 10333 13991
rect 10367 13988 10379 13991
rect 11701 13991 11759 13997
rect 10367 13960 11468 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 7156 13892 7420 13920
rect 7469 13923 7527 13929
rect 7156 13880 7162 13892
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7834 13920 7840 13932
rect 7515 13892 7840 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9079 13892 9873 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9861 13889 9873 13892
rect 9907 13920 9919 13923
rect 11054 13920 11060 13932
rect 9907 13892 11060 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 11146 13880 11152 13932
rect 11204 13880 11210 13932
rect 7558 13852 7564 13864
rect 5092 13824 7564 13852
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 11330 13852 11336 13864
rect 7668 13824 11336 13852
rect 7668 13784 7696 13824
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11440 13852 11468 13960
rect 11701 13957 11713 13991
rect 11747 13988 11759 13991
rect 12066 13988 12072 14000
rect 11747 13960 12072 13988
rect 11747 13957 11759 13960
rect 11701 13951 11759 13957
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 12176 13988 12204 14028
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 13265 14059 13323 14065
rect 13265 14056 13277 14059
rect 12308 14028 13277 14056
rect 12308 14016 12314 14028
rect 13265 14025 13277 14028
rect 13311 14025 13323 14059
rect 13265 14019 13323 14025
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14240 14028 15485 14056
rect 14240 14016 14246 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16264 14028 16681 14056
rect 16264 14016 16270 14028
rect 16669 14025 16681 14028
rect 16715 14056 16727 14059
rect 17218 14056 17224 14068
rect 16715 14028 17224 14056
rect 16715 14025 16727 14028
rect 16669 14019 16727 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 17920 14028 19334 14056
rect 17920 14016 17926 14028
rect 13630 13988 13636 14000
rect 12176 13960 13636 13988
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 14274 13988 14280 14000
rect 13740 13960 14280 13988
rect 11974 13880 11980 13932
rect 12032 13880 12038 13932
rect 12618 13880 12624 13932
rect 12676 13880 12682 13932
rect 13740 13929 13768 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 14550 13948 14556 14000
rect 14608 13948 14614 14000
rect 16022 13948 16028 14000
rect 16080 13988 16086 14000
rect 18233 13991 18291 13997
rect 16080 13960 18092 13988
rect 16080 13948 16086 13960
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 15286 13880 15292 13932
rect 15344 13920 15350 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 15344 13892 16129 13920
rect 15344 13880 15350 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 18064 13920 18092 13960
rect 18233 13957 18245 13991
rect 18279 13988 18291 13991
rect 18414 13988 18420 14000
rect 18279 13960 18420 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 18414 13948 18420 13960
rect 18472 13988 18478 14000
rect 19058 13988 19064 14000
rect 18472 13960 19064 13988
rect 18472 13948 18478 13960
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 19306 13988 19334 14028
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19484 14028 19533 14056
rect 19484 14016 19490 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20349 14059 20407 14065
rect 20349 14025 20361 14059
rect 20395 14056 20407 14059
rect 20806 14056 20812 14068
rect 20395 14028 20812 14056
rect 20395 14025 20407 14028
rect 20349 14019 20407 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 21140 14028 21189 14056
rect 21140 14016 21146 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 24670 14056 24676 14068
rect 21416 14028 24676 14056
rect 21416 14016 21422 14028
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 25038 14016 25044 14068
rect 25096 14056 25102 14068
rect 25590 14056 25596 14068
rect 25096 14028 25596 14056
rect 25096 14016 25102 14028
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 21450 13988 21456 14000
rect 19306 13960 21456 13988
rect 21450 13948 21456 13960
rect 21508 13988 21514 14000
rect 22097 13991 22155 13997
rect 22097 13988 22109 13991
rect 21508 13960 22109 13988
rect 21508 13948 21514 13960
rect 22097 13957 22109 13960
rect 22143 13957 22155 13991
rect 23382 13988 23388 14000
rect 22097 13951 22155 13957
rect 22204 13960 23388 13988
rect 20533 13923 20591 13929
rect 20533 13920 20545 13923
rect 18064 13892 20545 13920
rect 20533 13889 20545 13892
rect 20579 13920 20591 13923
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20579 13892 21097 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 22204 13920 22232 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 24946 13948 24952 14000
rect 25004 13988 25010 14000
rect 25133 13991 25191 13997
rect 25133 13988 25145 13991
rect 25004 13960 25145 13988
rect 25004 13948 25010 13960
rect 25133 13957 25145 13960
rect 25179 13988 25191 13991
rect 25866 13988 25872 14000
rect 25179 13960 25872 13988
rect 25179 13957 25191 13960
rect 25133 13951 25191 13957
rect 25866 13948 25872 13960
rect 25924 13948 25930 14000
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 21085 13883 21143 13889
rect 21192 13892 22232 13920
rect 22296 13892 22845 13920
rect 13538 13852 13544 13864
rect 11440 13824 13544 13852
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 16022 13852 16028 13864
rect 13832 13824 16028 13852
rect 5000 13756 7696 13784
rect 3881 13747 3939 13753
rect 7742 13744 7748 13796
rect 7800 13784 7806 13796
rect 7800 13756 11744 13784
rect 7800 13744 7806 13756
rect 1578 13676 1584 13728
rect 1636 13716 1642 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 1636 13688 6561 13716
rect 1636 13676 1642 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6549 13679 6607 13685
rect 9674 13676 9680 13728
rect 9732 13676 9738 13728
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11606 13716 11612 13728
rect 11112 13688 11612 13716
rect 11112 13676 11118 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11716 13716 11744 13756
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 13832 13784 13860 13824
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16264 13824 16313 13852
rect 16264 13812 16270 13824
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 16301 13815 16359 13821
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13821 17647 13855
rect 17589 13815 17647 13821
rect 11848 13756 13860 13784
rect 11848 13744 11854 13756
rect 17034 13744 17040 13796
rect 17092 13744 17098 13796
rect 17494 13744 17500 13796
rect 17552 13784 17558 13796
rect 17604 13784 17632 13815
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 21192 13852 21220 13892
rect 17920 13824 21220 13852
rect 21361 13855 21419 13861
rect 17920 13812 17926 13824
rect 21361 13821 21373 13855
rect 21407 13852 21419 13855
rect 21634 13852 21640 13864
rect 21407 13824 21640 13852
rect 21407 13821 21419 13824
rect 21361 13815 21419 13821
rect 21634 13812 21640 13824
rect 21692 13812 21698 13864
rect 22186 13812 22192 13864
rect 22244 13852 22250 13864
rect 22296 13852 22324 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 25958 13880 25964 13932
rect 26016 13880 26022 13932
rect 22244 13824 22324 13852
rect 23109 13855 23167 13861
rect 22244 13812 22250 13824
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 23155 13824 24440 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 22281 13787 22339 13793
rect 17552 13756 17632 13784
rect 17696 13756 20852 13784
rect 17552 13744 17558 13756
rect 12434 13716 12440 13728
rect 11716 13688 12440 13716
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 13988 13719 14046 13725
rect 13988 13685 14000 13719
rect 14034 13716 14046 13719
rect 15378 13716 15384 13728
rect 14034 13688 15384 13716
rect 14034 13685 14046 13688
rect 13988 13679 14046 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 16758 13676 16764 13728
rect 16816 13716 16822 13728
rect 17696 13716 17724 13756
rect 16816 13688 17724 13716
rect 16816 13676 16822 13688
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 19242 13716 19248 13728
rect 18564 13688 19248 13716
rect 18564 13676 18570 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 20824 13716 20852 13756
rect 22281 13753 22293 13787
rect 22327 13753 22339 13787
rect 24412 13784 24440 13824
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24544 13824 24593 13852
rect 24544 13812 24550 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 25317 13855 25375 13861
rect 25317 13821 25329 13855
rect 25363 13852 25375 13855
rect 25590 13852 25596 13864
rect 25363 13824 25596 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 25682 13812 25688 13864
rect 25740 13852 25746 13864
rect 25866 13852 25872 13864
rect 25740 13824 25872 13852
rect 25740 13812 25746 13824
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 24946 13784 24952 13796
rect 24412 13756 24952 13784
rect 22281 13747 22339 13753
rect 21726 13716 21732 13728
rect 20824 13688 21732 13716
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22296 13716 22324 13747
rect 24946 13744 24952 13756
rect 25004 13744 25010 13796
rect 22922 13716 22928 13728
rect 22296 13688 22928 13716
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 2593 13515 2651 13521
rect 2593 13481 2605 13515
rect 2639 13512 2651 13515
rect 3142 13512 3148 13524
rect 2639 13484 3148 13512
rect 2639 13481 2651 13484
rect 2593 13475 2651 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 3237 13515 3295 13521
rect 3237 13481 3249 13515
rect 3283 13512 3295 13515
rect 5902 13512 5908 13524
rect 3283 13484 5908 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 11790 13512 11796 13524
rect 9180 13484 11796 13512
rect 9180 13472 9186 13484
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 13541 13515 13599 13521
rect 11900 13484 13492 13512
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 5442 13444 5448 13456
rect 1627 13416 5448 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 5442 13404 5448 13416
rect 5500 13404 5506 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 11900 13444 11928 13484
rect 8352 13416 11928 13444
rect 13464 13444 13492 13484
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13998 13512 14004 13524
rect 13587 13484 14004 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15562 13512 15568 13524
rect 15252 13484 15568 13512
rect 15252 13472 15258 13484
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 17494 13512 17500 13524
rect 16080 13484 17500 13512
rect 16080 13472 16086 13484
rect 17494 13472 17500 13484
rect 17552 13512 17558 13524
rect 18233 13515 18291 13521
rect 18233 13512 18245 13515
rect 17552 13484 18245 13512
rect 17552 13472 17558 13484
rect 18233 13481 18245 13484
rect 18279 13481 18291 13515
rect 20162 13512 20168 13524
rect 18233 13475 18291 13481
rect 18432 13484 20168 13512
rect 13464 13416 14412 13444
rect 8352 13404 8358 13416
rect 2130 13336 2136 13388
rect 2188 13336 2194 13388
rect 9674 13376 9680 13388
rect 3344 13348 9680 13376
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13308 1823 13311
rect 2148 13308 2176 13336
rect 1811 13280 2176 13308
rect 2785 13311 2843 13317
rect 1811 13277 1823 13280
rect 1765 13271 1823 13277
rect 2785 13277 2797 13311
rect 2831 13308 2843 13311
rect 3344 13308 3372 13348
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 10928 13348 11805 13376
rect 10928 13336 10934 13348
rect 11793 13345 11805 13348
rect 11839 13345 11851 13379
rect 11793 13339 11851 13345
rect 13814 13336 13820 13388
rect 13872 13336 13878 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14384 13376 14412 13416
rect 14384 13348 15884 13376
rect 2831 13280 3372 13308
rect 2831 13277 2843 13280
rect 2785 13271 2843 13277
rect 2317 13243 2375 13249
rect 2317 13209 2329 13243
rect 2363 13240 2375 13243
rect 2792 13240 2820 13271
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 13832 13308 13860 13336
rect 4663 13280 11744 13308
rect 13202 13280 13860 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 2363 13212 2820 13240
rect 3973 13243 4031 13249
rect 2363 13209 2375 13212
rect 2317 13203 2375 13209
rect 3973 13209 3985 13243
rect 4019 13240 4031 13243
rect 9398 13240 9404 13252
rect 4019 13212 9404 13240
rect 4019 13209 4031 13212
rect 3973 13203 4031 13209
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 11606 13240 11612 13252
rect 9631 13212 11612 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 11606 13200 11612 13212
rect 11664 13200 11670 13252
rect 11716 13240 11744 13280
rect 11716 13212 11928 13240
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10870 13172 10876 13184
rect 10100 13144 10876 13172
rect 10100 13132 10106 13144
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11900 13172 11928 13212
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 13722 13200 13728 13252
rect 13780 13240 13786 13252
rect 14553 13243 14611 13249
rect 14553 13240 14565 13243
rect 13780 13212 14565 13240
rect 13780 13200 13786 13212
rect 14553 13209 14565 13212
rect 14599 13209 14611 13243
rect 14553 13203 14611 13209
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 15856 13240 15884 13348
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18322 13376 18328 13388
rect 16807 13348 18328 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18322 13336 18328 13348
rect 18380 13336 18386 13388
rect 16758 13240 16764 13252
rect 15856 13212 16764 13240
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17218 13200 17224 13252
rect 17276 13200 17282 13252
rect 15194 13172 15200 13184
rect 11900 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13132 15258 13184
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 16025 13175 16083 13181
rect 16025 13172 16037 13175
rect 15620 13144 16037 13172
rect 15620 13132 15626 13144
rect 16025 13141 16037 13144
rect 16071 13172 16083 13175
rect 18432 13172 18460 13484
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 21453 13515 21511 13521
rect 21453 13481 21465 13515
rect 21499 13512 21511 13515
rect 21634 13512 21640 13524
rect 21499 13484 21640 13512
rect 21499 13481 21511 13484
rect 21453 13475 21511 13481
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 23661 13515 23719 13521
rect 23661 13481 23673 13515
rect 23707 13512 23719 13515
rect 23934 13512 23940 13524
rect 23707 13484 23940 13512
rect 23707 13481 23719 13484
rect 23661 13475 23719 13481
rect 23934 13472 23940 13484
rect 23992 13472 23998 13524
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 24394 13512 24400 13524
rect 24176 13484 24400 13512
rect 24176 13472 24182 13484
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 24029 13447 24087 13453
rect 24029 13444 24041 13447
rect 23308 13416 24041 13444
rect 18693 13379 18751 13385
rect 18693 13345 18705 13379
rect 18739 13376 18751 13379
rect 18782 13376 18788 13388
rect 18739 13348 18788 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 21910 13376 21916 13388
rect 19720 13348 21916 13376
rect 19720 13320 19748 13348
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22646 13336 22652 13388
rect 22704 13376 22710 13388
rect 22922 13376 22928 13388
rect 22704 13348 22928 13376
rect 22704 13336 22710 13348
rect 22922 13336 22928 13348
rect 22980 13336 22986 13388
rect 19702 13268 19708 13320
rect 19760 13268 19766 13320
rect 23308 13294 23336 13416
rect 24029 13413 24041 13416
rect 24075 13444 24087 13447
rect 24210 13444 24216 13456
rect 24075 13416 24216 13444
rect 24075 13413 24087 13416
rect 24029 13407 24087 13413
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 23808 13348 25145 13376
rect 23808 13336 23814 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 25406 13308 25412 13320
rect 24136 13280 25412 13308
rect 19978 13200 19984 13252
rect 20036 13200 20042 13252
rect 21634 13240 21640 13252
rect 21206 13212 21640 13240
rect 16071 13144 18460 13172
rect 19337 13175 19395 13181
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 21284 13172 21312 13212
rect 21634 13200 21640 13212
rect 21692 13200 21698 13252
rect 22189 13243 22247 13249
rect 22189 13209 22201 13243
rect 22235 13209 22247 13243
rect 22189 13203 22247 13209
rect 19383 13144 21312 13172
rect 22204 13172 22232 13203
rect 24136 13172 24164 13280
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 24949 13243 25007 13249
rect 24949 13209 24961 13243
rect 24995 13240 25007 13243
rect 25866 13240 25872 13252
rect 24995 13212 25872 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 22204 13144 24164 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 24210 13132 24216 13184
rect 24268 13172 24274 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24268 13144 24593 13172
rect 24268 13132 24274 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 25041 13175 25099 13181
rect 25041 13141 25053 13175
rect 25087 13172 25099 13175
rect 25314 13172 25320 13184
rect 25087 13144 25320 13172
rect 25087 13141 25099 13144
rect 25041 13135 25099 13141
rect 25314 13132 25320 13144
rect 25372 13132 25378 13184
rect 25976 13172 26004 13880
rect 25884 13144 26004 13172
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12937 2007 12971
rect 1949 12931 2007 12937
rect 1964 12900 1992 12931
rect 2498 12928 2504 12980
rect 2556 12968 2562 12980
rect 2593 12971 2651 12977
rect 2593 12968 2605 12971
rect 2556 12940 2605 12968
rect 2556 12928 2562 12940
rect 2593 12937 2605 12940
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3200 12940 8432 12968
rect 3200 12928 3206 12940
rect 8294 12900 8300 12912
rect 1964 12872 8300 12900
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 8404 12900 8432 12940
rect 10594 12928 10600 12980
rect 10652 12928 10658 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11204 12940 11529 12968
rect 11204 12928 11210 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 12124 12940 12541 12968
rect 12124 12928 12130 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 12529 12931 12587 12937
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14274 12968 14280 12980
rect 13872 12940 14280 12968
rect 13872 12928 13878 12940
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15105 12971 15163 12977
rect 15105 12937 15117 12971
rect 15151 12968 15163 12971
rect 18414 12968 18420 12980
rect 15151 12940 18420 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 11238 12900 11244 12912
rect 8404 12872 11244 12900
rect 11238 12860 11244 12872
rect 11296 12860 11302 12912
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 11664 12872 13001 12900
rect 11664 12860 11670 12872
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 15120 12900 15148 12931
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 19521 12971 19579 12977
rect 19521 12968 19533 12971
rect 18656 12940 19533 12968
rect 18656 12928 18662 12940
rect 19521 12937 19533 12940
rect 19567 12937 19579 12971
rect 19521 12931 19579 12937
rect 19794 12928 19800 12980
rect 19852 12968 19858 12980
rect 19852 12940 19932 12968
rect 19852 12928 19858 12940
rect 13035 12872 15148 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 16301 12903 16359 12909
rect 16301 12900 16313 12903
rect 15436 12872 16313 12900
rect 15436 12860 15442 12872
rect 16301 12869 16313 12872
rect 16347 12869 16359 12903
rect 16301 12863 16359 12869
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 17218 12900 17224 12912
rect 16540 12872 17224 12900
rect 16540 12860 16546 12872
rect 17218 12860 17224 12872
rect 17276 12900 17282 12912
rect 19904 12900 19932 12940
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 20036 12940 24869 12968
rect 20036 12928 20042 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 24857 12931 24915 12937
rect 25130 12928 25136 12980
rect 25188 12968 25194 12980
rect 25314 12968 25320 12980
rect 25188 12940 25320 12968
rect 25188 12928 25194 12940
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 20717 12903 20775 12909
rect 20717 12900 20729 12903
rect 17276 12872 17618 12900
rect 18432 12872 19840 12900
rect 19904 12872 20729 12900
rect 17276 12860 17282 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2130 12832 2136 12844
rect 1719 12804 2136 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 7190 12832 7196 12844
rect 2823 12804 7196 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11698 12832 11704 12844
rect 11195 12804 11704 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 13446 12832 13452 12844
rect 12400 12804 13452 12832
rect 12400 12792 12406 12804
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 15068 12804 15301 12832
rect 15068 12792 15074 12804
rect 15289 12801 15301 12804
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 3191 12736 3249 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 3252 12696 3280 12727
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 12710 12764 12716 12776
rect 3476 12736 12716 12764
rect 3476 12724 3482 12736
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 17126 12724 17132 12776
rect 17184 12724 17190 12776
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 17678 12764 17684 12776
rect 17276 12736 17684 12764
rect 17276 12724 17282 12736
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 18432 12764 18460 12872
rect 18598 12792 18604 12844
rect 18656 12832 18662 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 18656 12804 19441 12832
rect 18656 12792 18662 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19812 12832 19840 12872
rect 20717 12869 20729 12872
rect 20763 12869 20775 12903
rect 22554 12900 22560 12912
rect 20717 12863 20775 12869
rect 21744 12872 22560 12900
rect 20530 12832 20536 12844
rect 19429 12795 19487 12801
rect 19536 12804 19748 12832
rect 19812 12804 20536 12832
rect 18156 12736 18460 12764
rect 11054 12696 11060 12708
rect 3252 12668 11060 12696
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 11698 12656 11704 12708
rect 11756 12696 11762 12708
rect 15746 12696 15752 12708
rect 11756 12668 15752 12696
rect 11756 12656 11762 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 10962 12588 10968 12640
rect 11020 12588 11026 12640
rect 15562 12588 15568 12640
rect 15620 12628 15626 12640
rect 18156 12628 18184 12736
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 19536 12764 19564 12804
rect 19300 12736 19564 12764
rect 19613 12767 19671 12773
rect 19300 12724 19306 12736
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19720 12764 19748 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 20622 12792 20628 12844
rect 20680 12792 20686 12844
rect 21744 12832 21772 12872
rect 22554 12860 22560 12872
rect 22612 12860 22618 12912
rect 23506 12872 24348 12900
rect 24320 12844 24348 12872
rect 20732 12804 21772 12832
rect 20732 12764 20760 12804
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 23934 12792 23940 12844
rect 23992 12832 23998 12844
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23992 12804 24225 12832
rect 23992 12792 23998 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24360 12804 25145 12832
rect 24360 12792 24366 12804
rect 25133 12801 25145 12804
rect 25179 12832 25191 12835
rect 25317 12835 25375 12841
rect 25317 12832 25329 12835
rect 25179 12804 25329 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 25317 12801 25329 12804
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 19720 12736 20760 12764
rect 20809 12767 20867 12773
rect 19613 12727 19671 12733
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 18601 12699 18659 12705
rect 18601 12696 18613 12699
rect 18472 12668 18613 12696
rect 18472 12656 18478 12668
rect 18601 12665 18613 12668
rect 18647 12696 18659 12699
rect 19628 12696 19656 12727
rect 18647 12668 19656 12696
rect 18647 12665 18659 12668
rect 18601 12659 18659 12665
rect 20530 12656 20536 12708
rect 20588 12696 20594 12708
rect 20824 12696 20852 12727
rect 20990 12724 20996 12776
rect 21048 12764 21054 12776
rect 21358 12764 21364 12776
rect 21048 12736 21364 12764
rect 21048 12724 21054 12736
rect 21358 12724 21364 12736
rect 21416 12724 21422 12776
rect 21450 12724 21456 12776
rect 21508 12764 21514 12776
rect 21545 12767 21603 12773
rect 21545 12764 21557 12767
rect 21508 12736 21557 12764
rect 21508 12724 21514 12736
rect 21545 12733 21557 12736
rect 21591 12733 21603 12767
rect 21545 12727 21603 12733
rect 22278 12724 22284 12776
rect 22336 12724 22342 12776
rect 23750 12724 23756 12776
rect 23808 12724 23814 12776
rect 20588 12668 20852 12696
rect 20588 12656 20594 12668
rect 23382 12656 23388 12708
rect 23440 12696 23446 12708
rect 23842 12696 23848 12708
rect 23440 12668 23848 12696
rect 23440 12656 23446 12668
rect 23842 12656 23848 12668
rect 23900 12656 23906 12708
rect 15620 12600 18184 12628
rect 15620 12588 15626 12600
rect 19058 12588 19064 12640
rect 19116 12588 19122 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 20257 12631 20315 12637
rect 20257 12628 20269 12631
rect 19576 12600 20269 12628
rect 19576 12588 19582 12600
rect 20257 12597 20269 12600
rect 20303 12597 20315 12631
rect 20257 12591 20315 12597
rect 21361 12631 21419 12637
rect 21361 12597 21373 12631
rect 21407 12628 21419 12631
rect 21634 12628 21640 12640
rect 21407 12600 21640 12628
rect 21407 12597 21419 12600
rect 21361 12591 21419 12597
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22646 12628 22652 12640
rect 22152 12600 22652 12628
rect 22152 12588 22158 12600
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 23014 12588 23020 12640
rect 23072 12628 23078 12640
rect 23934 12628 23940 12640
rect 23072 12600 23940 12628
rect 23072 12588 23078 12600
rect 23934 12588 23940 12600
rect 23992 12588 23998 12640
rect 25682 12588 25688 12640
rect 25740 12628 25746 12640
rect 25884 12628 25912 13144
rect 25740 12600 25912 12628
rect 25740 12588 25746 12600
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 11517 12427 11575 12433
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 11606 12424 11612 12436
rect 11563 12396 11612 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11698 12384 11704 12436
rect 11756 12384 11762 12436
rect 11808 12396 12434 12424
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 11808 12356 11836 12396
rect 6972 12328 11836 12356
rect 12406 12356 12434 12396
rect 13722 12384 13728 12436
rect 13780 12384 13786 12436
rect 13832 12396 20760 12424
rect 13832 12356 13860 12396
rect 12406 12328 13860 12356
rect 6972 12316 6978 12328
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18601 12359 18659 12365
rect 18601 12356 18613 12359
rect 18288 12328 18613 12356
rect 18288 12316 18294 12328
rect 18601 12325 18613 12328
rect 18647 12325 18659 12359
rect 20732 12356 20760 12396
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 23290 12424 23296 12436
rect 21048 12396 23296 12424
rect 21048 12384 21054 12396
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 25225 12427 25283 12433
rect 25225 12393 25237 12427
rect 25271 12424 25283 12427
rect 25314 12424 25320 12436
rect 25271 12396 25320 12424
rect 25271 12393 25283 12396
rect 25225 12387 25283 12393
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 21818 12356 21824 12368
rect 18601 12319 18659 12325
rect 18708 12328 19564 12356
rect 20732 12328 21824 12356
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 7524 12260 15393 12288
rect 7524 12248 7530 12260
rect 15381 12257 15393 12260
rect 15427 12288 15439 12291
rect 15470 12288 15476 12300
rect 15427 12260 15476 12288
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16758 12288 16764 12300
rect 15795 12260 16764 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 18708 12288 18736 12328
rect 17736 12260 18736 12288
rect 17736 12248 17742 12260
rect 19426 12248 19432 12300
rect 19484 12248 19490 12300
rect 19536 12288 19564 12328
rect 21818 12316 21824 12328
rect 21876 12316 21882 12368
rect 19536 12260 21036 12288
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11940 12192 11989 12220
rect 11940 12180 11946 12192
rect 11977 12189 11989 12192
rect 12023 12220 12035 12223
rect 12342 12220 12348 12232
rect 12023 12192 12348 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12220 13139 12223
rect 13354 12220 13360 12232
rect 13127 12192 13360 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 13722 12220 13728 12232
rect 13412 12192 13728 12220
rect 13412 12180 13418 12192
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14056 12192 14289 12220
rect 14056 12180 14062 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18506 12220 18512 12232
rect 18003 12192 18512 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 14458 12152 14464 12164
rect 12636 12124 14464 12152
rect 1946 12044 1952 12096
rect 2004 12044 2010 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 12526 12084 12532 12096
rect 9916 12056 12532 12084
rect 9916 12044 9922 12056
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12636 12093 12664 12124
rect 14458 12112 14464 12124
rect 14516 12112 14522 12164
rect 15289 12155 15347 12161
rect 15289 12121 15301 12155
rect 15335 12152 15347 12155
rect 15470 12152 15476 12164
rect 15335 12124 15476 12152
rect 15335 12121 15347 12124
rect 15289 12115 15347 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16298 12152 16304 12164
rect 16071 12124 16304 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16298 12112 16304 12124
rect 16356 12112 16362 12164
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 18877 12155 18935 12161
rect 18877 12152 18889 12155
rect 17920 12124 18889 12152
rect 17920 12112 17926 12124
rect 18877 12121 18889 12124
rect 18923 12121 18935 12155
rect 18877 12115 18935 12121
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12152 19763 12155
rect 19978 12152 19984 12164
rect 19751 12124 19984 12152
rect 19751 12121 19763 12124
rect 19705 12115 19763 12121
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20438 12112 20444 12164
rect 20496 12112 20502 12164
rect 21008 12152 21036 12260
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21910 12288 21916 12300
rect 21416 12260 21916 12288
rect 21416 12248 21422 12260
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 22603 12260 25268 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 25240 12232 25268 12260
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21637 12223 21695 12229
rect 21637 12220 21649 12223
rect 21140 12192 21649 12220
rect 21140 12180 21146 12192
rect 21637 12189 21649 12192
rect 21683 12189 21695 12223
rect 21637 12183 21695 12189
rect 24118 12180 24124 12232
rect 24176 12220 24182 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24176 12192 24593 12220
rect 24176 12180 24182 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 25222 12180 25228 12232
rect 25280 12180 25286 12232
rect 23842 12152 23848 12164
rect 21008 12124 22094 12152
rect 23782 12124 23848 12152
rect 12621 12087 12679 12093
rect 12621 12053 12633 12087
rect 12667 12053 12679 12087
rect 12621 12047 12679 12053
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 13136 12056 14933 12084
rect 13136 12044 13142 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 17368 12056 17509 12084
rect 17368 12044 17374 12056
rect 17497 12053 17509 12056
rect 17543 12084 17555 12087
rect 17586 12084 17592 12096
rect 17543 12056 17592 12084
rect 17543 12053 17555 12056
rect 17497 12047 17555 12053
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 19058 12084 19064 12096
rect 18564 12056 19064 12084
rect 18564 12044 18570 12056
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 20070 12084 20076 12096
rect 19484 12056 20076 12084
rect 19484 12044 19490 12056
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20588 12056 21189 12084
rect 20588 12044 20594 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 22066 12084 22094 12124
rect 23842 12112 23848 12124
rect 23900 12152 23906 12164
rect 24302 12152 24308 12164
rect 23900 12124 24308 12152
rect 23900 12112 23906 12124
rect 24302 12112 24308 12124
rect 24360 12112 24366 12164
rect 22646 12084 22652 12096
rect 22066 12056 22652 12084
rect 21177 12047 21235 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 23934 12084 23940 12096
rect 23440 12056 23940 12084
rect 23440 12044 23446 12056
rect 23934 12044 23940 12056
rect 23992 12084 23998 12096
rect 24029 12087 24087 12093
rect 24029 12084 24041 12087
rect 23992 12056 24041 12084
rect 23992 12044 23998 12056
rect 24029 12053 24041 12056
rect 24075 12053 24087 12087
rect 24029 12047 24087 12053
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 11882 11840 11888 11892
rect 11940 11840 11946 11892
rect 12250 11840 12256 11892
rect 12308 11840 12314 11892
rect 13814 11880 13820 11892
rect 12820 11852 13820 11880
rect 12820 11753 12848 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 16761 11883 16819 11889
rect 16761 11880 16773 11883
rect 16540 11852 16773 11880
rect 16540 11840 16546 11852
rect 16761 11849 16773 11852
rect 16807 11849 16819 11883
rect 16761 11843 16819 11849
rect 18877 11883 18935 11889
rect 18877 11849 18889 11883
rect 18923 11880 18935 11883
rect 19426 11880 19432 11892
rect 18923 11852 19432 11880
rect 18923 11849 18935 11852
rect 18877 11843 18935 11849
rect 13078 11772 13084 11824
rect 13136 11772 13142 11824
rect 15010 11812 15016 11824
rect 14306 11784 15016 11812
rect 15010 11772 15016 11784
rect 15068 11772 15074 11824
rect 16776 11812 16804 11843
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20496 11852 21036 11880
rect 20496 11840 20502 11852
rect 17862 11812 17868 11824
rect 16776 11784 17868 11812
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11676 12587 11679
rect 13538 11676 13544 11688
rect 12575 11648 13544 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 13780 11648 14565 11676
rect 13780 11636 13786 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15102 11676 15108 11688
rect 15059 11648 15108 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 16390 11676 16396 11688
rect 15335 11648 16396 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 16868 11676 16896 11784
rect 17862 11772 17868 11784
rect 17920 11772 17926 11824
rect 19702 11812 19708 11824
rect 19444 11784 19708 11812
rect 19444 11753 19472 11784
rect 19702 11772 19708 11784
rect 19760 11772 19766 11824
rect 21008 11812 21036 11852
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 26234 11880 26240 11892
rect 22152 11852 26240 11880
rect 22152 11840 22158 11852
rect 26234 11840 26240 11852
rect 26292 11840 26298 11892
rect 21634 11812 21640 11824
rect 20930 11784 21640 11812
rect 21634 11772 21640 11784
rect 21692 11772 21698 11824
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25130 11772 25136 11824
rect 25188 11772 25194 11824
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 23937 11747 23995 11753
rect 23937 11713 23949 11747
rect 23983 11713 23995 11747
rect 23937 11707 23995 11713
rect 16942 11676 16948 11688
rect 16868 11648 16948 11676
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 19058 11676 19064 11688
rect 17451 11648 19064 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 16301 11611 16359 11617
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 16482 11608 16488 11620
rect 16347 11580 16488 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 17144 11608 17172 11639
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 21174 11676 21180 11688
rect 19751 11648 21180 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 22738 11676 22744 11688
rect 21284 11648 22744 11676
rect 21284 11608 21312 11648
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 16632 11580 17172 11608
rect 21008 11580 21312 11608
rect 16632 11568 16638 11580
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 21008 11540 21036 11580
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 23952 11608 23980 11707
rect 21876 11580 23980 11608
rect 21876 11568 21882 11580
rect 18932 11512 21036 11540
rect 18932 11500 18938 11512
rect 21082 11500 21088 11552
rect 21140 11540 21146 11552
rect 21177 11543 21235 11549
rect 21177 11540 21189 11543
rect 21140 11512 21189 11540
rect 21140 11500 21146 11512
rect 21177 11509 21189 11512
rect 21223 11509 21235 11543
rect 21177 11503 21235 11509
rect 21634 11500 21640 11552
rect 21692 11500 21698 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 22094 11336 22100 11348
rect 4488 11308 22100 11336
rect 4488 11296 4494 11308
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 22281 11339 22339 11345
rect 22281 11305 22293 11339
rect 22327 11336 22339 11339
rect 22646 11336 22652 11348
rect 22327 11308 22652 11336
rect 22327 11305 22339 11308
rect 22281 11299 22339 11305
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12492 11240 13185 11268
rect 12492 11228 12498 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 14185 11271 14243 11277
rect 14185 11237 14197 11271
rect 14231 11268 14243 11271
rect 14366 11268 14372 11280
rect 14231 11240 14372 11268
rect 14231 11237 14243 11240
rect 14185 11231 14243 11237
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 15286 11268 15292 11280
rect 14507 11240 15292 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 15378 11228 15384 11280
rect 15436 11228 15442 11280
rect 16298 11228 16304 11280
rect 16356 11228 16362 11280
rect 16669 11271 16727 11277
rect 16669 11237 16681 11271
rect 16715 11268 16727 11271
rect 17218 11268 17224 11280
rect 16715 11240 17224 11268
rect 16715 11237 16727 11240
rect 16669 11231 16727 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 17957 11271 18015 11277
rect 17957 11237 17969 11271
rect 18003 11268 18015 11271
rect 18322 11268 18328 11280
rect 18003 11240 18328 11268
rect 18003 11237 18015 11240
rect 17957 11231 18015 11237
rect 18322 11228 18328 11240
rect 18380 11228 18386 11280
rect 18432 11240 18828 11268
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 18432 11200 18460 11240
rect 12584 11172 18460 11200
rect 12584 11160 12590 11172
rect 18690 11160 18696 11212
rect 18748 11160 18754 11212
rect 18800 11200 18828 11240
rect 19978 11228 19984 11280
rect 20036 11268 20042 11280
rect 20073 11271 20131 11277
rect 20073 11268 20085 11271
rect 20036 11240 20085 11268
rect 20036 11228 20042 11240
rect 20073 11237 20085 11240
rect 20119 11237 20131 11271
rect 20073 11231 20131 11237
rect 21174 11228 21180 11280
rect 21232 11228 21238 11280
rect 21634 11228 21640 11280
rect 21692 11268 21698 11280
rect 22296 11268 22324 11299
rect 22646 11296 22652 11308
rect 22704 11336 22710 11348
rect 23842 11336 23848 11348
rect 22704 11308 23848 11336
rect 22704 11296 22710 11308
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 25038 11296 25044 11348
rect 25096 11336 25102 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 25096 11308 25237 11336
rect 25096 11296 25102 11308
rect 25225 11305 25237 11308
rect 25271 11305 25283 11339
rect 25225 11299 25283 11305
rect 21692 11240 22324 11268
rect 21692 11228 21698 11240
rect 20254 11200 20260 11212
rect 18800 11172 20260 11200
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20990 11200 20996 11212
rect 20864 11172 20996 11200
rect 20864 11160 20870 11172
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24854 11200 24860 11212
rect 23891 11172 24860 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11132 14703 11135
rect 15657 11135 15715 11141
rect 14691 11104 15240 11132
rect 14691 11101 14703 11104
rect 14645 11095 14703 11101
rect 15212 11073 15240 11104
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 16022 11132 16028 11144
rect 15703 11104 16028 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16758 11092 16764 11144
rect 16816 11092 16822 11144
rect 16942 11092 16948 11144
rect 17000 11092 17006 11144
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 18708 11132 18736 11160
rect 17359 11104 18736 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 20036 11104 20484 11132
rect 20036 11092 20042 11104
rect 15197 11067 15255 11073
rect 13556 11036 15148 11064
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 11698 10996 11704 11008
rect 4120 10968 11704 10996
rect 4120 10956 4126 10968
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 13556 11005 13584 11036
rect 13541 10999 13599 11005
rect 13541 10965 13553 10999
rect 13587 10965 13599 10999
rect 13541 10959 13599 10965
rect 14918 10956 14924 11008
rect 14976 10956 14982 11008
rect 15120 10996 15148 11036
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 17678 11064 17684 11076
rect 15243 11036 17684 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18380 11036 18705 11064
rect 18380 11024 18386 11036
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 18693 11027 18751 11033
rect 18877 11067 18935 11073
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 20070 11064 20076 11076
rect 18923 11036 20076 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 20456 11064 20484 11104
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 22738 11092 22744 11144
rect 22796 11092 22802 11144
rect 24578 11092 24584 11144
rect 24636 11092 24642 11144
rect 21818 11064 21824 11076
rect 20456 11036 21824 11064
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 21910 11024 21916 11076
rect 21968 11024 21974 11076
rect 23382 11064 23388 11076
rect 22066 11036 23388 11064
rect 16574 10996 16580 11008
rect 15120 10968 16580 10996
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 19702 10956 19708 11008
rect 19760 10996 19766 11008
rect 22066 10996 22094 11036
rect 23382 11024 23388 11036
rect 23440 11024 23446 11076
rect 19760 10968 22094 10996
rect 19760 10956 19766 10968
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 13630 10752 13636 10804
rect 13688 10752 13694 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13872 10764 13921 10792
rect 13872 10752 13878 10764
rect 13909 10761 13921 10764
rect 13955 10792 13967 10795
rect 14918 10792 14924 10804
rect 13955 10764 14924 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 16666 10792 16672 10804
rect 16163 10764 16672 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 16666 10752 16672 10764
rect 16724 10752 16730 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 16850 10792 16856 10804
rect 16807 10764 16856 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 17126 10752 17132 10804
rect 17184 10792 17190 10804
rect 17957 10795 18015 10801
rect 17957 10792 17969 10795
rect 17184 10764 17969 10792
rect 17184 10752 17190 10764
rect 17957 10761 17969 10764
rect 18003 10761 18015 10795
rect 17957 10755 18015 10761
rect 19058 10752 19064 10804
rect 19116 10752 19122 10804
rect 20349 10795 20407 10801
rect 20349 10761 20361 10795
rect 20395 10792 20407 10795
rect 22278 10792 22284 10804
rect 20395 10764 22284 10792
rect 20395 10761 20407 10764
rect 20349 10755 20407 10761
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 23293 10727 23351 10733
rect 11756 10696 15056 10724
rect 11756 10684 11762 10696
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 14384 10520 14412 10619
rect 14458 10548 14464 10600
rect 14516 10588 14522 10600
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14516 10560 14841 10588
rect 14516 10548 14522 10560
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 15028 10588 15056 10696
rect 15120 10696 23060 10724
rect 15120 10665 15148 10696
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16850 10656 16856 10668
rect 16347 10628 16856 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 18414 10616 18420 10668
rect 18472 10616 18478 10668
rect 19702 10616 19708 10668
rect 19760 10616 19766 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 18322 10588 18328 10600
rect 15028 10560 18328 10588
rect 14829 10551 14887 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 20824 10588 20852 10619
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 21542 10616 21548 10668
rect 21600 10656 21606 10668
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 21600 10628 22109 10656
rect 21600 10616 21606 10628
rect 22097 10625 22109 10628
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22554 10656 22560 10668
rect 22336 10628 22560 10656
rect 22336 10616 22342 10628
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 23032 10656 23060 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23032 10628 23949 10656
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 22370 10588 22376 10600
rect 18432 10560 19840 10588
rect 20824 10560 22376 10588
rect 18432 10532 18460 10560
rect 15562 10520 15568 10532
rect 14384 10492 15568 10520
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 16482 10480 16488 10532
rect 16540 10520 16546 10532
rect 16540 10492 18368 10520
rect 16540 10480 16546 10492
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 16942 10452 16948 10464
rect 14231 10424 16948 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 17126 10452 17132 10464
rect 17083 10424 17132 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 18340 10452 18368 10492
rect 18414 10480 18420 10532
rect 18472 10480 18478 10532
rect 19058 10480 19064 10532
rect 19116 10480 19122 10532
rect 19334 10480 19340 10532
rect 19392 10520 19398 10532
rect 19702 10520 19708 10532
rect 19392 10492 19708 10520
rect 19392 10480 19398 10492
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 19812 10520 19840 10560
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 22002 10520 22008 10532
rect 19812 10492 22008 10520
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 26510 10520 26516 10532
rect 22480 10492 26516 10520
rect 19076 10452 19104 10480
rect 18340 10424 19104 10452
rect 19429 10455 19487 10461
rect 19429 10421 19441 10455
rect 19475 10452 19487 10455
rect 20162 10452 20168 10464
rect 19475 10424 20168 10452
rect 19475 10421 19487 10424
rect 19429 10415 19487 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 22480 10452 22508 10492
rect 26510 10480 26516 10492
rect 26568 10480 26574 10532
rect 20312 10424 22508 10452
rect 20312 10412 20318 10424
rect 22554 10412 22560 10464
rect 22612 10452 22618 10464
rect 23290 10452 23296 10464
rect 22612 10424 23296 10452
rect 22612 10412 22618 10424
rect 23290 10412 23296 10424
rect 23348 10412 23354 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 14458 10208 14464 10260
rect 14516 10208 14522 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14884 10220 15117 10248
rect 14884 10208 14890 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15252 10220 15761 10248
rect 15252 10208 15258 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 17037 10251 17095 10257
rect 17037 10217 17049 10251
rect 17083 10248 17095 10251
rect 17218 10248 17224 10260
rect 17083 10220 17224 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 18414 10248 18420 10260
rect 17644 10220 18420 10248
rect 17644 10208 17650 10220
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 18693 10251 18751 10257
rect 18693 10217 18705 10251
rect 18739 10248 18751 10251
rect 19610 10248 19616 10260
rect 18739 10220 19616 10248
rect 18739 10217 18751 10220
rect 18693 10211 18751 10217
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 22370 10248 22376 10260
rect 20947 10220 22376 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 22370 10208 22376 10220
rect 22428 10208 22434 10260
rect 12406 10152 21496 10180
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 12406 10112 12434 10152
rect 11020 10084 12434 10112
rect 11020 10072 11026 10084
rect 16390 10072 16396 10124
rect 16448 10112 16454 10124
rect 16448 10084 17356 10112
rect 16448 10072 16454 10084
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16482 10044 16488 10056
rect 15979 10016 16488 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16666 10044 16672 10056
rect 16623 10016 16672 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17126 10004 17132 10056
rect 17184 10044 17190 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 17184 10016 17233 10044
rect 17184 10004 17190 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17328 10044 17356 10084
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17460 10084 17969 10112
rect 17460 10072 17466 10084
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 19613 10115 19671 10121
rect 19613 10081 19625 10115
rect 19659 10112 19671 10115
rect 20990 10112 20996 10124
rect 19659 10084 20996 10112
rect 19659 10081 19671 10084
rect 19613 10075 19671 10081
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21468 10112 21496 10152
rect 23198 10140 23204 10192
rect 23256 10180 23262 10192
rect 23256 10152 25176 10180
rect 23256 10140 23262 10152
rect 25148 10121 25176 10152
rect 25133 10115 25191 10121
rect 21468 10084 23888 10112
rect 18877 10047 18935 10053
rect 17328 10016 18828 10044
rect 17221 10007 17279 10013
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 16393 9911 16451 9917
rect 16393 9908 16405 9911
rect 12860 9880 16405 9908
rect 12860 9868 12866 9880
rect 16393 9877 16405 9880
rect 16439 9877 16451 9911
rect 16393 9871 16451 9877
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17586 9908 17592 9920
rect 16724 9880 17592 9908
rect 16724 9868 16730 9880
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 18800 9908 18828 10016
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 18923 10016 19380 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19352 9985 19380 10016
rect 20254 10004 20260 10056
rect 20312 10004 20318 10056
rect 23860 10053 23888 10084
rect 25133 10081 25145 10115
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25774 10044 25780 10056
rect 25087 10016 25780 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25774 10004 25780 10016
rect 25832 10004 25838 10056
rect 19337 9979 19395 9985
rect 19337 9945 19349 9979
rect 19383 9976 19395 9979
rect 20346 9976 20352 9988
rect 19383 9948 20352 9976
rect 19383 9945 19395 9948
rect 19337 9939 19395 9945
rect 20346 9936 20352 9948
rect 20404 9936 20410 9988
rect 21634 9936 21640 9988
rect 21692 9936 21698 9988
rect 22646 9936 22652 9988
rect 22704 9936 22710 9988
rect 23382 9936 23388 9988
rect 23440 9976 23446 9988
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 23440 9948 24961 9976
rect 23440 9936 23446 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 21542 9908 21548 9920
rect 18800 9880 21548 9908
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 23109 9911 23167 9917
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23198 9908 23204 9920
rect 23155 9880 23204 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 23934 9868 23940 9920
rect 23992 9868 23998 9920
rect 24578 9868 24584 9920
rect 24636 9868 24642 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 14642 9664 14648 9716
rect 14700 9704 14706 9716
rect 14737 9707 14795 9713
rect 14737 9704 14749 9707
rect 14700 9676 14749 9704
rect 14700 9664 14706 9676
rect 14737 9673 14749 9676
rect 14783 9673 14795 9707
rect 14737 9667 14795 9673
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15381 9707 15439 9713
rect 15381 9704 15393 9707
rect 15344 9676 15393 9704
rect 15344 9664 15350 9676
rect 15381 9673 15393 9676
rect 15427 9673 15439 9707
rect 15381 9667 15439 9673
rect 16942 9664 16948 9716
rect 17000 9704 17006 9716
rect 19610 9704 19616 9716
rect 17000 9676 19616 9704
rect 17000 9664 17006 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20220 9676 21036 9704
rect 20220 9664 20226 9676
rect 15654 9596 15660 9648
rect 15712 9596 15718 9648
rect 18141 9639 18199 9645
rect 18141 9605 18153 9639
rect 18187 9636 18199 9639
rect 18598 9636 18604 9648
rect 18187 9608 18604 9636
rect 18187 9605 18199 9608
rect 18141 9599 18199 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 20898 9636 20904 9648
rect 18984 9608 20904 9636
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 16298 9568 16304 9580
rect 15887 9540 16304 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 18984 9577 19012 9608
rect 20898 9596 20904 9608
rect 20956 9596 20962 9648
rect 21008 9636 21036 9676
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 22646 9704 22652 9716
rect 22152 9676 22652 9704
rect 22152 9664 22158 9676
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 21082 9636 21088 9648
rect 21008 9608 21088 9636
rect 21082 9596 21088 9608
rect 21140 9636 21146 9648
rect 22002 9636 22008 9648
rect 21140 9608 22008 9636
rect 21140 9596 21146 9608
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23842 9636 23848 9648
rect 23532 9608 23848 9636
rect 23532 9596 23538 9608
rect 23842 9596 23848 9608
rect 23900 9596 23906 9648
rect 25130 9596 25136 9648
rect 25188 9596 25194 9648
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9568 19671 9571
rect 20346 9568 20352 9580
rect 19659 9540 20352 9568
rect 19659 9537 19671 9540
rect 19613 9531 19671 9537
rect 17696 9500 17724 9531
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 20717 9572 20775 9577
rect 20717 9571 20852 9572
rect 20717 9537 20729 9571
rect 20763 9568 20852 9571
rect 20763 9544 21128 9568
rect 20763 9537 20775 9544
rect 20824 9540 21128 9544
rect 20717 9531 20775 9537
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 17696 9472 19993 9500
rect 19981 9469 19993 9472
rect 20027 9500 20039 9503
rect 21100 9500 21128 9540
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21232 9540 21373 9568
rect 21232 9528 21238 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 21542 9528 21548 9580
rect 21600 9568 21606 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 21600 9540 22109 9568
rect 21600 9528 21606 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22462 9528 22468 9580
rect 22520 9568 22526 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 22520 9540 23949 9568
rect 22520 9528 22526 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 21726 9500 21732 9512
rect 20027 9472 20668 9500
rect 21100 9472 21732 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 15068 9404 16129 9432
rect 15068 9392 15074 9404
rect 16117 9401 16129 9404
rect 16163 9401 16175 9435
rect 16117 9395 16175 9401
rect 18782 9392 18788 9444
rect 18840 9392 18846 9444
rect 19429 9435 19487 9441
rect 19429 9401 19441 9435
rect 19475 9432 19487 9435
rect 19794 9432 19800 9444
rect 19475 9404 19800 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 20530 9392 20536 9444
rect 20588 9392 20594 9444
rect 20640 9432 20668 9472
rect 21726 9460 21732 9472
rect 21784 9500 21790 9512
rect 24026 9500 24032 9512
rect 21784 9472 24032 9500
rect 21784 9460 21790 9472
rect 24026 9460 24032 9472
rect 24084 9460 24090 9512
rect 22002 9432 22008 9444
rect 20640 9404 22008 9432
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 26878 9432 26884 9444
rect 22152 9404 26884 9432
rect 22152 9392 22158 9404
rect 26878 9392 26884 9404
rect 26936 9392 26942 9444
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 19334 9364 19340 9376
rect 17543 9336 19340 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 21177 9367 21235 9373
rect 21177 9333 21189 9367
rect 21223 9364 21235 9367
rect 22370 9364 22376 9376
rect 21223 9336 22376 9364
rect 21223 9333 21235 9336
rect 21177 9327 21235 9333
rect 22370 9324 22376 9336
rect 22428 9324 22434 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 25958 9188 25964 9240
rect 26016 9228 26022 9240
rect 26602 9228 26608 9240
rect 26016 9200 26608 9228
rect 26016 9188 26022 9200
rect 26602 9188 26608 9200
rect 26660 9188 26666 9240
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 11882 9160 11888 9172
rect 11839 9132 11888 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 15838 9120 15844 9172
rect 15896 9160 15902 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 15896 9132 18061 9160
rect 15896 9120 15902 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 19150 9160 19156 9172
rect 18049 9123 18107 9129
rect 18616 9132 19156 9160
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8628 9064 10180 9092
rect 8628 9052 8634 9064
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10152 9024 10180 9064
rect 16117 9027 16175 9033
rect 16117 9024 16129 9027
rect 10152 8996 16129 9024
rect 16117 8993 16129 8996
rect 16163 8993 16175 9027
rect 16117 8987 16175 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 8993 16451 9027
rect 18616 9024 18644 9132
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19429 9163 19487 9169
rect 19429 9129 19441 9163
rect 19475 9160 19487 9163
rect 21542 9160 21548 9172
rect 19475 9132 21548 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 22097 9163 22155 9169
rect 22097 9160 22109 9163
rect 21692 9132 22109 9160
rect 21692 9120 21698 9132
rect 22097 9129 22109 9132
rect 22143 9129 22155 9163
rect 22097 9123 22155 9129
rect 25225 9163 25283 9169
rect 25225 9129 25237 9163
rect 25271 9160 25283 9163
rect 25406 9160 25412 9172
rect 25271 9132 25412 9160
rect 25271 9129 25283 9132
rect 25225 9123 25283 9129
rect 25406 9120 25412 9132
rect 25464 9120 25470 9172
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 20073 9095 20131 9101
rect 20073 9092 20085 9095
rect 18748 9064 20085 9092
rect 18748 9052 18754 9064
rect 20073 9061 20085 9064
rect 20119 9061 20131 9095
rect 20073 9055 20131 9061
rect 20162 9024 20168 9036
rect 16393 8987 16451 8993
rect 17604 8996 18644 9024
rect 18800 8996 20168 9024
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 6880 8860 10333 8888
rect 6880 8848 6886 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12161 8891 12219 8897
rect 12161 8888 12173 8891
rect 11546 8860 12173 8888
rect 10321 8851 10379 8857
rect 12161 8857 12173 8860
rect 12207 8888 12219 8891
rect 13814 8888 13820 8900
rect 12207 8860 13820 8888
rect 12207 8857 12219 8860
rect 12161 8851 12219 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 16408 8888 16436 8987
rect 17604 8965 17632 8996
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18800 8956 18828 8996
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 22830 9024 22836 9036
rect 21376 8996 22836 9024
rect 18279 8928 18828 8956
rect 18877 8959 18935 8965
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 19426 8956 19432 8968
rect 18923 8928 19432 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19610 8916 19616 8968
rect 19668 8916 19674 8968
rect 20257 8959 20315 8965
rect 20257 8925 20269 8959
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 19978 8888 19984 8900
rect 16408 8860 19984 8888
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 20272 8888 20300 8919
rect 20806 8916 20812 8968
rect 20864 8916 20870 8968
rect 21376 8956 21404 8996
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24854 9024 24860 9036
rect 23891 8996 24860 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 20916 8928 21404 8956
rect 21453 8959 21511 8965
rect 20916 8888 20944 8928
rect 21453 8925 21465 8959
rect 21499 8956 21511 8959
rect 21542 8956 21548 8968
rect 21499 8928 21548 8956
rect 21499 8925 21511 8928
rect 21453 8919 21511 8925
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 23808 8928 24593 8956
rect 23808 8916 23814 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 20272 8860 20944 8888
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 26326 8888 26332 8900
rect 21048 8860 26332 8888
rect 21048 8848 21054 8860
rect 26326 8848 26332 8860
rect 26384 8848 26390 8900
rect 17405 8823 17463 8829
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 18414 8820 18420 8832
rect 17451 8792 18420 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18693 8823 18751 8829
rect 18693 8789 18705 8823
rect 18739 8820 18751 8823
rect 18782 8820 18788 8832
rect 18739 8792 18788 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 20162 8780 20168 8832
rect 20220 8820 20226 8832
rect 22554 8820 22560 8832
rect 20220 8792 22560 8820
rect 20220 8780 20226 8792
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19153 8619 19211 8625
rect 19153 8585 19165 8619
rect 19199 8585 19211 8619
rect 19153 8579 19211 8585
rect 16574 8508 16580 8560
rect 16632 8548 16638 8560
rect 19168 8548 19196 8579
rect 19794 8576 19800 8628
rect 19852 8576 19858 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20864 8588 20913 8616
rect 20864 8576 20870 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21266 8576 21272 8628
rect 21324 8576 21330 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 22094 8616 22100 8628
rect 21416 8588 22100 8616
rect 21416 8576 21422 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 26694 8616 26700 8628
rect 22296 8588 26700 8616
rect 16632 8520 19104 8548
rect 19168 8520 22232 8548
rect 16632 8508 16638 8520
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 19076 8480 19104 8520
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 17451 8452 19012 8480
rect 19076 8452 19349 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17862 8372 17868 8424
rect 17920 8372 17926 8424
rect 18141 8415 18199 8421
rect 18141 8381 18153 8415
rect 18187 8412 18199 8415
rect 18874 8412 18880 8424
rect 18187 8384 18880 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 18984 8412 19012 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8480 20039 8483
rect 20254 8480 20260 8492
rect 20027 8452 20260 8480
rect 20027 8449 20039 8452
rect 19981 8443 20039 8449
rect 20254 8440 20260 8452
rect 20312 8480 20318 8492
rect 20438 8480 20444 8492
rect 20312 8452 20444 8480
rect 20312 8440 20318 8452
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 19058 8412 19064 8424
rect 18984 8384 19064 8412
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 20640 8412 20668 8443
rect 22204 8412 22232 8520
rect 22296 8489 22324 8588
rect 26694 8576 26700 8588
rect 26752 8576 26758 8628
rect 22388 8520 24072 8548
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22388 8412 22416 8520
rect 24044 8489 24072 8520
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24946 8480 24952 8492
rect 24029 8443 24087 8449
rect 24688 8452 24952 8480
rect 19628 8384 20576 8412
rect 20640 8384 22094 8412
rect 22204 8384 22416 8412
rect 23293 8415 23351 8421
rect 17221 8347 17279 8353
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 19628 8344 19656 8384
rect 17267 8316 19656 8344
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 20438 8304 20444 8356
rect 20496 8304 20502 8356
rect 20548 8344 20576 8384
rect 21358 8344 21364 8356
rect 20548 8316 21364 8344
rect 21358 8304 21364 8316
rect 21416 8304 21422 8356
rect 22066 8344 22094 8384
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 24688 8412 24716 8452
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 23339 8384 24716 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 24210 8344 24216 8356
rect 22066 8316 24216 8344
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20220 8044 20545 8072
rect 20220 8032 20226 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 20809 8075 20867 8081
rect 20809 8041 20821 8075
rect 20855 8072 20867 8075
rect 20898 8072 20904 8084
rect 20855 8044 20904 8072
rect 20855 8041 20867 8044
rect 20809 8035 20867 8041
rect 20898 8032 20904 8044
rect 20956 8072 20962 8084
rect 20956 8044 24256 8072
rect 20956 8032 20962 8044
rect 22186 8004 22192 8016
rect 17696 7976 22192 8004
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7936 17463 7939
rect 17494 7936 17500 7948
rect 17451 7908 17500 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 17696 7945 17724 7976
rect 22186 7964 22192 7976
rect 22244 7964 22250 8016
rect 24228 8004 24256 8044
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 26418 8004 26424 8016
rect 24228 7976 26424 8004
rect 26418 7964 26424 7976
rect 26476 7964 26482 8016
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 23474 7936 23480 7948
rect 18739 7908 23480 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24854 7936 24860 7948
rect 23891 7908 24860 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19628 7732 19656 7831
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 20680 7840 21281 7868
rect 20680 7828 20686 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 22094 7828 22100 7880
rect 22152 7828 22158 7880
rect 22370 7828 22376 7880
rect 22428 7868 22434 7880
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 22428 7840 22661 7868
rect 22428 7828 22434 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24544 7840 24593 7868
rect 24544 7828 24550 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 20073 7803 20131 7809
rect 20073 7769 20085 7803
rect 20119 7800 20131 7803
rect 23382 7800 23388 7812
rect 20119 7772 23388 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 23382 7760 23388 7772
rect 23440 7760 23446 7812
rect 20806 7732 20812 7744
rect 19628 7704 20812 7732
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 20993 7735 21051 7741
rect 20993 7701 21005 7735
rect 21039 7732 21051 7735
rect 21082 7732 21088 7744
rect 21039 7704 21088 7732
rect 21039 7701 21051 7704
rect 20993 7695 21051 7701
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 21913 7735 21971 7741
rect 21913 7701 21925 7735
rect 21959 7732 21971 7735
rect 22186 7732 22192 7744
rect 21959 7704 22192 7732
rect 21959 7701 21971 7704
rect 21913 7695 21971 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17862 7528 17868 7540
rect 17451 7500 17868 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 17957 7531 18015 7537
rect 17957 7497 17969 7531
rect 18003 7528 18015 7531
rect 18322 7528 18328 7540
rect 18003 7500 18328 7528
rect 18003 7497 18015 7500
rect 17957 7491 18015 7497
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17972 7392 18000 7491
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 22646 7528 22652 7540
rect 18555 7500 22652 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 23750 7528 23756 7540
rect 23032 7500 23756 7528
rect 18414 7420 18420 7472
rect 18472 7460 18478 7472
rect 23032 7460 23060 7500
rect 23750 7488 23756 7500
rect 23808 7488 23814 7540
rect 18472 7432 19196 7460
rect 18472 7420 18478 7432
rect 17635 7364 18000 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 18690 7352 18696 7404
rect 18748 7352 18754 7404
rect 19168 7401 19196 7432
rect 19444 7432 23060 7460
rect 23293 7463 23351 7469
rect 19444 7401 19472 7432
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 19760 7364 20392 7392
rect 19760 7352 19766 7364
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 20257 7327 20315 7333
rect 20257 7324 20269 7327
rect 19392 7296 20269 7324
rect 19392 7284 19398 7296
rect 20257 7293 20269 7296
rect 20303 7293 20315 7327
rect 20364 7324 20392 7364
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20772 7364 20821 7392
rect 20772 7352 20778 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 21468 7324 21496 7355
rect 20364 7296 21496 7324
rect 20257 7287 20315 7293
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 22112 7256 22140 7355
rect 23474 7352 23480 7404
rect 23532 7392 23538 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23532 7364 23949 7392
rect 23532 7352 23538 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 16264 7228 22140 7256
rect 16264 7216 16270 7228
rect 20622 7148 20628 7200
rect 20680 7148 20686 7200
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 25038 7188 25044 7200
rect 21315 7160 25044 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 20717 6919 20775 6925
rect 20717 6885 20729 6919
rect 20763 6885 20775 6919
rect 20717 6879 20775 6885
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 17218 6848 17224 6860
rect 6328 6820 17224 6848
rect 6328 6808 6334 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 20732 6848 20760 6879
rect 22462 6848 22468 6860
rect 20732 6820 22468 6848
rect 22462 6808 22468 6820
rect 22520 6808 22526 6860
rect 24486 6808 24492 6860
rect 24544 6808 24550 6860
rect 24670 6808 24676 6860
rect 24728 6808 24734 6860
rect 19242 6740 19248 6792
rect 19300 6780 19306 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19300 6752 19625 6780
rect 19300 6740 19306 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 20622 6780 20628 6792
rect 20303 6752 20628 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 20901 6783 20959 6789
rect 20901 6749 20913 6783
rect 20947 6780 20959 6783
rect 21266 6780 21272 6792
rect 20947 6752 21272 6780
rect 20947 6749 20959 6752
rect 20901 6743 20959 6749
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 21376 6752 22661 6780
rect 21376 6712 21404 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24946 6780 24952 6792
rect 23891 6752 24952 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 25133 6783 25191 6789
rect 25133 6749 25145 6783
rect 25179 6780 25191 6783
rect 25222 6780 25228 6792
rect 25179 6752 25228 6780
rect 25179 6749 25191 6752
rect 25133 6743 25191 6749
rect 20088 6684 21404 6712
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 20088 6653 20116 6684
rect 21450 6672 21456 6724
rect 21508 6672 21514 6724
rect 21637 6715 21695 6721
rect 21637 6681 21649 6715
rect 21683 6712 21695 6715
rect 21726 6712 21732 6724
rect 21683 6684 21732 6712
rect 21683 6681 21695 6684
rect 21637 6675 21695 6681
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 22005 6715 22063 6721
rect 22005 6712 22017 6715
rect 21876 6684 22017 6712
rect 21876 6672 21882 6684
rect 22005 6681 22017 6684
rect 22051 6681 22063 6715
rect 22005 6675 22063 6681
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25148 6712 25176 6743
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 24903 6684 25176 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25314 6672 25320 6724
rect 25372 6672 25378 6724
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 16172 6616 19441 6644
rect 16172 6604 16178 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 21174 6604 21180 6656
rect 21232 6604 21238 6656
rect 22094 6604 22100 6656
rect 22152 6604 22158 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 19300 6412 19717 6440
rect 19300 6400 19306 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 20254 6440 20260 6452
rect 20211 6412 20260 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 20898 6400 20904 6452
rect 20956 6400 20962 6452
rect 21266 6400 21272 6452
rect 21324 6400 21330 6452
rect 25498 6440 25504 6452
rect 22066 6412 25504 6440
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 21818 6372 21824 6384
rect 16908 6344 21824 6372
rect 16908 6332 16914 6344
rect 21818 6332 21824 6344
rect 21876 6332 21882 6384
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20496 6276 20637 6304
rect 20496 6264 20502 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6304 21511 6307
rect 22066 6304 22094 6412
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 21499 6276 22094 6304
rect 21499 6273 21511 6276
rect 21453 6267 21511 6273
rect 22186 6264 22192 6316
rect 22244 6264 22250 6316
rect 23842 6264 23848 6316
rect 23900 6304 23906 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 23900 6276 23949 6304
rect 23900 6264 23906 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17276 6208 24348 6236
rect 17276 6196 17282 6208
rect 20441 6171 20499 6177
rect 20441 6137 20453 6171
rect 20487 6168 20499 6171
rect 23474 6168 23480 6180
rect 20487 6140 23480 6168
rect 20487 6137 20499 6140
rect 20441 6131 20499 6137
rect 23474 6128 23480 6140
rect 23532 6128 23538 6180
rect 24320 6168 24348 6208
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 25222 6168 25228 6180
rect 24320 6140 25228 6168
rect 25222 6128 25228 6140
rect 25280 6128 25286 6180
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 25501 5899 25559 5905
rect 25501 5865 25513 5899
rect 25547 5896 25559 5899
rect 25682 5896 25688 5908
rect 25547 5868 25688 5896
rect 25547 5865 25559 5868
rect 25501 5859 25559 5865
rect 25682 5856 25688 5868
rect 25740 5856 25746 5908
rect 21085 5831 21143 5837
rect 21085 5797 21097 5831
rect 21131 5828 21143 5831
rect 23382 5828 23388 5840
rect 21131 5800 23388 5828
rect 21131 5797 21143 5800
rect 21085 5791 21143 5797
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 25317 5831 25375 5837
rect 25317 5797 25329 5831
rect 25363 5828 25375 5831
rect 25406 5828 25412 5840
rect 25363 5800 25412 5828
rect 25363 5797 25375 5800
rect 25317 5791 25375 5797
rect 25406 5788 25412 5800
rect 25464 5828 25470 5840
rect 26786 5828 26792 5840
rect 25464 5800 26792 5828
rect 25464 5788 25470 5800
rect 26786 5788 26792 5800
rect 26844 5788 26850 5840
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 22005 5763 22063 5769
rect 18564 5732 21312 5760
rect 18564 5720 18570 5732
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 21284 5701 21312 5732
rect 22005 5729 22017 5763
rect 22051 5760 22063 5763
rect 25866 5760 25872 5772
rect 22051 5732 25872 5760
rect 22051 5729 22063 5732
rect 22005 5723 22063 5729
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 19576 5664 20637 5692
rect 19576 5652 19582 5664
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 21269 5695 21327 5701
rect 21269 5661 21281 5695
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 25038 5692 25044 5704
rect 24903 5664 25044 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 22738 5624 22744 5636
rect 20456 5596 22744 5624
rect 20456 5565 20484 5596
rect 22738 5584 22744 5596
rect 22796 5584 22802 5636
rect 20441 5559 20499 5565
rect 20441 5525 20453 5559
rect 20487 5525 20499 5559
rect 22848 5556 22876 5655
rect 25038 5652 25044 5664
rect 25096 5652 25102 5704
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 22848 5528 24685 5556
rect 20441 5519 20499 5525
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 24578 5352 24584 5364
rect 22066 5324 24584 5352
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5216 21511 5219
rect 22066 5216 22094 5324
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 23293 5287 23351 5293
rect 23293 5253 23305 5287
rect 23339 5284 23351 5287
rect 24854 5284 24860 5296
rect 23339 5256 24860 5284
rect 23339 5253 23351 5256
rect 23293 5247 23351 5253
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 21499 5188 22094 5216
rect 21499 5185 21511 5188
rect 21453 5179 21511 5185
rect 22278 5176 22284 5228
rect 22336 5176 22342 5228
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23808 5188 23949 5216
rect 23808 5176 23814 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 24578 5012 24584 5024
rect 21315 4984 24584 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 24578 4972 24584 4984
rect 24636 4972 24642 5024
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 22005 4811 22063 4817
rect 22005 4808 22017 4811
rect 15988 4780 22017 4808
rect 15988 4768 15994 4780
rect 22005 4777 22017 4780
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 25501 4811 25559 4817
rect 25501 4777 25513 4811
rect 25547 4808 25559 4811
rect 25682 4808 25688 4820
rect 25547 4780 25688 4808
rect 25547 4777 25559 4780
rect 25501 4771 25559 4777
rect 25682 4768 25688 4780
rect 25740 4768 25746 4820
rect 25225 4743 25283 4749
rect 25225 4709 25237 4743
rect 25271 4740 25283 4743
rect 25958 4740 25964 4752
rect 25271 4712 25964 4740
rect 25271 4709 25283 4712
rect 25225 4703 25283 4709
rect 25958 4700 25964 4712
rect 26016 4700 26022 4752
rect 25130 4672 25136 4684
rect 22848 4644 25136 4672
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22186 4604 22192 4616
rect 21775 4576 22192 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 22848 4613 22876 4644
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 22833 4607 22891 4613
rect 22833 4573 22845 4607
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 23440 4576 24869 4604
rect 23440 4564 23446 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 25498 4536 25504 4548
rect 23891 4508 25504 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 24670 4428 24676 4480
rect 24728 4428 24734 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 20303 4100 21128 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20162 4060 20168 4072
rect 19024 4032 20168 4060
rect 19024 4020 19030 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21100 3992 21128 4100
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 23658 4088 23664 4140
rect 23716 4128 23722 4140
rect 23937 4131 23995 4137
rect 23937 4128 23949 4131
rect 23716 4100 23949 4128
rect 23716 4088 23722 4100
rect 23937 4097 23949 4100
rect 23983 4097 23995 4131
rect 23937 4091 23995 4097
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 22186 4060 22192 4072
rect 21315 4032 22192 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22186 4020 22192 4032
rect 22244 4020 22250 4072
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 21100 3964 22094 3992
rect 23308 3964 24952 3992
rect 22066 3924 22094 3964
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 25590 3924 25596 3936
rect 22066 3896 25596 3924
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 25222 3680 25228 3732
rect 25280 3680 25286 3732
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 22796 3556 24900 3584
rect 22796 3544 22802 3556
rect 20993 3519 21051 3525
rect 20993 3485 21005 3519
rect 21039 3516 21051 3519
rect 21910 3516 21916 3528
rect 21039 3488 21916 3516
rect 21039 3485 21051 3488
rect 20993 3479 21051 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 24670 3516 24676 3528
rect 22879 3488 24676 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24872 3525 24900 3556
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24946 3448 24952 3460
rect 23891 3420 24952 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24946 3408 24952 3420
rect 25004 3408 25010 3460
rect 22278 3340 22284 3392
rect 22336 3380 22342 3392
rect 24673 3383 24731 3389
rect 24673 3380 24685 3383
rect 22336 3352 24685 3380
rect 22336 3340 22342 3352
rect 24673 3349 24685 3352
rect 24719 3349 24731 3383
rect 24673 3343 24731 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 25314 3176 25320 3188
rect 22066 3148 25320 3176
rect 22066 3108 22094 3148
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 18432 3080 22094 3108
rect 23293 3111 23351 3117
rect 18432 3049 18460 3080
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25130 3068 25136 3120
rect 25188 3068 25194 3120
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 20070 3000 20076 3052
rect 20128 3000 20134 3052
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 23934 3000 23940 3052
rect 23992 3000 23998 3052
rect 19426 2932 19432 2984
rect 19484 2932 19490 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6822 2592 6828 2644
rect 6880 2592 6886 2644
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 22094 2632 22100 2644
rect 19484 2604 22100 2632
rect 19484 2592 19490 2604
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 23290 2564 23296 2576
rect 20272 2536 23296 2564
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 20272 2437 20300 2536
rect 23290 2524 23296 2536
rect 23348 2524 23354 2576
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 23382 2496 23388 2508
rect 21315 2468 23388 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7055 2400 7297 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 22848 2292 22876 2391
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24636 2400 24777 2428
rect 24636 2388 24642 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 22848 2264 24593 2292
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 5632 26324 5684 26376
rect 22376 26324 22428 26376
rect 3608 26256 3660 26308
rect 19616 26256 19668 26308
rect 3700 26188 3752 26240
rect 17960 26188 18012 26240
rect 6276 26120 6328 26172
rect 19800 26120 19852 26172
rect 3148 25644 3200 25696
rect 10692 25644 10744 25696
rect 7380 25508 7432 25560
rect 23756 25508 23808 25560
rect 4068 25440 4120 25492
rect 20812 25440 20864 25492
rect 6552 25372 6604 25424
rect 22560 25372 22612 25424
rect 3792 25304 3844 25356
rect 23848 25304 23900 25356
rect 5264 25236 5316 25288
rect 18604 25236 18656 25288
rect 6184 25168 6236 25220
rect 24400 25168 24452 25220
rect 7288 25100 7340 25152
rect 24216 25100 24268 25152
rect 14372 25032 14424 25084
rect 20720 25032 20772 25084
rect 13544 24964 13596 25016
rect 23480 24964 23532 25016
rect 7196 24896 7248 24948
rect 22284 24896 22336 24948
rect 9496 24828 9548 24880
rect 22468 24828 22520 24880
rect 7748 24760 7800 24812
rect 19984 24760 20036 24812
rect 3976 24624 4028 24676
rect 11244 24624 11296 24676
rect 12164 24624 12216 24676
rect 16396 24624 16448 24676
rect 4160 24556 4212 24608
rect 14740 24556 14792 24608
rect 22376 24556 22428 24608
rect 24768 24556 24820 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 3332 24352 3384 24404
rect 4068 24352 4120 24404
rect 6460 24216 6512 24268
rect 12624 24352 12676 24404
rect 14464 24352 14516 24404
rect 15292 24352 15344 24404
rect 19616 24352 19668 24404
rect 20720 24352 20772 24404
rect 2688 24080 2740 24132
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 4068 24012 4120 24064
rect 4160 24012 4212 24064
rect 4896 24148 4948 24200
rect 11520 24284 11572 24336
rect 12348 24284 12400 24336
rect 12532 24284 12584 24336
rect 9680 24216 9732 24268
rect 13728 24216 13780 24268
rect 18328 24216 18380 24268
rect 7104 24148 7156 24200
rect 8668 24080 8720 24132
rect 9864 24191 9916 24200
rect 9864 24157 9873 24191
rect 9873 24157 9907 24191
rect 9907 24157 9916 24191
rect 9864 24148 9916 24157
rect 10968 24191 11020 24200
rect 10968 24157 10977 24191
rect 10977 24157 11011 24191
rect 11011 24157 11020 24191
rect 10968 24148 11020 24157
rect 9680 24080 9732 24132
rect 15200 24148 15252 24200
rect 16764 24148 16816 24200
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 22100 24284 22152 24336
rect 18696 24259 18748 24268
rect 18696 24225 18705 24259
rect 18705 24225 18739 24259
rect 18739 24225 18748 24259
rect 18696 24216 18748 24225
rect 18788 24216 18840 24268
rect 22836 24216 22888 24268
rect 23664 24216 23716 24268
rect 8392 24012 8444 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 10968 24012 11020 24064
rect 11060 24012 11112 24064
rect 14004 24012 14056 24064
rect 14924 24055 14976 24064
rect 14924 24021 14933 24055
rect 14933 24021 14967 24055
rect 14967 24021 14976 24055
rect 14924 24012 14976 24021
rect 15108 24012 15160 24064
rect 16304 24055 16356 24064
rect 16304 24021 16313 24055
rect 16313 24021 16347 24055
rect 16347 24021 16356 24055
rect 16304 24012 16356 24021
rect 16488 24012 16540 24064
rect 19524 24148 19576 24200
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22192 24148 22244 24157
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 20904 24080 20956 24132
rect 22376 24080 22428 24132
rect 17684 24012 17736 24064
rect 18788 24012 18840 24064
rect 19156 24012 19208 24064
rect 22100 24055 22152 24064
rect 22100 24021 22109 24055
rect 22109 24021 22143 24055
rect 22143 24021 22152 24055
rect 22100 24012 22152 24021
rect 24124 24012 24176 24064
rect 24860 24012 24912 24064
rect 24952 24012 25004 24064
rect 25504 24012 25556 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 5356 23740 5408 23792
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 4896 23672 4948 23724
rect 10140 23740 10192 23792
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 11336 23808 11388 23860
rect 13636 23740 13688 23792
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 1952 23604 2004 23656
rect 7564 23604 7616 23656
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 9772 23715 9824 23724
rect 9772 23681 9781 23715
rect 9781 23681 9815 23715
rect 9815 23681 9824 23715
rect 9772 23672 9824 23681
rect 10048 23672 10100 23724
rect 13820 23672 13872 23724
rect 15016 23740 15068 23792
rect 17592 23808 17644 23860
rect 20812 23808 20864 23860
rect 22284 23808 22336 23860
rect 18420 23740 18472 23792
rect 20904 23740 20956 23792
rect 22008 23740 22060 23792
rect 22836 23808 22888 23860
rect 24768 23740 24820 23792
rect 15292 23672 15344 23724
rect 16028 23672 16080 23724
rect 11336 23604 11388 23656
rect 11980 23604 12032 23656
rect 15200 23604 15252 23656
rect 15384 23604 15436 23656
rect 15476 23604 15528 23656
rect 16488 23672 16540 23724
rect 17408 23672 17460 23724
rect 23664 23672 23716 23724
rect 17960 23604 18012 23656
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 5172 23468 5224 23520
rect 7932 23468 7984 23520
rect 10416 23468 10468 23520
rect 10968 23468 11020 23520
rect 12256 23468 12308 23520
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 14648 23468 14700 23520
rect 15752 23468 15804 23520
rect 17040 23468 17092 23520
rect 17224 23468 17276 23520
rect 19432 23468 19484 23520
rect 24952 23536 25004 23588
rect 20720 23468 20772 23520
rect 24032 23511 24084 23520
rect 24032 23477 24041 23511
rect 24041 23477 24075 23511
rect 24075 23477 24084 23511
rect 24032 23468 24084 23477
rect 25136 23468 25188 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 3884 23264 3936 23316
rect 4896 23264 4948 23316
rect 8392 23264 8444 23316
rect 11612 23264 11664 23316
rect 4620 23128 4672 23180
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 11152 23196 11204 23248
rect 12440 23264 12492 23316
rect 12624 23196 12676 23248
rect 13636 23196 13688 23248
rect 7656 23128 7708 23180
rect 9404 23128 9456 23180
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 5448 23103 5500 23112
rect 5448 23069 5457 23103
rect 5457 23069 5491 23103
rect 5491 23069 5500 23103
rect 5448 23060 5500 23069
rect 1584 23035 1636 23044
rect 1584 23001 1593 23035
rect 1593 23001 1627 23035
rect 1627 23001 1636 23035
rect 1584 22992 1636 23001
rect 4988 22992 5040 23044
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 10140 23060 10192 23112
rect 12256 23060 12308 23112
rect 13912 23128 13964 23180
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 17040 23264 17092 23316
rect 17684 23264 17736 23316
rect 17776 23264 17828 23316
rect 18328 23307 18380 23316
rect 18328 23273 18337 23307
rect 18337 23273 18371 23307
rect 18371 23273 18380 23307
rect 18328 23264 18380 23273
rect 18604 23307 18656 23316
rect 18604 23273 18613 23307
rect 18613 23273 18647 23307
rect 18647 23273 18656 23307
rect 18604 23264 18656 23273
rect 16488 23196 16540 23248
rect 17500 23196 17552 23248
rect 21548 23264 21600 23316
rect 22008 23264 22060 23316
rect 23664 23264 23716 23316
rect 17776 23171 17828 23180
rect 17776 23137 17785 23171
rect 17785 23137 17819 23171
rect 17819 23137 17828 23171
rect 17776 23128 17828 23137
rect 17868 23128 17920 23180
rect 19800 23128 19852 23180
rect 20904 23128 20956 23180
rect 22284 23128 22336 23180
rect 23296 23128 23348 23180
rect 23664 23128 23716 23180
rect 24032 23128 24084 23180
rect 13820 23060 13872 23112
rect 14280 23060 14332 23112
rect 17132 23060 17184 23112
rect 17500 23060 17552 23112
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 17960 23060 18012 23112
rect 19340 23060 19392 23112
rect 9864 22992 9916 23044
rect 1768 22967 1820 22976
rect 1768 22933 1777 22967
rect 1777 22933 1811 22967
rect 1811 22933 1820 22967
rect 1768 22924 1820 22933
rect 2688 22924 2740 22976
rect 7840 22924 7892 22976
rect 8944 22924 8996 22976
rect 11980 22992 12032 23044
rect 12624 23035 12676 23044
rect 12624 23001 12633 23035
rect 12633 23001 12667 23035
rect 12667 23001 12676 23035
rect 12624 22992 12676 23001
rect 14832 22992 14884 23044
rect 15752 22992 15804 23044
rect 17316 22992 17368 23044
rect 18328 22992 18380 23044
rect 10324 22924 10376 22976
rect 12348 22924 12400 22976
rect 16672 22924 16724 22976
rect 16764 22967 16816 22976
rect 16764 22933 16773 22967
rect 16773 22933 16807 22967
rect 16807 22933 16816 22967
rect 16764 22924 16816 22933
rect 17040 22924 17092 22976
rect 17592 22924 17644 22976
rect 18696 22992 18748 23044
rect 19800 22992 19852 23044
rect 18972 22967 19024 22976
rect 18972 22933 18981 22967
rect 18981 22933 19015 22967
rect 19015 22933 19024 22967
rect 18972 22924 19024 22933
rect 19432 22924 19484 22976
rect 24768 22992 24820 23044
rect 26792 22992 26844 23044
rect 22744 22924 22796 22976
rect 23572 22924 23624 22976
rect 23940 22924 23992 22976
rect 25044 22967 25096 22976
rect 25044 22933 25053 22967
rect 25053 22933 25087 22967
rect 25087 22933 25096 22967
rect 25044 22924 25096 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 2228 22720 2280 22772
rect 1768 22652 1820 22704
rect 3700 22652 3752 22704
rect 4252 22652 4304 22704
rect 5356 22652 5408 22704
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 5908 22652 5960 22704
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 6644 22627 6696 22636
rect 6644 22593 6653 22627
rect 6653 22593 6687 22627
rect 6687 22593 6696 22627
rect 6644 22584 6696 22593
rect 6920 22584 6972 22636
rect 7288 22627 7340 22636
rect 7288 22593 7297 22627
rect 7297 22593 7331 22627
rect 7331 22593 7340 22627
rect 7288 22584 7340 22593
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 11152 22652 11204 22704
rect 10784 22584 10836 22636
rect 6736 22516 6788 22568
rect 9036 22516 9088 22568
rect 1308 22380 1360 22432
rect 6736 22423 6788 22432
rect 6736 22389 6745 22423
rect 6745 22389 6779 22423
rect 6779 22389 6788 22423
rect 6736 22380 6788 22389
rect 7748 22448 7800 22500
rect 9772 22516 9824 22568
rect 11888 22584 11940 22636
rect 11152 22559 11204 22568
rect 11152 22525 11161 22559
rect 11161 22525 11195 22559
rect 11195 22525 11204 22559
rect 11152 22516 11204 22525
rect 12348 22584 12400 22636
rect 12440 22584 12492 22636
rect 13820 22652 13872 22704
rect 14556 22652 14608 22704
rect 15384 22763 15436 22772
rect 15384 22729 15393 22763
rect 15393 22729 15427 22763
rect 15427 22729 15436 22763
rect 15384 22720 15436 22729
rect 15936 22695 15988 22704
rect 15936 22661 15945 22695
rect 15945 22661 15979 22695
rect 15979 22661 15988 22695
rect 15936 22652 15988 22661
rect 16304 22652 16356 22704
rect 16120 22584 16172 22636
rect 17868 22720 17920 22772
rect 17960 22720 18012 22772
rect 18972 22720 19024 22772
rect 19524 22720 19576 22772
rect 20904 22720 20956 22772
rect 21548 22720 21600 22772
rect 24308 22720 24360 22772
rect 17132 22695 17184 22704
rect 17132 22661 17141 22695
rect 17141 22661 17175 22695
rect 17175 22661 17184 22695
rect 17132 22652 17184 22661
rect 17684 22652 17736 22704
rect 19892 22652 19944 22704
rect 22284 22652 22336 22704
rect 23480 22652 23532 22704
rect 19708 22584 19760 22636
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 16764 22516 16816 22568
rect 15108 22448 15160 22500
rect 15200 22448 15252 22500
rect 11704 22423 11756 22432
rect 11704 22389 11713 22423
rect 11713 22389 11747 22423
rect 11747 22389 11756 22423
rect 11704 22380 11756 22389
rect 11980 22380 12032 22432
rect 16396 22423 16448 22432
rect 16396 22389 16405 22423
rect 16405 22389 16439 22423
rect 16439 22389 16448 22423
rect 16396 22380 16448 22389
rect 18420 22448 18472 22500
rect 19248 22448 19300 22500
rect 20720 22559 20772 22568
rect 20720 22525 20729 22559
rect 20729 22525 20763 22559
rect 20763 22525 20772 22559
rect 20720 22516 20772 22525
rect 20352 22448 20404 22500
rect 22468 22559 22520 22568
rect 22468 22525 22477 22559
rect 22477 22525 22511 22559
rect 22511 22525 22520 22559
rect 22468 22516 22520 22525
rect 22284 22448 22336 22500
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 24768 22516 24820 22568
rect 25412 22448 25464 22500
rect 17592 22380 17644 22432
rect 17776 22380 17828 22432
rect 18972 22380 19024 22432
rect 20720 22380 20772 22432
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 22836 22380 22888 22432
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 2228 22176 2280 22228
rect 2504 22176 2556 22228
rect 3976 22176 4028 22228
rect 9588 22176 9640 22228
rect 9680 22176 9732 22228
rect 11704 22176 11756 22228
rect 12716 22176 12768 22228
rect 14188 22176 14240 22228
rect 14924 22176 14976 22228
rect 15016 22176 15068 22228
rect 1860 22108 1912 22160
rect 10140 22108 10192 22160
rect 1492 22040 1544 22092
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 2504 21972 2556 22024
rect 2596 21972 2648 22024
rect 3976 21904 4028 21956
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 10600 22040 10652 22092
rect 10968 22083 11020 22092
rect 10968 22049 10977 22083
rect 10977 22049 11011 22083
rect 11011 22049 11020 22083
rect 10968 22040 11020 22049
rect 11336 22040 11388 22092
rect 14280 22083 14332 22092
rect 14280 22049 14289 22083
rect 14289 22049 14323 22083
rect 14323 22049 14332 22083
rect 14280 22040 14332 22049
rect 16028 22151 16080 22160
rect 16028 22117 16037 22151
rect 16037 22117 16071 22151
rect 16071 22117 16080 22151
rect 16028 22108 16080 22117
rect 15752 22040 15804 22092
rect 17684 22176 17736 22228
rect 19064 22176 19116 22228
rect 19984 22176 20036 22228
rect 21916 22176 21968 22228
rect 26884 22176 26936 22228
rect 9036 21972 9088 22024
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 16856 22040 16908 22092
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18236 22040 18288 22049
rect 18696 22040 18748 22092
rect 21272 22040 21324 22092
rect 23480 22108 23532 22160
rect 24124 22108 24176 22160
rect 23756 22040 23808 22092
rect 25228 22083 25280 22092
rect 25228 22049 25237 22083
rect 25237 22049 25271 22083
rect 25271 22049 25280 22083
rect 25228 22040 25280 22049
rect 8576 21904 8628 21956
rect 10876 21904 10928 21956
rect 12348 21904 12400 21956
rect 3700 21836 3752 21888
rect 4252 21836 4304 21888
rect 5448 21836 5500 21888
rect 6460 21836 6512 21888
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 9312 21836 9364 21888
rect 9404 21836 9456 21888
rect 11796 21836 11848 21888
rect 11980 21836 12032 21888
rect 12256 21836 12308 21888
rect 12532 21836 12584 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 14556 21904 14608 21956
rect 16028 21904 16080 21956
rect 16212 21904 16264 21956
rect 16488 21972 16540 22024
rect 16580 21972 16632 22024
rect 18972 21972 19024 22024
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 19616 21972 19668 22024
rect 21640 21972 21692 22024
rect 22008 21972 22060 22024
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 25596 21972 25648 22024
rect 17500 21904 17552 21956
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17960 21836 18012 21888
rect 19064 21836 19116 21888
rect 21088 21904 21140 21956
rect 25780 21904 25832 21956
rect 19616 21879 19668 21888
rect 19616 21845 19625 21879
rect 19625 21845 19659 21879
rect 19659 21845 19668 21879
rect 19616 21836 19668 21845
rect 20720 21836 20772 21888
rect 22008 21836 22060 21888
rect 22468 21836 22520 21888
rect 22652 21836 22704 21888
rect 23756 21836 23808 21888
rect 26608 21836 26660 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 1584 21632 1636 21684
rect 3976 21632 4028 21684
rect 1952 21564 2004 21616
rect 2872 21564 2924 21616
rect 1768 21496 1820 21548
rect 6736 21564 6788 21616
rect 7840 21564 7892 21616
rect 10784 21564 10836 21616
rect 11244 21632 11296 21684
rect 12256 21632 12308 21684
rect 12532 21632 12584 21684
rect 14096 21632 14148 21684
rect 14188 21675 14240 21684
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 17684 21632 17736 21684
rect 3700 21496 3752 21548
rect 4620 21496 4672 21548
rect 5264 21496 5316 21548
rect 7104 21496 7156 21548
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 14464 21564 14516 21616
rect 15752 21564 15804 21616
rect 11520 21496 11572 21548
rect 12532 21496 12584 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 2872 21360 2924 21412
rect 6460 21360 6512 21412
rect 7472 21428 7524 21480
rect 12164 21428 12216 21480
rect 12256 21428 12308 21480
rect 14556 21496 14608 21548
rect 14924 21496 14976 21548
rect 10600 21360 10652 21412
rect 12808 21471 12860 21480
rect 12808 21437 12817 21471
rect 12817 21437 12851 21471
rect 12851 21437 12860 21471
rect 12808 21428 12860 21437
rect 13084 21428 13136 21480
rect 15292 21428 15344 21480
rect 16304 21496 16356 21548
rect 18696 21632 18748 21684
rect 21088 21632 21140 21684
rect 21640 21632 21692 21684
rect 22192 21632 22244 21684
rect 22744 21632 22796 21684
rect 24952 21632 25004 21684
rect 25780 21632 25832 21684
rect 17040 21496 17092 21548
rect 19064 21496 19116 21548
rect 20812 21539 20864 21548
rect 20812 21505 20821 21539
rect 20821 21505 20855 21539
rect 20855 21505 20864 21539
rect 20812 21496 20864 21505
rect 20996 21496 21048 21548
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 15568 21471 15620 21480
rect 15568 21437 15577 21471
rect 15577 21437 15611 21471
rect 15611 21437 15620 21471
rect 15568 21428 15620 21437
rect 4712 21292 4764 21344
rect 6092 21292 6144 21344
rect 8484 21292 8536 21344
rect 9404 21292 9456 21344
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 14188 21360 14240 21412
rect 15384 21360 15436 21412
rect 15752 21360 15804 21412
rect 13636 21292 13688 21344
rect 14372 21292 14424 21344
rect 17316 21428 17368 21480
rect 17408 21428 17460 21480
rect 17500 21471 17552 21480
rect 17500 21437 17509 21471
rect 17509 21437 17543 21471
rect 17543 21437 17552 21471
rect 17500 21428 17552 21437
rect 16948 21360 17000 21412
rect 18420 21428 18472 21480
rect 19616 21428 19668 21480
rect 19708 21428 19760 21480
rect 18604 21360 18656 21412
rect 20720 21360 20772 21412
rect 20904 21471 20956 21480
rect 20904 21437 20913 21471
rect 20913 21437 20947 21471
rect 20947 21437 20956 21471
rect 20904 21428 20956 21437
rect 21364 21428 21416 21480
rect 23296 21496 23348 21548
rect 24768 21496 24820 21548
rect 22744 21360 22796 21412
rect 16580 21292 16632 21344
rect 16764 21292 16816 21344
rect 17868 21292 17920 21344
rect 19340 21292 19392 21344
rect 19984 21292 20036 21344
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 21916 21292 21968 21344
rect 24768 21292 24820 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 1768 21088 1820 21140
rect 4712 21088 4764 21140
rect 14188 21088 14240 21140
rect 17592 21088 17644 21140
rect 18328 21088 18380 21140
rect 20812 21088 20864 21140
rect 6920 21020 6972 21072
rect 9312 21020 9364 21072
rect 10232 21020 10284 21072
rect 15016 21020 15068 21072
rect 4896 20995 4948 21004
rect 4896 20961 4905 20995
rect 4905 20961 4939 20995
rect 4939 20961 4948 20995
rect 4896 20952 4948 20961
rect 6828 20952 6880 21004
rect 8576 20952 8628 21004
rect 8852 20952 8904 21004
rect 9036 20952 9088 21004
rect 11796 20952 11848 21004
rect 16764 21020 16816 21072
rect 17684 21020 17736 21072
rect 18420 21020 18472 21072
rect 2412 20884 2464 20936
rect 1952 20816 2004 20868
rect 1400 20748 1452 20800
rect 2688 20748 2740 20800
rect 4252 20884 4304 20936
rect 7288 20884 7340 20936
rect 7564 20884 7616 20936
rect 8392 20884 8444 20936
rect 9128 20927 9180 20936
rect 9128 20893 9137 20927
rect 9137 20893 9171 20927
rect 9171 20893 9180 20927
rect 9128 20884 9180 20893
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 11060 20884 11112 20936
rect 12900 20884 12952 20936
rect 14464 20884 14516 20936
rect 16120 20995 16172 21004
rect 16120 20961 16129 20995
rect 16129 20961 16163 20995
rect 16163 20961 16172 20995
rect 16120 20952 16172 20961
rect 16580 20952 16632 21004
rect 18328 20995 18380 21004
rect 18328 20961 18337 20995
rect 18337 20961 18371 20995
rect 18371 20961 18380 20995
rect 18328 20952 18380 20961
rect 18696 20952 18748 21004
rect 20720 21020 20772 21072
rect 19708 20952 19760 21004
rect 20352 20952 20404 21004
rect 22652 21088 22704 21140
rect 22928 21088 22980 21140
rect 22008 21020 22060 21072
rect 21916 20952 21968 21004
rect 22836 20952 22888 21004
rect 24860 20952 24912 21004
rect 25412 20952 25464 21004
rect 26792 20952 26844 21004
rect 8300 20816 8352 20868
rect 8576 20816 8628 20868
rect 11520 20816 11572 20868
rect 14096 20816 14148 20868
rect 15660 20884 15712 20936
rect 18604 20884 18656 20936
rect 19340 20884 19392 20936
rect 21088 20884 21140 20936
rect 22560 20884 22612 20936
rect 15476 20816 15528 20868
rect 16212 20816 16264 20868
rect 6460 20748 6512 20800
rect 6644 20748 6696 20800
rect 10600 20748 10652 20800
rect 14556 20748 14608 20800
rect 14924 20791 14976 20800
rect 14924 20757 14933 20791
rect 14933 20757 14967 20791
rect 14967 20757 14976 20791
rect 14924 20748 14976 20757
rect 15568 20748 15620 20800
rect 17040 20791 17092 20800
rect 17040 20757 17049 20791
rect 17049 20757 17083 20791
rect 17083 20757 17092 20791
rect 17040 20748 17092 20757
rect 19708 20859 19760 20868
rect 19708 20825 19717 20859
rect 19717 20825 19751 20859
rect 19751 20825 19760 20859
rect 19708 20816 19760 20825
rect 20168 20816 20220 20868
rect 21272 20748 21324 20800
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 22468 20816 22520 20868
rect 23572 20748 23624 20800
rect 23940 20791 23992 20800
rect 23940 20757 23949 20791
rect 23949 20757 23983 20791
rect 23983 20757 23992 20791
rect 23940 20748 23992 20757
rect 24032 20791 24084 20800
rect 24032 20757 24041 20791
rect 24041 20757 24075 20791
rect 24075 20757 24084 20791
rect 24032 20748 24084 20757
rect 24584 20791 24636 20800
rect 24584 20757 24593 20791
rect 24593 20757 24627 20791
rect 24627 20757 24636 20791
rect 24584 20748 24636 20757
rect 25412 20748 25464 20800
rect 25596 20748 25648 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 6920 20544 6972 20596
rect 7472 20587 7524 20596
rect 7472 20553 7481 20587
rect 7481 20553 7515 20587
rect 7515 20553 7524 20587
rect 7472 20544 7524 20553
rect 1860 20451 1912 20460
rect 1860 20417 1869 20451
rect 1869 20417 1903 20451
rect 1903 20417 1912 20451
rect 1860 20408 1912 20417
rect 7564 20476 7616 20528
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 2780 20340 2832 20392
rect 6000 20408 6052 20460
rect 6092 20408 6144 20460
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 6920 20408 6972 20460
rect 7748 20408 7800 20460
rect 12808 20544 12860 20596
rect 13360 20544 13412 20596
rect 14188 20544 14240 20596
rect 16488 20544 16540 20596
rect 8576 20519 8628 20528
rect 8576 20485 8585 20519
rect 8585 20485 8619 20519
rect 8619 20485 8628 20519
rect 8576 20476 8628 20485
rect 8116 20408 8168 20460
rect 9588 20476 9640 20528
rect 11520 20476 11572 20528
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 11060 20408 11112 20460
rect 11244 20408 11296 20460
rect 12624 20476 12676 20528
rect 13452 20408 13504 20460
rect 13820 20476 13872 20528
rect 16304 20519 16356 20528
rect 16304 20485 16313 20519
rect 16313 20485 16347 20519
rect 16347 20485 16356 20519
rect 16304 20476 16356 20485
rect 5448 20340 5500 20392
rect 9404 20340 9456 20392
rect 12256 20340 12308 20392
rect 8300 20272 8352 20324
rect 10416 20272 10468 20324
rect 11980 20272 12032 20324
rect 12624 20383 12676 20392
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 15108 20340 15160 20392
rect 3976 20204 4028 20256
rect 7932 20204 7984 20256
rect 11060 20204 11112 20256
rect 11428 20204 11480 20256
rect 11796 20204 11848 20256
rect 15016 20272 15068 20324
rect 16120 20451 16172 20460
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 17224 20519 17276 20528
rect 17224 20485 17233 20519
rect 17233 20485 17267 20519
rect 17267 20485 17276 20519
rect 17224 20476 17276 20485
rect 20168 20544 20220 20596
rect 21548 20544 21600 20596
rect 22008 20544 22060 20596
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 22100 20476 22152 20528
rect 24768 20476 24820 20528
rect 21456 20408 21508 20460
rect 22376 20408 22428 20460
rect 22836 20408 22888 20460
rect 23296 20408 23348 20460
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 20260 20340 20312 20392
rect 20812 20340 20864 20392
rect 16396 20272 16448 20324
rect 15476 20204 15528 20256
rect 19708 20204 19760 20256
rect 22284 20272 22336 20324
rect 22560 20272 22612 20324
rect 24216 20340 24268 20392
rect 21548 20247 21600 20256
rect 21548 20213 21557 20247
rect 21557 20213 21591 20247
rect 21591 20213 21600 20247
rect 21548 20204 21600 20213
rect 23848 20204 23900 20256
rect 25688 20204 25740 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 1492 20000 1544 20052
rect 4160 20000 4212 20052
rect 7656 20000 7708 20052
rect 8944 20043 8996 20052
rect 6000 19932 6052 19984
rect 8024 19932 8076 19984
rect 2320 19864 2372 19916
rect 6368 19864 6420 19916
rect 8944 20009 8953 20043
rect 8953 20009 8987 20043
rect 8987 20009 8996 20043
rect 8944 20000 8996 20009
rect 9772 20000 9824 20052
rect 10600 20000 10652 20052
rect 9312 19932 9364 19984
rect 10784 19932 10836 19984
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 4804 19796 4856 19848
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 9588 19864 9640 19916
rect 10416 19864 10468 19916
rect 15476 20000 15528 20052
rect 20168 20000 20220 20052
rect 20536 20000 20588 20052
rect 21456 20000 21508 20052
rect 21916 20000 21968 20052
rect 25044 20000 25096 20052
rect 25596 20000 25648 20052
rect 26056 20000 26108 20052
rect 3424 19728 3476 19780
rect 3792 19728 3844 19780
rect 1400 19660 1452 19712
rect 1952 19660 2004 19712
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 8024 19796 8076 19848
rect 5724 19728 5776 19780
rect 6000 19728 6052 19780
rect 6552 19771 6604 19780
rect 6552 19737 6561 19771
rect 6561 19737 6595 19771
rect 6595 19737 6604 19771
rect 6552 19728 6604 19737
rect 7012 19728 7064 19780
rect 7288 19728 7340 19780
rect 9772 19796 9824 19848
rect 10324 19796 10376 19848
rect 11060 19864 11112 19916
rect 13360 19907 13412 19916
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 15752 19932 15804 19984
rect 17592 19932 17644 19984
rect 18144 19932 18196 19984
rect 18420 19932 18472 19984
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 14004 19796 14056 19848
rect 14188 19796 14240 19848
rect 16028 19796 16080 19848
rect 16304 19796 16356 19848
rect 20812 19864 20864 19916
rect 23296 19864 23348 19916
rect 23664 19864 23716 19916
rect 24492 19864 24544 19916
rect 24860 19864 24912 19916
rect 18420 19796 18472 19848
rect 9588 19728 9640 19780
rect 13452 19728 13504 19780
rect 13544 19728 13596 19780
rect 19708 19728 19760 19780
rect 5540 19660 5592 19712
rect 5816 19660 5868 19712
rect 8392 19660 8444 19712
rect 8576 19703 8628 19712
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 9772 19660 9824 19712
rect 10600 19660 10652 19712
rect 10876 19660 10928 19712
rect 13176 19660 13228 19712
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 15108 19660 15160 19712
rect 15384 19703 15436 19712
rect 15384 19669 15393 19703
rect 15393 19669 15427 19703
rect 15427 19669 15436 19703
rect 15384 19660 15436 19669
rect 15476 19660 15528 19712
rect 16304 19660 16356 19712
rect 16764 19703 16816 19712
rect 16764 19669 16773 19703
rect 16773 19669 16807 19703
rect 16807 19669 16816 19703
rect 16764 19660 16816 19669
rect 17408 19660 17460 19712
rect 18144 19703 18196 19712
rect 18144 19669 18153 19703
rect 18153 19669 18187 19703
rect 18187 19669 18196 19703
rect 18144 19660 18196 19669
rect 18512 19660 18564 19712
rect 18880 19660 18932 19712
rect 19432 19703 19484 19712
rect 19432 19669 19441 19703
rect 19441 19669 19475 19703
rect 19475 19669 19484 19703
rect 19432 19660 19484 19669
rect 24952 19796 25004 19848
rect 21456 19728 21508 19780
rect 22744 19728 22796 19780
rect 20812 19660 20864 19712
rect 21272 19660 21324 19712
rect 21640 19660 21692 19712
rect 22376 19660 22428 19712
rect 23572 19660 23624 19712
rect 25412 19728 25464 19780
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 1492 19499 1544 19508
rect 1492 19465 1501 19499
rect 1501 19465 1535 19499
rect 1535 19465 1544 19499
rect 1492 19456 1544 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 4160 19456 4212 19508
rect 4344 19388 4396 19440
rect 4252 19320 4304 19372
rect 9680 19456 9732 19508
rect 11612 19456 11664 19508
rect 7472 19431 7524 19440
rect 7472 19397 7481 19431
rect 7481 19397 7515 19431
rect 7515 19397 7524 19431
rect 7472 19388 7524 19397
rect 8576 19388 8628 19440
rect 10876 19388 10928 19440
rect 4804 19320 4856 19372
rect 5816 19320 5868 19372
rect 7840 19320 7892 19372
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 13820 19456 13872 19508
rect 14556 19456 14608 19508
rect 14740 19456 14792 19508
rect 19432 19456 19484 19508
rect 21272 19456 21324 19508
rect 22100 19456 22152 19508
rect 22468 19499 22520 19508
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 23940 19456 23992 19508
rect 25228 19456 25280 19508
rect 26516 19456 26568 19508
rect 13452 19388 13504 19440
rect 14280 19388 14332 19440
rect 16396 19388 16448 19440
rect 20904 19388 20956 19440
rect 24952 19388 25004 19440
rect 14004 19320 14056 19372
rect 1676 19252 1728 19304
rect 3884 19252 3936 19304
rect 9404 19252 9456 19304
rect 10692 19252 10744 19304
rect 11612 19295 11664 19304
rect 11612 19261 11621 19295
rect 11621 19261 11655 19295
rect 11655 19261 11664 19295
rect 11612 19252 11664 19261
rect 11704 19252 11756 19304
rect 13728 19252 13780 19304
rect 8668 19184 8720 19236
rect 10968 19184 11020 19236
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 6828 19116 6880 19168
rect 7840 19116 7892 19168
rect 10048 19116 10100 19168
rect 10416 19116 10468 19168
rect 10876 19116 10928 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 14004 19184 14056 19236
rect 16488 19320 16540 19372
rect 13176 19116 13228 19168
rect 13360 19116 13412 19168
rect 16028 19252 16080 19304
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 17868 19252 17920 19304
rect 20168 19252 20220 19304
rect 20720 19252 20772 19304
rect 22652 19320 22704 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 25228 19320 25280 19372
rect 26056 19320 26108 19372
rect 26240 19320 26292 19372
rect 15016 19184 15068 19236
rect 15752 19184 15804 19236
rect 16396 19184 16448 19236
rect 17040 19184 17092 19236
rect 21180 19252 21232 19304
rect 22284 19252 22336 19304
rect 23664 19252 23716 19304
rect 14740 19116 14792 19168
rect 14924 19116 14976 19168
rect 15384 19116 15436 19168
rect 16212 19116 16264 19168
rect 16948 19116 17000 19168
rect 21548 19184 21600 19236
rect 21732 19184 21784 19236
rect 19340 19116 19392 19168
rect 19432 19116 19484 19168
rect 22100 19116 22152 19168
rect 22560 19116 22612 19168
rect 22744 19116 22796 19168
rect 25504 19252 25556 19304
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 2596 18955 2648 18964
rect 2596 18921 2605 18955
rect 2605 18921 2639 18955
rect 2639 18921 2648 18955
rect 2596 18912 2648 18921
rect 4620 18912 4672 18964
rect 5448 18955 5500 18964
rect 5448 18921 5457 18955
rect 5457 18921 5491 18955
rect 5491 18921 5500 18955
rect 5448 18912 5500 18921
rect 8760 18912 8812 18964
rect 9772 18912 9824 18964
rect 10232 18912 10284 18964
rect 11612 18912 11664 18964
rect 13636 18912 13688 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 14556 18912 14608 18964
rect 23388 18912 23440 18964
rect 25320 18912 25372 18964
rect 26056 18912 26108 18964
rect 2780 18844 2832 18896
rect 3792 18844 3844 18896
rect 3332 18776 3384 18828
rect 3976 18819 4028 18828
rect 3976 18785 3985 18819
rect 3985 18785 4019 18819
rect 4019 18785 4028 18819
rect 3976 18776 4028 18785
rect 5172 18776 5224 18828
rect 6552 18776 6604 18828
rect 8760 18776 8812 18828
rect 10048 18776 10100 18828
rect 11888 18776 11940 18828
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 6092 18708 6144 18760
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 7564 18640 7616 18692
rect 10324 18708 10376 18760
rect 11336 18708 11388 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 13820 18776 13872 18828
rect 14280 18776 14332 18828
rect 15384 18844 15436 18896
rect 15476 18844 15528 18896
rect 17224 18887 17276 18896
rect 17224 18853 17233 18887
rect 17233 18853 17267 18887
rect 17267 18853 17276 18887
rect 17224 18844 17276 18853
rect 16764 18776 16816 18828
rect 17592 18776 17644 18828
rect 11060 18640 11112 18692
rect 3056 18572 3108 18624
rect 3608 18572 3660 18624
rect 5172 18615 5224 18624
rect 5172 18581 5181 18615
rect 5181 18581 5215 18615
rect 5215 18581 5224 18615
rect 5172 18572 5224 18581
rect 6368 18615 6420 18624
rect 6368 18581 6377 18615
rect 6377 18581 6411 18615
rect 6411 18581 6420 18615
rect 6368 18572 6420 18581
rect 6828 18572 6880 18624
rect 7748 18572 7800 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 8668 18572 8720 18624
rect 9588 18615 9640 18624
rect 9588 18581 9597 18615
rect 9597 18581 9631 18615
rect 9631 18581 9640 18615
rect 9588 18572 9640 18581
rect 13268 18640 13320 18692
rect 13452 18683 13504 18692
rect 13452 18649 13461 18683
rect 13461 18649 13495 18683
rect 13495 18649 13504 18683
rect 13452 18640 13504 18649
rect 13636 18640 13688 18692
rect 13728 18640 13780 18692
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 12900 18572 12952 18624
rect 15016 18708 15068 18760
rect 17040 18708 17092 18760
rect 17868 18708 17920 18760
rect 19432 18844 19484 18896
rect 19616 18844 19668 18896
rect 19340 18776 19392 18828
rect 19248 18708 19300 18760
rect 21732 18708 21784 18760
rect 22744 18776 22796 18828
rect 25504 18844 25556 18896
rect 25688 18776 25740 18828
rect 16212 18640 16264 18692
rect 17776 18640 17828 18692
rect 15752 18572 15804 18624
rect 17040 18572 17092 18624
rect 18328 18572 18380 18624
rect 19156 18640 19208 18692
rect 19432 18640 19484 18692
rect 20628 18683 20680 18692
rect 20628 18649 20637 18683
rect 20637 18649 20671 18683
rect 20671 18649 20680 18683
rect 20628 18640 20680 18649
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 23020 18640 23072 18649
rect 24032 18640 24084 18692
rect 25136 18640 25188 18692
rect 20536 18572 20588 18624
rect 22376 18572 22428 18624
rect 22652 18572 22704 18624
rect 23388 18572 23440 18624
rect 23664 18572 23716 18624
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 25320 18572 25372 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 3056 18232 3108 18284
rect 8668 18368 8720 18420
rect 9312 18368 9364 18420
rect 4344 18232 4396 18284
rect 5632 18300 5684 18352
rect 6184 18343 6236 18352
rect 6184 18309 6193 18343
rect 6193 18309 6227 18343
rect 6227 18309 6236 18343
rect 6184 18300 6236 18309
rect 8300 18300 8352 18352
rect 8576 18300 8628 18352
rect 10876 18368 10928 18420
rect 11336 18368 11388 18420
rect 13544 18368 13596 18420
rect 13820 18368 13872 18420
rect 14004 18368 14056 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 14924 18368 14976 18420
rect 7380 18232 7432 18284
rect 1860 18207 1912 18216
rect 1860 18173 1869 18207
rect 1869 18173 1903 18207
rect 1903 18173 1912 18207
rect 1860 18164 1912 18173
rect 7656 18164 7708 18216
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 10876 18232 10928 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 13268 18300 13320 18352
rect 15292 18368 15344 18420
rect 15384 18368 15436 18420
rect 17316 18368 17368 18420
rect 13544 18232 13596 18284
rect 15384 18232 15436 18284
rect 16580 18300 16632 18352
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 17776 18232 17828 18284
rect 9956 18164 10008 18216
rect 10416 18164 10468 18216
rect 12072 18164 12124 18216
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 8208 18096 8260 18148
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 12440 18164 12492 18216
rect 12716 18164 12768 18216
rect 12900 18164 12952 18216
rect 13360 18164 13412 18216
rect 15016 18096 15068 18148
rect 15476 18164 15528 18216
rect 4896 18028 4948 18080
rect 6276 18028 6328 18080
rect 6644 18028 6696 18080
rect 7656 18028 7708 18080
rect 9956 18028 10008 18080
rect 11336 18028 11388 18080
rect 12716 18028 12768 18080
rect 15108 18028 15160 18080
rect 15476 18028 15528 18080
rect 16304 18096 16356 18148
rect 21548 18300 21600 18352
rect 22008 18343 22060 18352
rect 22008 18309 22017 18343
rect 22017 18309 22051 18343
rect 22051 18309 22060 18343
rect 22008 18300 22060 18309
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 23388 18368 23440 18420
rect 25412 18368 25464 18420
rect 25780 18368 25832 18420
rect 25228 18343 25280 18352
rect 25228 18309 25237 18343
rect 25237 18309 25271 18343
rect 25271 18309 25280 18343
rect 25228 18300 25280 18309
rect 18696 18232 18748 18284
rect 20720 18232 20772 18284
rect 21180 18232 21232 18284
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 18880 18164 18932 18216
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 19064 18096 19116 18148
rect 19340 18096 19392 18148
rect 20812 18096 20864 18148
rect 24032 18164 24084 18216
rect 21916 18096 21968 18148
rect 26700 18096 26752 18148
rect 16212 18028 16264 18080
rect 16764 18028 16816 18080
rect 17500 18028 17552 18080
rect 19800 18028 19852 18080
rect 21088 18028 21140 18080
rect 22192 18028 22244 18080
rect 22560 18028 22612 18080
rect 23296 18028 23348 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 6920 17824 6972 17876
rect 5908 17756 5960 17808
rect 8668 17756 8720 17808
rect 4160 17688 4212 17740
rect 4436 17688 4488 17740
rect 3976 17620 4028 17672
rect 6736 17688 6788 17740
rect 12624 17824 12676 17876
rect 13452 17824 13504 17876
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 11612 17756 11664 17808
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 6276 17620 6328 17672
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 7656 17620 7708 17672
rect 7840 17620 7892 17672
rect 8944 17620 8996 17672
rect 11704 17688 11756 17740
rect 14464 17756 14516 17808
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 16304 17756 16356 17808
rect 16488 17756 16540 17808
rect 23388 17824 23440 17876
rect 17316 17756 17368 17808
rect 16580 17688 16632 17740
rect 18328 17688 18380 17740
rect 19248 17688 19300 17740
rect 20076 17731 20128 17740
rect 20076 17697 20085 17731
rect 20085 17697 20119 17731
rect 20119 17697 20128 17731
rect 20076 17688 20128 17697
rect 22192 17688 22244 17740
rect 22928 17756 22980 17808
rect 23480 17756 23532 17808
rect 14556 17620 14608 17672
rect 16672 17620 16724 17672
rect 17776 17620 17828 17672
rect 20628 17620 20680 17672
rect 22468 17620 22520 17672
rect 23480 17620 23532 17672
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 1492 17552 1544 17604
rect 5448 17552 5500 17604
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 2780 17484 2832 17493
rect 3884 17484 3936 17536
rect 4160 17484 4212 17536
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 5632 17484 5684 17536
rect 8484 17552 8536 17604
rect 7840 17484 7892 17536
rect 9588 17484 9640 17536
rect 9956 17552 10008 17604
rect 10784 17552 10836 17604
rect 12992 17552 13044 17604
rect 15200 17595 15252 17604
rect 15200 17561 15209 17595
rect 15209 17561 15243 17595
rect 15243 17561 15252 17595
rect 15200 17552 15252 17561
rect 11428 17484 11480 17536
rect 12532 17484 12584 17536
rect 14004 17484 14056 17536
rect 14740 17484 14792 17536
rect 15016 17484 15068 17536
rect 16488 17552 16540 17604
rect 18972 17552 19024 17604
rect 16212 17484 16264 17536
rect 16948 17484 17000 17536
rect 17040 17484 17092 17536
rect 17684 17484 17736 17536
rect 19616 17484 19668 17536
rect 20996 17595 21048 17604
rect 20996 17561 21005 17595
rect 21005 17561 21039 17595
rect 21039 17561 21048 17595
rect 20996 17552 21048 17561
rect 21732 17552 21784 17604
rect 22928 17552 22980 17604
rect 22652 17484 22704 17536
rect 23204 17484 23256 17536
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 23480 17484 23532 17536
rect 24216 17484 24268 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 2136 17280 2188 17332
rect 7012 17280 7064 17332
rect 1768 17212 1820 17264
rect 4252 17212 4304 17264
rect 6920 17212 6972 17264
rect 2044 17144 2096 17196
rect 4620 17144 4672 17196
rect 4988 17144 5040 17196
rect 7196 17280 7248 17332
rect 10784 17212 10836 17264
rect 11428 17212 11480 17264
rect 12624 17280 12676 17332
rect 13728 17280 13780 17332
rect 14096 17323 14148 17332
rect 14096 17289 14105 17323
rect 14105 17289 14139 17323
rect 14139 17289 14148 17323
rect 14096 17280 14148 17289
rect 15200 17280 15252 17332
rect 15476 17280 15528 17332
rect 15844 17323 15896 17332
rect 15844 17289 15853 17323
rect 15853 17289 15887 17323
rect 15887 17289 15896 17323
rect 15844 17280 15896 17289
rect 17224 17280 17276 17332
rect 13544 17212 13596 17264
rect 20168 17212 20220 17264
rect 24584 17280 24636 17332
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 21732 17212 21784 17264
rect 22468 17212 22520 17264
rect 22928 17212 22980 17264
rect 24216 17212 24268 17264
rect 25228 17212 25280 17264
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 4528 17119 4580 17128
rect 4528 17085 4537 17119
rect 4537 17085 4571 17119
rect 4571 17085 4580 17119
rect 4528 17076 4580 17085
rect 8300 17076 8352 17128
rect 7288 17008 7340 17060
rect 3884 16940 3936 16992
rect 6000 16940 6052 16992
rect 8944 17144 8996 17196
rect 10876 17144 10928 17196
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 10048 17076 10100 17128
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 12716 17076 12768 17128
rect 12992 17076 13044 17128
rect 13636 17144 13688 17196
rect 14648 17144 14700 17196
rect 16948 17144 17000 17196
rect 17684 17144 17736 17196
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 14096 17076 14148 17128
rect 11520 17008 11572 17060
rect 13544 17008 13596 17060
rect 16212 17076 16264 17128
rect 16304 17008 16356 17060
rect 17776 17008 17828 17060
rect 11060 16940 11112 16992
rect 13360 16940 13412 16992
rect 14096 16940 14148 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 17868 16983 17920 16992
rect 17868 16949 17877 16983
rect 17877 16949 17911 16983
rect 17911 16949 17920 16983
rect 17868 16940 17920 16949
rect 18972 16940 19024 16992
rect 19248 16940 19300 16992
rect 20260 17144 20312 17196
rect 20628 17144 20680 17196
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 25412 17144 25464 17196
rect 26056 17144 26108 17196
rect 21456 17076 21508 17128
rect 22468 17076 22520 17128
rect 22928 17076 22980 17128
rect 24400 17076 24452 17128
rect 19708 17008 19760 17060
rect 22560 17008 22612 17060
rect 26700 17008 26752 17060
rect 20812 16940 20864 16992
rect 21732 16940 21784 16992
rect 22652 16940 22704 16992
rect 23388 16940 23440 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 2228 16532 2280 16584
rect 6920 16736 6972 16788
rect 7472 16736 7524 16788
rect 9128 16736 9180 16788
rect 9680 16736 9732 16788
rect 10048 16736 10100 16788
rect 11152 16736 11204 16788
rect 3884 16711 3936 16720
rect 3884 16677 3893 16711
rect 3893 16677 3927 16711
rect 3927 16677 3936 16711
rect 3884 16668 3936 16677
rect 4160 16711 4212 16720
rect 4160 16677 4169 16711
rect 4169 16677 4203 16711
rect 4203 16677 4212 16711
rect 4160 16668 4212 16677
rect 3056 16600 3108 16652
rect 6460 16668 6512 16720
rect 9220 16668 9272 16720
rect 10784 16668 10836 16720
rect 5356 16600 5408 16652
rect 5908 16600 5960 16652
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 6552 16600 6604 16652
rect 9404 16600 9456 16652
rect 10600 16600 10652 16652
rect 11060 16600 11112 16652
rect 14096 16736 14148 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 17868 16736 17920 16788
rect 19156 16736 19208 16788
rect 15660 16668 15712 16720
rect 16764 16668 16816 16720
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 14004 16600 14056 16652
rect 14924 16600 14976 16652
rect 19156 16600 19208 16652
rect 19708 16643 19760 16652
rect 19708 16609 19717 16643
rect 19717 16609 19751 16643
rect 19751 16609 19760 16643
rect 19708 16600 19760 16609
rect 5448 16464 5500 16516
rect 2044 16396 2096 16448
rect 5724 16396 5776 16448
rect 6000 16464 6052 16516
rect 7564 16396 7616 16448
rect 8668 16396 8720 16448
rect 8944 16396 8996 16448
rect 9404 16396 9456 16448
rect 9772 16396 9824 16448
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 10876 16396 10928 16448
rect 11704 16532 11756 16584
rect 16764 16532 16816 16584
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 18972 16532 19024 16584
rect 19248 16532 19300 16584
rect 20812 16532 20864 16584
rect 22284 16736 22336 16788
rect 23112 16736 23164 16788
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 25136 16600 25188 16652
rect 26148 16600 26200 16652
rect 12716 16464 12768 16516
rect 14464 16464 14516 16516
rect 15016 16464 15068 16516
rect 17316 16464 17368 16516
rect 17868 16464 17920 16516
rect 12348 16396 12400 16448
rect 14004 16396 14056 16448
rect 16212 16396 16264 16448
rect 19432 16464 19484 16516
rect 20352 16396 20404 16448
rect 20444 16396 20496 16448
rect 24216 16532 24268 16584
rect 21364 16396 21416 16448
rect 22652 16464 22704 16516
rect 24032 16439 24084 16448
rect 24032 16405 24041 16439
rect 24041 16405 24075 16439
rect 24075 16405 24084 16439
rect 24032 16396 24084 16405
rect 25228 16439 25280 16448
rect 25228 16405 25237 16439
rect 25237 16405 25271 16439
rect 25271 16405 25280 16439
rect 25228 16396 25280 16405
rect 25780 16396 25832 16448
rect 25964 16396 26016 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 26056 16328 26108 16380
rect 9128 16192 9180 16244
rect 9496 16192 9548 16244
rect 3516 16124 3568 16176
rect 6644 16167 6696 16176
rect 1860 16099 1912 16108
rect 1860 16065 1869 16099
rect 1869 16065 1903 16099
rect 1903 16065 1912 16099
rect 1860 16056 1912 16065
rect 3424 16056 3476 16108
rect 6644 16133 6653 16167
rect 6653 16133 6687 16167
rect 6687 16133 6696 16167
rect 6644 16124 6696 16133
rect 10876 16192 10928 16244
rect 11244 16192 11296 16244
rect 5356 16056 5408 16108
rect 6368 16056 6420 16108
rect 6552 16056 6604 16108
rect 10324 16124 10376 16176
rect 12716 16124 12768 16176
rect 15292 16124 15344 16176
rect 16396 16124 16448 16176
rect 7196 16056 7248 16108
rect 7564 16056 7616 16108
rect 3332 15988 3384 16040
rect 4160 15920 4212 15972
rect 9036 16056 9088 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 9588 16056 9640 16108
rect 10692 15988 10744 16040
rect 6644 15920 6696 15972
rect 7104 15852 7156 15904
rect 7196 15852 7248 15904
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 11980 15988 12032 16040
rect 14740 16056 14792 16108
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 18972 16056 19024 16108
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 19064 15988 19116 16040
rect 19248 15988 19300 16040
rect 19616 16056 19668 16108
rect 20168 15988 20220 16040
rect 20720 16056 20772 16108
rect 21732 16124 21784 16176
rect 23848 16235 23900 16244
rect 23848 16201 23857 16235
rect 23857 16201 23891 16235
rect 23891 16201 23900 16235
rect 23848 16192 23900 16201
rect 25228 16124 25280 16176
rect 20536 15988 20588 16040
rect 21180 16031 21232 16040
rect 21180 15997 21189 16031
rect 21189 15997 21223 16031
rect 21223 15997 21232 16031
rect 21180 15988 21232 15997
rect 16764 15920 16816 15972
rect 22100 15988 22152 16040
rect 22192 15988 22244 16040
rect 23112 16056 23164 16108
rect 23480 16056 23532 16108
rect 21640 15920 21692 15972
rect 13544 15852 13596 15904
rect 14188 15852 14240 15904
rect 14556 15852 14608 15904
rect 16212 15852 16264 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 20628 15852 20680 15904
rect 22376 15852 22428 15904
rect 24032 16031 24084 16040
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 22652 15920 22704 15972
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 4712 15648 4764 15700
rect 6092 15648 6144 15700
rect 6460 15691 6512 15700
rect 6460 15657 6469 15691
rect 6469 15657 6503 15691
rect 6503 15657 6512 15691
rect 6460 15648 6512 15657
rect 6828 15648 6880 15700
rect 8668 15648 8720 15700
rect 12624 15648 12676 15700
rect 2780 15512 2832 15564
rect 8208 15512 8260 15564
rect 10508 15580 10560 15632
rect 12072 15512 12124 15564
rect 16856 15648 16908 15700
rect 19156 15648 19208 15700
rect 23756 15648 23808 15700
rect 24216 15691 24268 15700
rect 24216 15657 24225 15691
rect 24225 15657 24259 15691
rect 24259 15657 24268 15691
rect 24216 15648 24268 15657
rect 16764 15580 16816 15632
rect 20536 15580 20588 15632
rect 13360 15555 13412 15564
rect 13360 15521 13369 15555
rect 13369 15521 13403 15555
rect 13403 15521 13412 15555
rect 13360 15512 13412 15521
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 16856 15512 16908 15564
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 4436 15444 4488 15496
rect 5540 15444 5592 15496
rect 6000 15487 6052 15496
rect 6000 15453 6009 15487
rect 6009 15453 6043 15487
rect 6043 15453 6052 15487
rect 6000 15444 6052 15453
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 7196 15444 7248 15496
rect 8760 15444 8812 15496
rect 9680 15444 9732 15496
rect 10232 15376 10284 15428
rect 12348 15444 12400 15496
rect 12716 15444 12768 15496
rect 13912 15444 13964 15496
rect 19984 15555 20036 15564
rect 19984 15521 19993 15555
rect 19993 15521 20027 15555
rect 20027 15521 20036 15555
rect 19984 15512 20036 15521
rect 20260 15512 20312 15564
rect 21272 15512 21324 15564
rect 21364 15555 21416 15564
rect 21364 15521 21373 15555
rect 21373 15521 21407 15555
rect 21407 15521 21416 15555
rect 21364 15512 21416 15521
rect 21456 15512 21508 15564
rect 23020 15580 23072 15632
rect 23480 15580 23532 15632
rect 19892 15444 19944 15496
rect 25780 15512 25832 15564
rect 24032 15444 24084 15496
rect 10876 15376 10928 15428
rect 4436 15308 4488 15360
rect 7196 15308 7248 15360
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 9772 15351 9824 15360
rect 9772 15317 9781 15351
rect 9781 15317 9815 15351
rect 9815 15317 9824 15351
rect 9772 15308 9824 15317
rect 10508 15308 10560 15360
rect 11428 15308 11480 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 14556 15419 14608 15428
rect 14556 15385 14565 15419
rect 14565 15385 14599 15419
rect 14599 15385 14608 15419
rect 14556 15376 14608 15385
rect 15016 15376 15068 15428
rect 17224 15376 17276 15428
rect 13636 15308 13688 15360
rect 14648 15308 14700 15360
rect 16212 15308 16264 15360
rect 21272 15376 21324 15428
rect 21824 15376 21876 15428
rect 23296 15376 23348 15428
rect 23480 15376 23532 15428
rect 19156 15308 19208 15360
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 21548 15308 21600 15360
rect 22560 15351 22612 15360
rect 22560 15317 22569 15351
rect 22569 15317 22603 15351
rect 22603 15317 22612 15351
rect 22560 15308 22612 15317
rect 23756 15308 23808 15360
rect 24032 15308 24084 15360
rect 24308 15308 24360 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 1308 15104 1360 15156
rect 2044 15104 2096 15156
rect 3792 15147 3844 15156
rect 3792 15113 3801 15147
rect 3801 15113 3835 15147
rect 3835 15113 3844 15147
rect 3792 15104 3844 15113
rect 4528 15104 4580 15156
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 5540 15079 5592 15088
rect 5540 15045 5549 15079
rect 5549 15045 5583 15079
rect 5583 15045 5592 15079
rect 5540 15036 5592 15045
rect 8576 15104 8628 15156
rect 9220 15147 9272 15156
rect 9220 15113 9229 15147
rect 9229 15113 9263 15147
rect 9263 15113 9272 15147
rect 9220 15104 9272 15113
rect 9956 15104 10008 15156
rect 11060 15104 11112 15156
rect 11888 15104 11940 15156
rect 13636 15104 13688 15156
rect 13820 15104 13872 15156
rect 14556 15104 14608 15156
rect 7840 15036 7892 15088
rect 3700 14900 3752 14952
rect 4344 14943 4396 14952
rect 4344 14909 4353 14943
rect 4353 14909 4387 14943
rect 4387 14909 4396 14943
rect 4344 14900 4396 14909
rect 6552 14943 6604 14952
rect 6552 14909 6561 14943
rect 6561 14909 6595 14943
rect 6595 14909 6604 14943
rect 6552 14900 6604 14909
rect 8300 14900 8352 14952
rect 8760 15011 8812 15020
rect 8760 14977 8769 15011
rect 8769 14977 8803 15011
rect 8803 14977 8812 15011
rect 8760 14968 8812 14977
rect 9220 14968 9272 15020
rect 9864 14968 9916 15020
rect 10140 14900 10192 14952
rect 10324 15036 10376 15088
rect 11612 15036 11664 15088
rect 12256 15036 12308 15088
rect 12624 15036 12676 15088
rect 15016 15036 15068 15088
rect 16212 15036 16264 15088
rect 17224 15036 17276 15088
rect 18972 15147 19024 15156
rect 18972 15113 18981 15147
rect 18981 15113 19015 15147
rect 19015 15113 19024 15147
rect 18972 15104 19024 15113
rect 22560 15104 22612 15156
rect 22008 15036 22060 15088
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 23020 15104 23072 15156
rect 23296 15104 23348 15156
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 10876 14968 10928 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 16580 14968 16632 15020
rect 16764 14968 16816 15020
rect 20720 14968 20772 15020
rect 6736 14832 6788 14884
rect 7564 14832 7616 14884
rect 8300 14764 8352 14816
rect 8576 14807 8628 14816
rect 8576 14773 8585 14807
rect 8585 14773 8619 14807
rect 8619 14773 8628 14807
rect 8576 14764 8628 14773
rect 10968 14764 11020 14816
rect 13636 14832 13688 14884
rect 15384 14832 15436 14884
rect 17868 14900 17920 14952
rect 19340 14943 19392 14952
rect 13728 14764 13780 14816
rect 14556 14764 14608 14816
rect 15200 14807 15252 14816
rect 15200 14773 15209 14807
rect 15209 14773 15243 14807
rect 15243 14773 15252 14807
rect 15200 14764 15252 14773
rect 16764 14764 16816 14816
rect 17132 14764 17184 14816
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 19248 14832 19300 14884
rect 23756 15036 23808 15088
rect 22284 14968 22336 15020
rect 24308 14900 24360 14952
rect 24492 14900 24544 14952
rect 22836 14832 22888 14884
rect 18880 14764 18932 14816
rect 21824 14764 21876 14816
rect 23756 14764 23808 14816
rect 25228 14807 25280 14816
rect 25228 14773 25237 14807
rect 25237 14773 25271 14807
rect 25271 14773 25280 14807
rect 25228 14764 25280 14773
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 2780 14560 2832 14612
rect 4252 14560 4304 14612
rect 4620 14560 4672 14612
rect 4804 14560 4856 14612
rect 6460 14560 6512 14612
rect 6552 14560 6604 14612
rect 5632 14492 5684 14544
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3516 14356 3568 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 7748 14492 7800 14544
rect 7840 14535 7892 14544
rect 7840 14501 7849 14535
rect 7849 14501 7883 14535
rect 7883 14501 7892 14535
rect 7840 14492 7892 14501
rect 8392 14492 8444 14544
rect 10416 14492 10468 14544
rect 6092 14424 6144 14476
rect 9956 14424 10008 14476
rect 12072 14560 12124 14612
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 7840 14356 7892 14408
rect 8852 14356 8904 14408
rect 10968 14467 11020 14476
rect 10968 14433 10977 14467
rect 10977 14433 11011 14467
rect 11011 14433 11020 14467
rect 10968 14424 11020 14433
rect 12624 14492 12676 14544
rect 16028 14560 16080 14612
rect 13820 14535 13872 14544
rect 13820 14501 13829 14535
rect 13829 14501 13863 14535
rect 13863 14501 13872 14535
rect 13820 14492 13872 14501
rect 14096 14424 14148 14476
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16764 14560 16816 14612
rect 18604 14560 18656 14612
rect 19524 14560 19576 14612
rect 20720 14560 20772 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 22836 14560 22888 14612
rect 19248 14492 19300 14544
rect 16488 14424 16540 14433
rect 17776 14424 17828 14476
rect 19800 14424 19852 14476
rect 20352 14492 20404 14544
rect 23388 14492 23440 14544
rect 20260 14424 20312 14476
rect 26148 14492 26200 14544
rect 23572 14424 23624 14476
rect 24492 14424 24544 14476
rect 10324 14356 10376 14408
rect 9680 14288 9732 14340
rect 12072 14356 12124 14408
rect 12348 14356 12400 14408
rect 13544 14356 13596 14408
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 19064 14356 19116 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 22008 14356 22060 14408
rect 10876 14288 10928 14340
rect 3424 14220 3476 14272
rect 5264 14220 5316 14272
rect 5448 14220 5500 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 7288 14220 7340 14229
rect 7748 14220 7800 14272
rect 9864 14220 9916 14272
rect 11152 14220 11204 14272
rect 13820 14220 13872 14272
rect 14556 14220 14608 14272
rect 15016 14288 15068 14340
rect 16580 14220 16632 14272
rect 17224 14288 17276 14340
rect 21364 14288 21416 14340
rect 21640 14288 21692 14340
rect 24032 14288 24084 14340
rect 24216 14288 24268 14340
rect 19340 14220 19392 14272
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 22836 14220 22888 14272
rect 23572 14220 23624 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 2320 14016 2372 14068
rect 4068 14016 4120 14068
rect 4804 14016 4856 14068
rect 5540 14016 5592 14068
rect 6092 14016 6144 14068
rect 6828 14016 6880 14068
rect 8484 14016 8536 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 10232 14016 10284 14068
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 3424 13923 3476 13932
rect 3424 13889 3433 13923
rect 3433 13889 3467 13923
rect 3467 13889 3476 13923
rect 3424 13880 3476 13889
rect 4160 13812 4212 13864
rect 7012 13948 7064 14000
rect 6092 13880 6144 13932
rect 7104 13880 7156 13932
rect 7656 13948 7708 14000
rect 7932 13948 7984 14000
rect 10140 13948 10192 14000
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 11060 13880 11112 13932
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 7564 13812 7616 13864
rect 11336 13812 11388 13864
rect 12072 13948 12124 14000
rect 12256 14016 12308 14068
rect 14188 14016 14240 14068
rect 16212 14016 16264 14068
rect 17224 14016 17276 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 17868 14016 17920 14068
rect 13636 13948 13688 14000
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 14280 13948 14332 14000
rect 14556 13948 14608 14000
rect 16028 13948 16080 14000
rect 15292 13880 15344 13932
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 18420 13948 18472 14000
rect 19064 13948 19116 14000
rect 19432 14016 19484 14068
rect 20812 14016 20864 14068
rect 21088 14016 21140 14068
rect 21364 14016 21416 14068
rect 24676 14016 24728 14068
rect 25044 14016 25096 14068
rect 25596 14016 25648 14068
rect 21456 13948 21508 14000
rect 23388 13948 23440 14000
rect 24952 13991 25004 14000
rect 24952 13957 24961 13991
rect 24961 13957 24995 13991
rect 24995 13957 25004 13991
rect 24952 13948 25004 13957
rect 25872 13948 25924 14000
rect 13544 13812 13596 13864
rect 7748 13744 7800 13796
rect 1584 13676 1636 13728
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 11060 13676 11112 13728
rect 11612 13676 11664 13728
rect 11796 13744 11848 13796
rect 16028 13812 16080 13864
rect 16212 13812 16264 13864
rect 17040 13787 17092 13796
rect 17040 13753 17049 13787
rect 17049 13753 17083 13787
rect 17083 13753 17092 13787
rect 17040 13744 17092 13753
rect 17500 13744 17552 13796
rect 17868 13812 17920 13864
rect 21640 13812 21692 13864
rect 22192 13812 22244 13864
rect 24216 13880 24268 13932
rect 25964 13880 26016 13932
rect 12440 13676 12492 13728
rect 15384 13676 15436 13728
rect 16764 13676 16816 13728
rect 18512 13676 18564 13728
rect 19248 13676 19300 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 24492 13812 24544 13864
rect 25596 13812 25648 13864
rect 25688 13812 25740 13864
rect 25872 13812 25924 13864
rect 21732 13676 21784 13728
rect 24952 13744 25004 13796
rect 22928 13676 22980 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 3148 13472 3200 13524
rect 5908 13472 5960 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 9128 13472 9180 13524
rect 11796 13472 11848 13524
rect 5448 13404 5500 13456
rect 8300 13404 8352 13456
rect 14004 13472 14056 13524
rect 15200 13472 15252 13524
rect 15568 13472 15620 13524
rect 16028 13472 16080 13524
rect 17500 13472 17552 13524
rect 2136 13379 2188 13388
rect 2136 13345 2145 13379
rect 2145 13345 2179 13379
rect 2179 13345 2188 13379
rect 2136 13336 2188 13345
rect 9680 13336 9732 13388
rect 10876 13336 10928 13388
rect 13820 13379 13872 13388
rect 13820 13345 13829 13379
rect 13829 13345 13863 13379
rect 13863 13345 13872 13379
rect 13820 13336 13872 13345
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 9404 13200 9456 13252
rect 11612 13200 11664 13252
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 10048 13132 10100 13184
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12072 13243 12124 13252
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 13728 13200 13780 13252
rect 15016 13200 15068 13252
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 18328 13336 18380 13388
rect 16764 13200 16816 13252
rect 17224 13200 17276 13252
rect 15200 13132 15252 13184
rect 15568 13132 15620 13184
rect 20168 13472 20220 13524
rect 21640 13472 21692 13524
rect 23940 13472 23992 13524
rect 24124 13472 24176 13524
rect 24400 13472 24452 13524
rect 18788 13336 18840 13388
rect 21916 13379 21968 13388
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22652 13336 22704 13388
rect 22928 13336 22980 13388
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 24216 13447 24268 13456
rect 24216 13413 24225 13447
rect 24225 13413 24259 13447
rect 24259 13413 24268 13447
rect 24216 13404 24268 13413
rect 23756 13336 23808 13388
rect 19984 13243 20036 13252
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 21640 13200 21692 13252
rect 25412 13268 25464 13320
rect 25872 13200 25924 13252
rect 24216 13132 24268 13184
rect 25320 13132 25372 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 2504 12928 2556 12980
rect 3148 12928 3200 12980
rect 8300 12860 8352 12912
rect 10600 12971 10652 12980
rect 10600 12937 10609 12971
rect 10609 12937 10643 12971
rect 10643 12937 10652 12971
rect 10600 12928 10652 12937
rect 11152 12928 11204 12980
rect 12072 12928 12124 12980
rect 13820 12928 13872 12980
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 11244 12860 11296 12912
rect 11612 12860 11664 12912
rect 18420 12928 18472 12980
rect 18604 12928 18656 12980
rect 19800 12928 19852 12980
rect 15384 12860 15436 12912
rect 16488 12860 16540 12912
rect 17224 12860 17276 12912
rect 19984 12928 20036 12980
rect 25136 12928 25188 12980
rect 25320 12928 25372 12980
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 7196 12792 7248 12844
rect 11704 12792 11756 12844
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 12348 12792 12400 12844
rect 13452 12792 13504 12844
rect 15016 12792 15068 12844
rect 15568 12792 15620 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 3424 12724 3476 12776
rect 12716 12724 12768 12776
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 17224 12724 17276 12776
rect 17684 12724 17736 12776
rect 18604 12792 18656 12844
rect 11060 12656 11112 12708
rect 11704 12656 11756 12708
rect 15752 12656 15804 12708
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 15568 12588 15620 12640
rect 19248 12724 19300 12776
rect 20536 12792 20588 12844
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 22560 12860 22612 12912
rect 21916 12792 21968 12844
rect 23940 12792 23992 12844
rect 24308 12792 24360 12844
rect 18420 12656 18472 12708
rect 20536 12656 20588 12708
rect 20996 12724 21048 12776
rect 21364 12724 21416 12776
rect 21456 12724 21508 12776
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 23756 12767 23808 12776
rect 23756 12733 23765 12767
rect 23765 12733 23799 12767
rect 23799 12733 23808 12767
rect 23756 12724 23808 12733
rect 23388 12656 23440 12708
rect 23848 12656 23900 12708
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 19524 12588 19576 12640
rect 21640 12588 21692 12640
rect 22100 12588 22152 12640
rect 22652 12588 22704 12640
rect 23020 12588 23072 12640
rect 23940 12588 23992 12640
rect 25688 12588 25740 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 11612 12384 11664 12436
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 6920 12316 6972 12368
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 18236 12316 18288 12368
rect 20996 12384 21048 12436
rect 23296 12384 23348 12436
rect 25320 12384 25372 12436
rect 7472 12248 7524 12300
rect 15476 12248 15528 12300
rect 16764 12248 16816 12300
rect 17684 12248 17736 12300
rect 19432 12291 19484 12300
rect 19432 12257 19441 12291
rect 19441 12257 19475 12291
rect 19475 12257 19484 12291
rect 19432 12248 19484 12257
rect 21824 12316 21876 12368
rect 11888 12180 11940 12232
rect 12348 12180 12400 12232
rect 13360 12180 13412 12232
rect 13728 12180 13780 12232
rect 14004 12180 14056 12232
rect 18512 12180 18564 12232
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 9864 12044 9916 12096
rect 12532 12044 12584 12096
rect 14464 12112 14516 12164
rect 15476 12112 15528 12164
rect 16304 12112 16356 12164
rect 16488 12112 16540 12164
rect 17868 12112 17920 12164
rect 19984 12112 20036 12164
rect 20444 12112 20496 12164
rect 21364 12248 21416 12300
rect 21916 12248 21968 12300
rect 21088 12180 21140 12232
rect 24124 12180 24176 12232
rect 25228 12180 25280 12232
rect 13084 12044 13136 12096
rect 17316 12044 17368 12096
rect 17592 12044 17644 12096
rect 18512 12044 18564 12096
rect 19064 12044 19116 12096
rect 19432 12044 19484 12096
rect 20076 12044 20128 12096
rect 20536 12044 20588 12096
rect 23848 12112 23900 12164
rect 24308 12112 24360 12164
rect 22652 12044 22704 12096
rect 23388 12044 23440 12096
rect 23940 12044 23992 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12256 11883 12308 11892
rect 12256 11849 12265 11883
rect 12265 11849 12299 11883
rect 12299 11849 12308 11883
rect 12256 11840 12308 11849
rect 13820 11840 13872 11892
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 13084 11815 13136 11824
rect 13084 11781 13093 11815
rect 13093 11781 13127 11815
rect 13127 11781 13136 11815
rect 13084 11772 13136 11781
rect 15016 11772 15068 11824
rect 19432 11840 19484 11892
rect 20444 11840 20496 11892
rect 13544 11636 13596 11688
rect 13728 11636 13780 11688
rect 15108 11636 15160 11688
rect 16396 11636 16448 11688
rect 17868 11772 17920 11824
rect 19708 11772 19760 11824
rect 22100 11840 22152 11892
rect 26240 11840 26292 11892
rect 21640 11772 21692 11824
rect 24860 11772 24912 11824
rect 25136 11815 25188 11824
rect 25136 11781 25145 11815
rect 25145 11781 25179 11815
rect 25179 11781 25188 11815
rect 25136 11772 25188 11781
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 16948 11636 17000 11688
rect 16488 11568 16540 11620
rect 16580 11568 16632 11620
rect 19064 11636 19116 11688
rect 21180 11636 21232 11688
rect 22744 11636 22796 11688
rect 18880 11500 18932 11552
rect 21824 11568 21876 11620
rect 21088 11500 21140 11552
rect 21640 11543 21692 11552
rect 21640 11509 21649 11543
rect 21649 11509 21683 11543
rect 21683 11509 21692 11543
rect 21640 11500 21692 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 4436 11296 4488 11348
rect 22100 11296 22152 11348
rect 12440 11228 12492 11280
rect 14372 11228 14424 11280
rect 15292 11228 15344 11280
rect 15384 11271 15436 11280
rect 15384 11237 15393 11271
rect 15393 11237 15427 11271
rect 15427 11237 15436 11271
rect 15384 11228 15436 11237
rect 16304 11271 16356 11280
rect 16304 11237 16313 11271
rect 16313 11237 16347 11271
rect 16347 11237 16356 11271
rect 16304 11228 16356 11237
rect 17224 11228 17276 11280
rect 18328 11228 18380 11280
rect 12532 11160 12584 11212
rect 18696 11160 18748 11212
rect 19984 11228 20036 11280
rect 21180 11271 21232 11280
rect 21180 11237 21189 11271
rect 21189 11237 21223 11271
rect 21223 11237 21232 11271
rect 21180 11228 21232 11237
rect 21640 11228 21692 11280
rect 22652 11296 22704 11348
rect 23848 11296 23900 11348
rect 25044 11296 25096 11348
rect 20260 11160 20312 11212
rect 20812 11160 20864 11212
rect 20996 11160 21048 11212
rect 24860 11160 24912 11212
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 16028 11092 16080 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 19984 11092 20036 11144
rect 4068 10956 4120 11008
rect 11704 10956 11756 11008
rect 14924 10999 14976 11008
rect 14924 10965 14933 10999
rect 14933 10965 14967 10999
rect 14967 10965 14976 10999
rect 14924 10956 14976 10965
rect 17684 11024 17736 11076
rect 18328 11067 18380 11076
rect 18328 11033 18337 11067
rect 18337 11033 18371 11067
rect 18371 11033 18380 11067
rect 18328 11024 18380 11033
rect 20076 11024 20128 11076
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 22744 11135 22796 11144
rect 22744 11101 22753 11135
rect 22753 11101 22787 11135
rect 22787 11101 22796 11135
rect 22744 11092 22796 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 21824 11024 21876 11076
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 21916 11024 21968 11033
rect 16580 10956 16632 11008
rect 19708 10956 19760 11008
rect 23388 11024 23440 11076
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 13820 10752 13872 10804
rect 14924 10752 14976 10804
rect 16672 10752 16724 10804
rect 16856 10752 16908 10804
rect 17132 10752 17184 10804
rect 19064 10795 19116 10804
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 22284 10752 22336 10804
rect 11704 10684 11756 10736
rect 14464 10548 14516 10600
rect 16856 10616 16908 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 18328 10548 18380 10600
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 21548 10616 21600 10668
rect 22284 10616 22336 10668
rect 22560 10616 22612 10668
rect 24860 10684 24912 10736
rect 15568 10480 15620 10532
rect 16488 10480 16540 10532
rect 16948 10412 17000 10464
rect 17132 10412 17184 10464
rect 18420 10480 18472 10532
rect 19064 10480 19116 10532
rect 19340 10480 19392 10532
rect 19708 10480 19760 10532
rect 22376 10548 22428 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 22008 10480 22060 10532
rect 20168 10412 20220 10464
rect 20260 10412 20312 10464
rect 26516 10480 26568 10532
rect 22560 10412 22612 10464
rect 23296 10412 23348 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 14832 10208 14884 10260
rect 15200 10208 15252 10260
rect 17224 10208 17276 10260
rect 17592 10251 17644 10260
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 18420 10208 18472 10260
rect 19616 10208 19668 10260
rect 22376 10208 22428 10260
rect 10968 10072 11020 10124
rect 16396 10072 16448 10124
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 16488 10004 16540 10056
rect 16672 10004 16724 10056
rect 17132 10004 17184 10056
rect 17408 10072 17460 10124
rect 20996 10072 21048 10124
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 23204 10140 23256 10192
rect 12808 9868 12860 9920
rect 16672 9868 16724 9920
rect 17592 9868 17644 9920
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 25780 10004 25832 10056
rect 20352 9936 20404 9988
rect 21640 9979 21692 9988
rect 21640 9945 21649 9979
rect 21649 9945 21683 9979
rect 21683 9945 21692 9979
rect 21640 9936 21692 9945
rect 22652 9936 22704 9988
rect 23388 9936 23440 9988
rect 21548 9868 21600 9920
rect 23204 9868 23256 9920
rect 23940 9911 23992 9920
rect 23940 9877 23949 9911
rect 23949 9877 23983 9911
rect 23983 9877 23992 9911
rect 23940 9868 23992 9877
rect 24584 9911 24636 9920
rect 24584 9877 24593 9911
rect 24593 9877 24627 9911
rect 24627 9877 24636 9911
rect 24584 9868 24636 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 14648 9664 14700 9716
rect 15292 9664 15344 9716
rect 16948 9664 17000 9716
rect 19616 9664 19668 9716
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 15660 9639 15712 9648
rect 15660 9605 15669 9639
rect 15669 9605 15703 9639
rect 15703 9605 15712 9639
rect 15660 9596 15712 9605
rect 18604 9596 18656 9648
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 20904 9596 20956 9648
rect 22100 9664 22152 9716
rect 22652 9664 22704 9716
rect 21088 9596 21140 9648
rect 22008 9596 22060 9648
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 23480 9596 23532 9648
rect 23848 9596 23900 9648
rect 25136 9639 25188 9648
rect 25136 9605 25145 9639
rect 25145 9605 25179 9639
rect 25179 9605 25188 9639
rect 25136 9596 25188 9605
rect 20352 9528 20404 9580
rect 21180 9528 21232 9580
rect 21548 9528 21600 9580
rect 22468 9528 22520 9580
rect 15016 9392 15068 9444
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 19800 9392 19852 9444
rect 20536 9435 20588 9444
rect 20536 9401 20545 9435
rect 20545 9401 20579 9435
rect 20579 9401 20588 9435
rect 20536 9392 20588 9401
rect 21732 9460 21784 9512
rect 24032 9460 24084 9512
rect 22008 9392 22060 9444
rect 22100 9392 22152 9444
rect 26884 9392 26936 9444
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 19340 9324 19392 9376
rect 22376 9324 22428 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 25964 9188 26016 9240
rect 26608 9188 26660 9240
rect 11888 9120 11940 9172
rect 15844 9120 15896 9172
rect 8576 9052 8628 9104
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 19156 9120 19208 9172
rect 21548 9120 21600 9172
rect 21640 9120 21692 9172
rect 25412 9120 25464 9172
rect 18696 9052 18748 9104
rect 6828 8848 6880 8900
rect 13820 8848 13872 8900
rect 20168 8984 20220 9036
rect 19432 8916 19484 8968
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 19984 8848 20036 8900
rect 20812 8959 20864 8968
rect 20812 8925 20821 8959
rect 20821 8925 20855 8959
rect 20855 8925 20864 8959
rect 20812 8916 20864 8925
rect 22836 8984 22888 9036
rect 24860 8984 24912 9036
rect 21548 8916 21600 8968
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 23756 8916 23808 8968
rect 20996 8848 21048 8900
rect 26332 8848 26384 8900
rect 18420 8780 18472 8832
rect 18788 8780 18840 8832
rect 20168 8780 20220 8832
rect 22560 8780 22612 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 16580 8508 16632 8560
rect 19800 8619 19852 8628
rect 19800 8585 19809 8619
rect 19809 8585 19843 8619
rect 19843 8585 19852 8619
rect 19800 8576 19852 8585
rect 20812 8576 20864 8628
rect 21272 8619 21324 8628
rect 21272 8585 21281 8619
rect 21281 8585 21315 8619
rect 21315 8585 21324 8619
rect 21272 8576 21324 8585
rect 21364 8576 21416 8628
rect 22100 8576 22152 8628
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 18880 8372 18932 8424
rect 20260 8440 20312 8492
rect 20444 8440 20496 8492
rect 19064 8372 19116 8424
rect 26700 8576 26752 8628
rect 20444 8347 20496 8356
rect 20444 8313 20453 8347
rect 20453 8313 20487 8347
rect 20487 8313 20496 8347
rect 20444 8304 20496 8313
rect 21364 8304 21416 8356
rect 24952 8440 25004 8492
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 24216 8304 24268 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 20168 8032 20220 8084
rect 20904 8032 20956 8084
rect 17500 7896 17552 7948
rect 22192 7964 22244 8016
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 26424 7964 26476 8016
rect 23480 7896 23532 7948
rect 24860 7896 24912 7948
rect 20628 7828 20680 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 22376 7828 22428 7880
rect 24492 7828 24544 7880
rect 23388 7760 23440 7812
rect 20812 7692 20864 7744
rect 21088 7692 21140 7744
rect 22192 7692 22244 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 17868 7488 17920 7540
rect 18328 7488 18380 7540
rect 22652 7488 22704 7540
rect 18420 7420 18472 7472
rect 23756 7488 23808 7540
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 24860 7420 24912 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 19708 7352 19760 7404
rect 19340 7284 19392 7336
rect 20720 7352 20772 7404
rect 16212 7216 16264 7268
rect 23480 7352 23532 7404
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 25044 7148 25096 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 6276 6808 6328 6860
rect 17224 6808 17276 6860
rect 22468 6808 22520 6860
rect 24492 6851 24544 6860
rect 24492 6817 24501 6851
rect 24501 6817 24535 6851
rect 24535 6817 24544 6851
rect 24492 6808 24544 6817
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 19248 6740 19300 6792
rect 20628 6740 20680 6792
rect 21272 6740 21324 6792
rect 24952 6740 25004 6792
rect 16120 6604 16172 6656
rect 21456 6715 21508 6724
rect 21456 6681 21465 6715
rect 21465 6681 21499 6715
rect 21499 6681 21508 6715
rect 21456 6672 21508 6681
rect 21732 6672 21784 6724
rect 21824 6672 21876 6724
rect 25228 6740 25280 6792
rect 25320 6715 25372 6724
rect 25320 6681 25329 6715
rect 25329 6681 25363 6715
rect 25363 6681 25372 6715
rect 25320 6672 25372 6681
rect 21180 6647 21232 6656
rect 21180 6613 21189 6647
rect 21189 6613 21223 6647
rect 21223 6613 21232 6647
rect 21180 6604 21232 6613
rect 22100 6647 22152 6656
rect 22100 6613 22109 6647
rect 22109 6613 22143 6647
rect 22143 6613 22152 6647
rect 22100 6604 22152 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 19248 6400 19300 6452
rect 20260 6400 20312 6452
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 21272 6443 21324 6452
rect 21272 6409 21281 6443
rect 21281 6409 21315 6443
rect 21315 6409 21324 6443
rect 21272 6400 21324 6409
rect 16856 6332 16908 6384
rect 21824 6332 21876 6384
rect 20444 6264 20496 6316
rect 25504 6400 25556 6452
rect 24860 6332 24912 6384
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 23848 6264 23900 6316
rect 17224 6196 17276 6248
rect 23480 6128 23532 6180
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 25228 6128 25280 6180
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 25688 5856 25740 5908
rect 23388 5788 23440 5840
rect 25412 5788 25464 5840
rect 26792 5788 26844 5840
rect 18512 5720 18564 5772
rect 19524 5652 19576 5704
rect 25872 5720 25924 5772
rect 22744 5584 22796 5636
rect 25044 5652 25096 5704
rect 24952 5584 25004 5636
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 24584 5312 24636 5364
rect 24860 5244 24912 5296
rect 22284 5219 22336 5228
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 23756 5176 23808 5228
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 24584 4972 24636 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 15936 4768 15988 4820
rect 25688 4768 25740 4820
rect 25964 4700 26016 4752
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 25136 4632 25188 4684
rect 23388 4564 23440 4616
rect 25504 4496 25556 4548
rect 24676 4471 24728 4480
rect 24676 4437 24685 4471
rect 24685 4437 24719 4471
rect 24719 4437 24728 4471
rect 24676 4428 24728 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18972 4020 19024 4072
rect 20168 4020 20220 4072
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 23664 4088 23716 4140
rect 22192 4020 22244 4072
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 25596 3884 25648 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 25228 3723 25280 3732
rect 25228 3689 25237 3723
rect 25237 3689 25271 3723
rect 25271 3689 25280 3723
rect 25228 3680 25280 3689
rect 22744 3544 22796 3596
rect 21916 3476 21968 3528
rect 24676 3476 24728 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24952 3408 25004 3460
rect 22284 3340 22336 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 25320 3136 25372 3188
rect 24860 3068 24912 3120
rect 25136 3111 25188 3120
rect 25136 3077 25145 3111
rect 25145 3077 25179 3111
rect 25179 3077 25188 3111
rect 25136 3068 25188 3077
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 25044 2932 25096 2984
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 6828 2635 6880 2644
rect 6828 2601 6837 2635
rect 6837 2601 6871 2635
rect 6871 2601 6880 2635
rect 6828 2592 6880 2601
rect 19432 2592 19484 2644
rect 22100 2592 22152 2644
rect 6920 2388 6972 2440
rect 23296 2524 23348 2576
rect 23388 2456 23440 2508
rect 24584 2388 24636 2440
rect 24952 2320 25004 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 2042 26330 2098 27000
rect 2042 26302 2360 26330
rect 2042 26200 2098 26302
rect 2134 26208 2190 26217
rect 1490 24848 1546 24857
rect 1490 24783 1546 24792
rect 1308 22432 1360 22438
rect 1308 22374 1360 22380
rect 1320 15162 1348 22374
rect 1504 22098 1532 24783
rect 1582 23080 1638 23089
rect 1582 23015 1584 23024
rect 1636 23015 1638 23024
rect 1584 22986 1636 22992
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1596 21690 1624 22986
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 19718 1440 20742
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1492 20052 1544 20058
rect 1492 19994 1544 20000
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1412 19394 1440 19654
rect 1504 19514 1532 19994
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1412 19366 1532 19394
rect 1504 18630 1532 19366
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 17610 1532 18566
rect 1492 17604 1544 17610
rect 1492 17546 1544 17552
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1596 13734 1624 20334
rect 1688 19310 1716 26200
rect 2134 26143 2190 26152
rect 2042 23896 2098 23905
rect 2042 23831 2098 23840
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1780 22710 1808 22918
rect 1768 22704 1820 22710
rect 1768 22646 1820 22652
rect 1860 22160 1912 22166
rect 1860 22102 1912 22108
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 21146 1808 21490
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1780 17270 1808 21082
rect 1872 20466 1900 22102
rect 1964 21622 1992 23598
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 1952 20868 2004 20874
rect 1952 20810 2004 20816
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1964 19718 1992 20810
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1768 17264 1820 17270
rect 1768 17206 1820 17212
rect 1872 16574 1900 18158
rect 2056 17202 2084 23831
rect 2148 19854 2176 26143
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22778 2268 23054
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2134 18864 2190 18873
rect 2134 18799 2190 18808
rect 2148 18766 2176 18799
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 17338 2176 18702
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1780 16546 1900 16574
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1780 9625 1808 16546
rect 1858 16144 1914 16153
rect 1858 16079 1860 16088
rect 1912 16079 1914 16088
rect 1860 16050 1912 16056
rect 1964 15178 1992 17070
rect 2240 16590 2268 22170
rect 2332 19922 2360 26302
rect 2410 26200 2466 27000
rect 2502 26208 2558 26217
rect 2424 20942 2452 26200
rect 2778 26200 2834 27000
rect 3146 26330 3202 27000
rect 2884 26302 3202 26330
rect 2502 26143 2558 26152
rect 2516 22234 2544 26143
rect 2688 24132 2740 24138
rect 2688 24074 2740 24080
rect 2700 22982 2728 24074
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2504 22024 2556 22030
rect 2504 21966 2556 21972
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2228 16584 2280 16590
rect 2042 16552 2098 16561
rect 2228 16526 2280 16532
rect 2042 16487 2098 16496
rect 2056 16454 2084 16487
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1964 15162 2084 15178
rect 1964 15156 2096 15162
rect 1964 15150 2044 15156
rect 2044 15098 2096 15104
rect 2318 14512 2374 14521
rect 2318 14447 2374 14456
rect 2332 14414 2360 14447
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 14074 2360 14350
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2318 13968 2374 13977
rect 2318 13903 2320 13912
rect 2372 13903 2374 13912
rect 2320 13874 2372 13880
rect 2134 13424 2190 13433
rect 2134 13359 2136 13368
rect 2188 13359 2190 13368
rect 2136 13330 2188 13336
rect 2516 12986 2544 21966
rect 2608 18970 2636 21966
rect 2700 20806 2728 22918
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2792 20398 2820 26200
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 3514 26200 3570 27000
rect 3608 26308 3660 26314
rect 3608 26250 3660 26256
rect 3146 25936 3202 25945
rect 3146 25871 3202 25880
rect 3160 25702 3188 25871
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 2962 24168 3018 24177
rect 2962 24103 3018 24112
rect 2976 23730 3004 24103
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2872 21616 2924 21622
rect 2872 21558 2924 21564
rect 2884 21418 2912 21558
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2792 17898 2820 18838
rect 2700 17870 2820 17898
rect 2700 16674 2728 17870
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17105 2820 17478
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2884 16674 2912 21354
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3344 18834 3372 24346
rect 3528 21486 3556 26200
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3514 21312 3570 21321
rect 3514 21247 3570 21256
rect 3424 19780 3476 19786
rect 3424 19722 3476 19728
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3068 18290 3096 18566
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3436 18170 3464 19722
rect 3344 18142 3464 18170
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2700 16646 2820 16674
rect 2884 16658 3096 16674
rect 2884 16652 3108 16658
rect 2884 16646 3056 16652
rect 2792 15570 2820 16646
rect 3056 16594 3108 16600
rect 3344 16046 3372 18142
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3436 16114 3464 18022
rect 3528 16182 3556 21247
rect 3620 18630 3648 26250
rect 3700 26240 3752 26246
rect 3882 26200 3938 27000
rect 4250 26200 4306 27000
rect 4618 26200 4674 27000
rect 4986 26330 5042 27000
rect 4986 26302 5120 26330
rect 4986 26200 5042 26302
rect 3700 26182 3752 26188
rect 3712 23066 3740 26182
rect 3792 25356 3844 25362
rect 3792 25298 3844 25304
rect 3804 23202 3832 25298
rect 3896 23322 3924 26200
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 3976 24676 4028 24682
rect 3976 24618 4028 24624
rect 3988 23633 4016 24618
rect 4080 24410 4108 25434
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 4172 24206 4200 24550
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 3974 23624 4030 23633
rect 3974 23559 4030 23568
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 3804 23174 3924 23202
rect 3712 23038 3832 23066
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3712 22001 3740 22646
rect 3698 21992 3754 22001
rect 3698 21927 3754 21936
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3712 21554 3740 21830
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3698 20768 3754 20777
rect 3698 20703 3754 20712
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2778 15056 2834 15065
rect 2778 14991 2780 15000
rect 2832 14991 2834 15000
rect 2780 14962 2832 14968
rect 2792 14618 2820 14962
rect 3712 14958 3740 20703
rect 3804 19786 3832 23038
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 3896 19666 3924 23174
rect 3974 22672 4030 22681
rect 3974 22607 4030 22616
rect 3988 22234 4016 22607
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3988 21690 4016 21898
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3804 19638 3924 19666
rect 3804 18902 3832 19638
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3896 19417 3924 19450
rect 3882 19408 3938 19417
rect 3882 19343 3938 19352
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3792 18896 3844 18902
rect 3792 18838 3844 18844
rect 3896 17542 3924 19246
rect 3988 18834 4016 20198
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3896 16726 3924 16934
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3790 15192 3846 15201
rect 3790 15127 3792 15136
rect 3844 15127 3846 15136
rect 3792 15098 3844 15104
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 13938 3464 14214
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3160 12986 3188 13466
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2134 12880 2190 12889
rect 2134 12815 2136 12824
rect 2188 12815 2190 12824
rect 2136 12786 2188 12792
rect 3436 12782 3464 13262
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3528 12345 3556 14350
rect 3514 12336 3570 12345
rect 3514 12271 3570 12280
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11665 1992 12038
rect 1950 11656 2006 11665
rect 1950 11591 2006 11600
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3988 10713 4016 17614
rect 4080 14414 4108 24006
rect 4172 22522 4200 24006
rect 4264 22710 4292 26200
rect 4434 23624 4490 23633
rect 4434 23559 4490 23568
rect 4342 23216 4398 23225
rect 4342 23151 4398 23160
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4172 22494 4292 22522
rect 4158 22128 4214 22137
rect 4158 22063 4214 22072
rect 4172 20058 4200 22063
rect 4264 22001 4292 22494
rect 4250 21992 4306 22001
rect 4250 21927 4306 21936
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4264 20942 4292 21830
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4172 17746 4200 19450
rect 4356 19446 4384 23151
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4264 17542 4292 19314
rect 4342 18320 4398 18329
rect 4342 18255 4344 18264
rect 4396 18255 4398 18264
rect 4344 18226 4396 18232
rect 4448 17746 4476 23559
rect 4632 23186 4660 26200
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4908 23730 4936 24142
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4816 22545 4844 22578
rect 4802 22536 4858 22545
rect 4802 22471 4858 22480
rect 4526 21992 4582 22001
rect 4526 21927 4582 21936
rect 4540 19553 4568 21927
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4526 19544 4582 19553
rect 4526 19479 4582 19488
rect 4632 18970 4660 21490
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4724 21146 4752 21286
rect 4802 21176 4858 21185
rect 4712 21140 4764 21146
rect 4802 21111 4858 21120
rect 4712 21082 4764 21088
rect 4816 19854 4844 21111
rect 4908 21010 4936 23258
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4894 19952 4950 19961
rect 4894 19887 4950 19896
rect 4908 19854 4936 19887
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4816 19378 4844 19790
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4908 18086 4936 19790
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4172 16726 4200 17478
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4080 11014 4108 14010
rect 4172 13870 4200 15914
rect 4264 14618 4292 17206
rect 5000 17202 5028 22986
rect 5092 21486 5120 26302
rect 5354 26200 5410 27000
rect 5446 26888 5502 26897
rect 5446 26823 5502 26832
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4448 15366 4476 15438
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4356 14793 4384 14894
rect 4342 14784 4398 14793
rect 4342 14719 4398 14728
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4448 11354 4476 15302
rect 4540 15162 4568 17070
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4632 14618 4660 17138
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4724 15706 4752 16526
rect 4894 15736 4950 15745
rect 4712 15700 4764 15706
rect 4894 15671 4950 15680
rect 4712 15642 4764 15648
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4816 14074 4844 14554
rect 4908 14414 4936 15671
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 5092 12434 5120 19110
rect 5184 18834 5212 23462
rect 5276 21554 5304 25230
rect 5368 23798 5396 26200
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5460 23118 5488 26823
rect 5632 26376 5684 26382
rect 5632 26318 5684 26324
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5356 22704 5408 22710
rect 5356 22646 5408 22652
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5262 18728 5318 18737
rect 5262 18663 5318 18672
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 18329 5212 18566
rect 5170 18320 5226 18329
rect 5170 18255 5226 18264
rect 5276 14278 5304 18663
rect 5368 16658 5396 22646
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5460 20398 5488 21830
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5446 19136 5502 19145
rect 5446 19071 5502 19080
rect 5460 18970 5488 19071
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5460 16522 5488 17546
rect 5448 16516 5500 16522
rect 5448 16458 5500 16464
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5368 12753 5396 16050
rect 5446 15872 5502 15881
rect 5446 15807 5502 15816
rect 5460 14278 5488 15807
rect 5552 15502 5580 19654
rect 5644 18358 5672 26318
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26200 6514 27000
rect 6826 26200 6882 27000
rect 7194 26330 7250 27000
rect 7194 26302 7512 26330
rect 7194 26200 7250 26302
rect 5736 22710 5764 26200
rect 5814 25528 5870 25537
rect 5814 25463 5870 25472
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5722 21856 5778 21865
rect 5722 21791 5778 21800
rect 5736 19786 5764 21791
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5828 19718 5856 25463
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5920 19530 5948 22646
rect 6104 22098 6132 26200
rect 6276 26172 6328 26178
rect 6276 26114 6328 26120
rect 6184 25220 6236 25226
rect 6184 25162 6236 25168
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6090 21992 6146 22001
rect 6090 21927 6146 21936
rect 6104 21350 6132 21927
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6104 20466 6132 21286
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6012 19990 6040 20402
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 5736 19502 5948 19530
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5644 16697 5672 17478
rect 5630 16688 5686 16697
rect 5630 16623 5686 16632
rect 5736 16454 5764 19502
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15094 5580 15438
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5632 14544 5684 14550
rect 5538 14512 5594 14521
rect 5632 14486 5684 14492
rect 5538 14447 5594 14456
rect 5552 14414 5580 14447
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5552 14074 5580 14350
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5460 13297 5488 13398
rect 5446 13288 5502 13297
rect 5446 13223 5502 13232
rect 5354 12744 5410 12753
rect 5354 12679 5410 12688
rect 5000 12406 5120 12434
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 1766 9616 1822 9625
rect 1766 9551 1822 9560
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 5000 7993 5028 12406
rect 5644 11121 5672 14486
rect 5828 11257 5856 19314
rect 5908 17808 5960 17814
rect 5908 17750 5960 17756
rect 5920 17105 5948 17750
rect 5906 17096 5962 17105
rect 5906 17031 5962 17040
rect 6012 16998 6040 19722
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5920 13530 5948 16594
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 6012 15502 6040 16458
rect 6104 15706 6132 18702
rect 6196 18358 6224 25162
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 6196 17762 6224 18294
rect 6288 18086 6316 26114
rect 6472 24274 6500 26200
rect 6552 25424 6604 25430
rect 6552 25366 6604 25372
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6564 23866 6592 25366
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6564 22094 6592 23802
rect 6734 22672 6790 22681
rect 6644 22636 6696 22642
rect 6734 22607 6790 22616
rect 6644 22578 6696 22584
rect 6380 22066 6592 22094
rect 6380 19922 6408 22066
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21418 6500 21830
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6656 20806 6684 22578
rect 6748 22574 6776 22607
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 21622 6776 22374
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6840 21010 6868 26200
rect 7380 25560 7432 25566
rect 7380 25502 7432 25508
rect 7288 25152 7340 25158
rect 7010 25120 7066 25129
rect 7288 25094 7340 25100
rect 7010 25055 7066 25064
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6932 21078 6960 22578
rect 7024 21865 7052 25055
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7010 21856 7066 21865
rect 7010 21791 7066 21800
rect 7116 21706 7144 24142
rect 7024 21678 7144 21706
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 7024 20924 7052 21678
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6932 20896 7052 20924
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6644 20800 6696 20806
rect 6932 20754 6960 20896
rect 6644 20742 6696 20748
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6472 18714 6500 20742
rect 6840 20726 6960 20754
rect 6840 20584 6868 20726
rect 6748 20556 6868 20584
rect 6920 20596 6972 20602
rect 6748 20346 6776 20556
rect 6920 20538 6972 20544
rect 6826 20496 6882 20505
rect 6932 20466 6960 20538
rect 6826 20431 6828 20440
rect 6880 20431 6882 20440
rect 6920 20460 6972 20466
rect 6828 20402 6880 20408
rect 6920 20402 6972 20408
rect 6748 20318 6960 20346
rect 6550 19816 6606 19825
rect 6550 19751 6552 19760
rect 6604 19751 6606 19760
rect 6552 19722 6604 19728
rect 6564 18834 6592 19722
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6840 18766 6868 19110
rect 6828 18760 6880 18766
rect 6472 18686 6592 18714
rect 6828 18702 6880 18708
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6196 17734 6316 17762
rect 6288 17678 6316 17734
rect 6184 17672 6236 17678
rect 6182 17640 6184 17649
rect 6276 17672 6328 17678
rect 6236 17640 6238 17649
rect 6276 17614 6328 17620
rect 6182 17575 6238 17584
rect 6380 16402 6408 18566
rect 6460 16720 6512 16726
rect 6460 16662 6512 16668
rect 6288 16374 6408 16402
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6288 14498 6316 16374
rect 6366 16280 6422 16289
rect 6366 16215 6422 16224
rect 6380 16114 6408 16215
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6472 15706 6500 16662
rect 6564 16658 6592 18686
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6656 16182 6684 18022
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6564 15042 6592 16050
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6656 15502 6684 15914
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6748 15178 6776 17682
rect 6840 15706 6868 18566
rect 6932 17882 6960 20318
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7024 17338 7052 19722
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6920 17264 6972 17270
rect 6918 17232 6920 17241
rect 6972 17232 6974 17241
rect 6918 17167 6974 17176
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6748 15150 6868 15178
rect 6472 15014 6592 15042
rect 6734 15056 6790 15065
rect 6472 14618 6500 15014
rect 6734 14991 6790 15000
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6564 14618 6592 14894
rect 6748 14890 6776 14991
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6092 14476 6144 14482
rect 6288 14470 6408 14498
rect 6092 14418 6144 14424
rect 6104 14074 6132 14418
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6104 13938 6132 14010
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5814 11248 5870 11257
rect 5814 11183 5870 11192
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 4986 7984 5042 7993
rect 4986 7919 5042 7928
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 6288 6866 6316 14350
rect 6380 13569 6408 14470
rect 6840 14074 6868 15150
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6366 13560 6422 13569
rect 6366 13495 6422 13504
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12889 6592 13126
rect 6550 12880 6606 12889
rect 6550 12815 6606 12824
rect 6932 12374 6960 16730
rect 7116 15910 7144 21490
rect 7208 17338 7236 24890
rect 7300 22642 7328 25094
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7392 22030 7420 25502
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7484 21486 7512 26302
rect 7562 26200 7618 27000
rect 7930 26330 7986 27000
rect 7668 26302 7986 26330
rect 7576 23662 7604 26200
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7668 23186 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26200 8722 27000
rect 9034 26330 9090 27000
rect 8772 26302 9090 26330
rect 7930 25664 7986 25673
rect 7930 25599 7986 25608
rect 7944 25265 7972 25599
rect 7930 25256 7986 25265
rect 7930 25191 7986 25200
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7656 23180 7708 23186
rect 7656 23122 7708 23128
rect 7760 23066 7788 24754
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7944 23526 7972 23666
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7668 23038 7788 23066
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7288 20936 7340 20942
rect 7564 20936 7616 20942
rect 7288 20878 7340 20884
rect 7470 20904 7526 20913
rect 7300 19786 7328 20878
rect 7564 20878 7616 20884
rect 7470 20839 7526 20848
rect 7484 20602 7512 20839
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7576 20534 7604 20878
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 7470 20088 7526 20097
rect 7668 20058 7696 23038
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 20466 7788 22442
rect 7852 21622 7880 22918
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22098 8340 26200
rect 8574 24984 8630 24993
rect 8574 24919 8630 24928
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23322 8432 24006
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8300 22092 8352 22098
rect 8588 22080 8616 24919
rect 8680 24138 8708 26200
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9692 26302 9826 26330
rect 9218 25256 9274 25265
rect 9218 25191 9274 25200
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23497 9168 24006
rect 9126 23488 9182 23497
rect 9126 23423 9182 23432
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8588 22052 8708 22080
rect 8300 22034 8352 22040
rect 8576 21956 8628 21962
rect 8680 21944 8708 22052
rect 8680 21916 8800 21944
rect 8576 21898 8628 21904
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 21616 7892 21622
rect 7840 21558 7892 21564
rect 8298 21584 8354 21593
rect 8298 21519 8354 21528
rect 8312 20874 8340 21519
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8404 20641 8432 20878
rect 8390 20632 8446 20641
rect 8390 20567 8446 20576
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 7838 20360 7894 20369
rect 7838 20295 7894 20304
rect 7746 20224 7802 20233
rect 7746 20159 7802 20168
rect 7470 20023 7526 20032
rect 7656 20052 7708 20058
rect 7288 19780 7340 19786
rect 7288 19722 7340 19728
rect 7286 19544 7342 19553
rect 7286 19479 7342 19488
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7300 17218 7328 19479
rect 7484 19446 7512 20023
rect 7656 19994 7708 20000
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7208 17190 7328 17218
rect 7208 16114 7236 17190
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15609 7236 15846
rect 7194 15600 7250 15609
rect 7194 15535 7250 15544
rect 7208 15502 7236 15535
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 7024 12209 7052 13942
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7116 13530 7144 13874
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7208 12850 7236 15302
rect 7300 14770 7328 17002
rect 7392 16674 7420 18226
rect 7470 18048 7526 18057
rect 7470 17983 7526 17992
rect 7484 17678 7512 17983
rect 7576 17785 7604 18634
rect 7760 18630 7788 20159
rect 7852 19378 7880 20295
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19854 7972 20198
rect 8024 19984 8076 19990
rect 8128 19961 8156 20402
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8312 19961 8340 20266
rect 8024 19926 8076 19932
rect 8114 19952 8170 19961
rect 8036 19854 8064 19926
rect 8114 19887 8170 19896
rect 8298 19952 8354 19961
rect 8298 19887 8354 19896
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7654 18456 7710 18465
rect 7654 18391 7710 18400
rect 7668 18222 7696 18391
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 18086 7696 18158
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7562 17776 7618 17785
rect 7562 17711 7618 17720
rect 7852 17678 7880 19110
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8404 18465 8432 19654
rect 8390 18456 8446 18465
rect 8390 18391 8446 18400
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8206 18184 8262 18193
rect 8206 18119 8208 18128
rect 8260 18119 8262 18128
rect 8208 18090 8260 18096
rect 8312 18057 8340 18294
rect 8496 18204 8524 21286
rect 8588 21010 8616 21898
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8588 20534 8616 20810
rect 8666 20768 8722 20777
rect 8666 20703 8722 20712
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19446 8616 19654
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8680 19242 8708 20703
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8772 18970 8800 21916
rect 8956 21894 8984 22918
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9048 22030 9076 22510
rect 9126 22264 9182 22273
rect 9126 22199 9182 22208
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 9048 21554 9076 21966
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 21010 9076 21490
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 9036 21004 9088 21010
rect 9036 20946 9088 20952
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8588 18358 8616 18566
rect 8680 18426 8708 18566
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8496 18176 8616 18204
rect 8298 18048 8354 18057
rect 8298 17983 8354 17992
rect 8298 17912 8354 17921
rect 8298 17847 8354 17856
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7484 16794 7512 17614
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7392 16646 7512 16674
rect 7300 14742 7420 14770
rect 7286 14376 7342 14385
rect 7286 14311 7342 14320
rect 7300 14278 7328 14311
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7010 12200 7066 12209
rect 7010 12135 7066 12144
rect 7392 11801 7420 14742
rect 7484 12306 7512 16646
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7576 16114 7604 16390
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 13870 7604 14826
rect 7668 14006 7696 17614
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 15094 7880 17478
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17134 8340 17847
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8496 17513 8524 17546
rect 8482 17504 8538 17513
rect 8482 17439 8538 17448
rect 8300 17128 8352 17134
rect 8352 17088 8524 17116
rect 8300 17070 8352 17076
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8206 15600 8262 15609
rect 8206 15535 8208 15544
rect 8260 15535 8262 15544
rect 8208 15506 8260 15512
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8390 15192 8446 15201
rect 8390 15127 8446 15136
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14822 8340 14894
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7760 14278 7788 14486
rect 7852 14414 7880 14486
rect 7840 14408 7892 14414
rect 7840 14350 7892 14356
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7760 13802 7788 14214
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7932 14000 7984 14006
rect 7838 13968 7894 13977
rect 7932 13942 7984 13948
rect 7838 13903 7840 13912
rect 7892 13903 7894 13912
rect 7840 13874 7892 13880
rect 7944 13841 7972 13942
rect 7930 13832 7986 13841
rect 7748 13796 7800 13802
rect 7930 13767 7986 13776
rect 7748 13738 7800 13744
rect 8312 13462 8340 14758
rect 8404 14550 8432 15127
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8496 14074 8524 17088
rect 8588 15162 8616 18176
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8680 17377 8708 17750
rect 8666 17368 8722 17377
rect 8666 17303 8722 17312
rect 8666 16552 8722 16561
rect 8666 16487 8722 16496
rect 8680 16454 8708 16487
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8680 15706 8708 15846
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8772 15502 8800 18770
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8772 14929 8800 14962
rect 8758 14920 8814 14929
rect 8758 14855 8814 14864
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8312 12481 8340 12854
rect 8298 12472 8354 12481
rect 8298 12407 8354 12416
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7378 11792 7434 11801
rect 7378 11727 7434 11736
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8588 9110 8616 14758
rect 8864 14414 8892 20946
rect 9048 20466 9076 20946
rect 9140 20942 9168 22199
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8956 19689 8984 19994
rect 8942 19680 8998 19689
rect 8942 19615 8998 19624
rect 9048 19378 9076 20402
rect 9036 19372 9088 19378
rect 9088 19320 9168 19334
rect 9036 19314 9168 19320
rect 9048 19306 9168 19314
rect 9140 18578 9168 19306
rect 8956 18550 9168 18578
rect 8956 18290 8984 18550
rect 9034 18456 9090 18465
rect 9034 18391 9090 18400
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17678 8984 18226
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 17202 8984 17614
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9048 16810 9076 18391
rect 9232 17898 9260 25191
rect 9416 23186 9444 26200
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9324 21078 9352 21830
rect 9416 21350 9444 21830
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9402 21040 9458 21049
rect 9324 20233 9352 21014
rect 9402 20975 9458 20984
rect 9416 20942 9444 20975
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9402 20632 9458 20641
rect 9402 20567 9458 20576
rect 9416 20398 9444 20567
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9310 20224 9366 20233
rect 9310 20159 9366 20168
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9324 19689 9352 19926
rect 9310 19680 9366 19689
rect 9310 19615 9366 19624
rect 9404 19304 9456 19310
rect 9402 19272 9404 19281
rect 9456 19272 9458 19281
rect 9402 19207 9458 19216
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 8956 16782 9076 16810
rect 9140 17870 9260 17898
rect 9140 16794 9168 17870
rect 9128 16788 9180 16794
rect 8956 16454 8984 16782
rect 9128 16730 9180 16736
rect 8944 16448 8996 16454
rect 9140 16402 9168 16730
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 8944 16390 8996 16396
rect 9048 16374 9168 16402
rect 9048 16114 9076 16374
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9140 16017 9168 16186
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 9140 13530 9168 15302
rect 9232 15162 9260 16662
rect 9324 16114 9352 18362
rect 9508 17218 9536 24822
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26330 11298 27000
rect 11072 26302 11298 26330
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9692 23905 9720 24074
rect 9678 23896 9734 23905
rect 9678 23831 9734 23840
rect 9770 23760 9826 23769
rect 9770 23695 9772 23704
rect 9824 23695 9826 23704
rect 9772 23666 9824 23672
rect 9876 23633 9904 24142
rect 10152 23798 10180 26200
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10048 23724 10100 23730
rect 10048 23666 10100 23672
rect 9862 23624 9918 23633
rect 9862 23559 9918 23568
rect 10060 23497 10088 23666
rect 10230 23624 10286 23633
rect 10230 23559 10286 23568
rect 10046 23488 10102 23497
rect 10046 23423 10102 23432
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9864 23044 9916 23050
rect 9864 22986 9916 22992
rect 9772 22568 9824 22574
rect 9600 22516 9772 22522
rect 9600 22510 9824 22516
rect 9600 22494 9812 22510
rect 9600 22234 9628 22494
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9600 20233 9628 20470
rect 9586 20224 9642 20233
rect 9586 20159 9642 20168
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9600 19786 9628 19858
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9692 19514 9720 22170
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9784 19854 9812 19994
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9784 18970 9812 19654
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 17626 9628 18566
rect 9600 17598 9720 17626
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9416 17190 9536 17218
rect 9416 16658 9444 17190
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 14074 9260 14962
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 12209 9260 14010
rect 9416 13258 9444 16390
rect 9508 16250 9536 17070
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9600 16114 9628 17478
rect 9692 16946 9720 17598
rect 9876 17252 9904 22986
rect 9968 18952 9996 23054
rect 10152 22166 10180 23054
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10244 21078 10272 23559
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 10336 19938 10364 22918
rect 10428 22094 10456 23462
rect 10520 23186 10548 26200
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10428 22066 10548 22094
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10060 19910 10364 19938
rect 10428 19922 10456 20266
rect 10416 19916 10468 19922
rect 10060 19174 10088 19910
rect 10416 19858 10468 19864
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10336 19122 10364 19790
rect 10416 19168 10468 19174
rect 10336 19116 10416 19122
rect 10336 19110 10468 19116
rect 10336 19094 10456 19110
rect 10232 18964 10284 18970
rect 9968 18924 10180 18952
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 18216 10008 18222
rect 10060 18204 10088 18770
rect 10008 18176 10088 18204
rect 9956 18158 10008 18164
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 17610 9996 18022
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9876 17224 9996 17252
rect 9692 16918 9812 16946
rect 9678 16824 9734 16833
rect 9678 16759 9680 16768
rect 9732 16759 9734 16768
rect 9680 16730 9732 16736
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9692 15502 9720 16730
rect 9784 16454 9812 16918
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9784 15366 9812 15399
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9968 15162 9996 17224
rect 10060 17134 10088 18176
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 13977 9720 14282
rect 9876 14278 9904 14962
rect 10060 14498 10088 16730
rect 10152 14958 10180 18924
rect 10232 18906 10284 18912
rect 10244 15434 10272 18906
rect 10336 18766 10364 19094
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10520 18306 10548 22066
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10612 21418 10640 22034
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10612 20058 10640 20742
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10336 18278 10548 18306
rect 10336 17241 10364 18278
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10322 17232 10378 17241
rect 10322 17167 10378 17176
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 16182 10364 16390
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 9968 14482 10088 14498
rect 9956 14476 10088 14482
rect 10008 14470 10088 14476
rect 9956 14418 10008 14424
rect 10336 14414 10364 15030
rect 10428 14550 10456 18158
rect 10612 17320 10640 19654
rect 10704 19310 10732 25638
rect 10888 23798 10916 26200
rect 11072 24324 11100 26302
rect 11242 26200 11298 26302
rect 11610 26200 11666 27000
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26200 12770 27000
rect 13082 26330 13138 27000
rect 12820 26302 13138 26330
rect 11244 24676 11296 24682
rect 11244 24618 11296 24624
rect 10980 24296 11100 24324
rect 10980 24206 11008 24296
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10980 23526 11008 24006
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 11072 23338 11100 24006
rect 10980 23310 11100 23338
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10796 21944 10824 22578
rect 10980 22098 11008 23310
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11164 22710 11192 23190
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 11164 22574 11192 22646
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11150 22400 11206 22409
rect 11150 22335 11206 22344
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10876 21956 10928 21962
rect 10796 21916 10876 21944
rect 10796 21622 10824 21916
rect 10876 21898 10928 21904
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20466 11100 20878
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10784 19984 10836 19990
rect 10836 19944 10916 19972
rect 10784 19926 10836 19932
rect 10888 19718 10916 19944
rect 11072 19922 11100 20198
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10888 19174 10916 19382
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10876 19168 10928 19174
rect 10980 19145 11008 19178
rect 10876 19110 10928 19116
rect 10966 19136 11022 19145
rect 10888 18426 10916 19110
rect 10966 19071 11022 19080
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10888 18290 10916 18362
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10784 17604 10836 17610
rect 10888 17592 10916 18226
rect 10836 17564 10916 17592
rect 10784 17546 10836 17552
rect 10520 17292 10640 17320
rect 10520 15638 10548 17292
rect 10784 17264 10836 17270
rect 10784 17206 10836 17212
rect 10796 16726 10824 17206
rect 10888 17202 10916 17564
rect 11072 17241 11100 18634
rect 11058 17232 11114 17241
rect 10876 17196 10928 17202
rect 11058 17167 11114 17176
rect 10876 17138 10928 17144
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15026 10548 15302
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 10138 14240 10194 14249
rect 9678 13968 9734 13977
rect 9678 13903 9734 13912
rect 9678 13832 9734 13841
rect 9678 13767 9734 13776
rect 9692 13734 9720 13767
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9586 13560 9642 13569
rect 9586 13495 9642 13504
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9600 12889 9628 13495
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 13161 9720 13330
rect 9678 13152 9734 13161
rect 9678 13087 9734 13096
rect 9586 12880 9642 12889
rect 9586 12815 9642 12824
rect 9218 12200 9274 12209
rect 9218 12135 9274 12144
rect 9876 12102 9904 14214
rect 10138 14175 10194 14184
rect 10152 14006 10180 14175
rect 10232 14068 10284 14074
rect 10336 14056 10364 14350
rect 10284 14028 10364 14056
rect 10232 14010 10284 14016
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 10060 9042 10088 13126
rect 10612 12986 10640 16594
rect 10888 16538 10916 17138
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16658 11100 16934
rect 11164 16794 11192 22335
rect 11256 22080 11284 24618
rect 11520 24336 11572 24342
rect 11520 24278 11572 24284
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11348 23662 11376 23802
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11336 22092 11388 22098
rect 11256 22052 11336 22080
rect 11256 21690 11284 22052
rect 11336 22034 11388 22040
rect 11532 21876 11560 24278
rect 11624 23322 11652 26200
rect 11992 23662 12020 26200
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12070 23352 12126 23361
rect 11612 23316 11664 23322
rect 12070 23287 12126 23296
rect 11612 23258 11664 23264
rect 11980 23044 12032 23050
rect 11980 22986 12032 22992
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11716 22234 11744 22374
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11796 21888 11848 21894
rect 11532 21848 11744 21876
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11532 20874 11560 21490
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11532 20534 11560 20810
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10704 16510 10916 16538
rect 10704 16046 10732 16510
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16250 10916 16390
rect 11150 16280 11206 16289
rect 10876 16244 10928 16250
rect 11256 16250 11284 20402
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18766 11376 19110
rect 11440 19009 11468 20198
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11518 19680 11574 19689
rect 11518 19615 11574 19624
rect 11426 19000 11482 19009
rect 11426 18935 11482 18944
rect 11336 18760 11388 18766
rect 11440 18737 11468 18935
rect 11336 18702 11388 18708
rect 11426 18728 11482 18737
rect 11348 18426 11376 18702
rect 11426 18663 11482 18672
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11150 16215 11206 16224
rect 11244 16244 11296 16250
rect 10876 16186 10928 16192
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10888 15026 10916 15370
rect 11072 15162 11100 15982
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10888 14346 10916 14962
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14482 11008 14758
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 11164 14362 11192 16215
rect 11244 16186 11296 16192
rect 11242 15328 11298 15337
rect 11242 15263 11298 15272
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 11072 14334 11192 14362
rect 10888 13394 10916 14282
rect 11072 13938 11100 14334
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13938 11192 14214
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 13190 10916 13330
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 11072 12714 11100 13670
rect 11164 12986 11192 13874
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11256 12918 11284 15263
rect 11348 13870 11376 18022
rect 11532 17814 11560 19615
rect 11624 19514 11652 19790
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11716 19310 11744 21848
rect 11796 21830 11848 21836
rect 11808 21010 11836 21830
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11624 18970 11652 19246
rect 11612 18964 11664 18970
rect 11612 18906 11664 18912
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11612 17808 11664 17814
rect 11612 17750 11664 17756
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17270 11468 17478
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11532 17066 11560 17750
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11518 16824 11574 16833
rect 11518 16759 11574 16768
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 15366 11468 16594
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11532 13410 11560 16759
rect 11624 15094 11652 17750
rect 11716 17746 11744 18566
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17202 11744 17682
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16046 11744 16526
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11716 15026 11744 15982
rect 11808 15745 11836 20198
rect 11900 18834 11928 22578
rect 11992 22438 12020 22986
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11992 20330 12020 21830
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 12084 20097 12112 23287
rect 12176 22273 12204 24618
rect 12360 24342 12388 26200
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12348 24336 12400 24342
rect 12532 24336 12584 24342
rect 12348 24278 12400 24284
rect 12452 24296 12532 24324
rect 12256 23520 12308 23526
rect 12452 23474 12480 24296
rect 12532 24278 12584 24284
rect 12256 23462 12308 23468
rect 12268 23118 12296 23462
rect 12360 23446 12480 23474
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12360 22982 12388 23446
rect 12636 23338 12664 24346
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12544 23310 12664 23338
rect 12452 23225 12480 23258
rect 12438 23216 12494 23225
rect 12438 23151 12494 23160
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12162 22264 12218 22273
rect 12162 22199 12218 22208
rect 12268 21894 12296 22510
rect 12360 21962 12388 22578
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12268 21486 12296 21626
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12256 21480 12308 21486
rect 12308 21440 12388 21468
rect 12256 21422 12308 21428
rect 12070 20088 12126 20097
rect 12070 20023 12126 20032
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 12084 18222 12112 19314
rect 12176 18290 12204 21422
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 20398 12296 21286
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12360 18306 12388 21440
rect 12452 19938 12480 22578
rect 12544 22094 12572 23310
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12636 23050 12664 23190
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12728 22409 12756 26200
rect 12820 22953 12848 26302
rect 13082 26200 13138 26302
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26200 14242 27000
rect 14554 26200 14610 27000
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15658 26200 15714 27000
rect 16026 26330 16082 27000
rect 15856 26302 16082 26330
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13266 23216 13322 23225
rect 13464 23202 13492 26200
rect 13544 25016 13596 25022
rect 13544 24958 13596 24964
rect 13322 23174 13492 23202
rect 13266 23151 13322 23160
rect 12806 22944 12862 22953
rect 12806 22879 12862 22888
rect 12714 22400 12770 22409
rect 12714 22335 12770 22344
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12544 22066 12664 22094
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12544 21690 12572 21830
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12544 21554 12572 21626
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12636 20534 12664 22066
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12624 20392 12676 20398
rect 12530 20360 12586 20369
rect 12624 20334 12676 20340
rect 12530 20295 12586 20304
rect 12544 20097 12572 20295
rect 12530 20088 12586 20097
rect 12530 20023 12586 20032
rect 12452 19910 12572 19938
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12268 18278 12388 18306
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12268 17490 12296 18278
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 11900 17462 12296 17490
rect 11794 15736 11850 15745
rect 11794 15671 11850 15680
rect 11900 15314 11928 17462
rect 12360 16454 12388 18158
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11808 15286 11928 15314
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11808 14634 11836 15286
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11624 14606 11836 14634
rect 11624 13734 11652 14606
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11808 13530 11836 13738
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11532 13382 11836 13410
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11624 12918 11652 13194
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 10130 11008 12582
rect 11624 12442 11652 12854
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12714 11744 12786
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11716 12442 11744 12650
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11704 12436 11756 12442
rect 11808 12434 11836 13382
rect 11900 12850 11928 15098
rect 11992 13938 12020 15982
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12084 14618 12112 15506
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 14006 12112 14350
rect 12268 14074 12296 15030
rect 12360 14414 12388 15438
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12452 13734 12480 18158
rect 12544 17542 12572 19910
rect 12636 17882 12664 20334
rect 12728 18222 12756 22170
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21486 13124 21966
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12820 20602 12848 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12912 20312 12940 20878
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 12820 20284 12940 20312
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12636 17338 12664 17818
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12728 17218 12756 18022
rect 12636 17190 12756 17218
rect 12530 16688 12586 16697
rect 12530 16623 12586 16632
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12544 13546 12572 16623
rect 12636 15706 12664 17190
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16522 12756 17070
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12728 16182 12756 16458
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12728 15502 12756 16118
rect 12716 15496 12768 15502
rect 12636 15456 12716 15484
rect 12636 15094 12664 15456
rect 12716 15438 12768 15444
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12636 13938 12664 14486
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12452 13518 12572 13546
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12084 12986 12112 13194
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11808 12406 12296 12434
rect 11704 12378 11756 12384
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11898 11928 12174
rect 12268 11898 12296 12406
rect 12360 12238 12388 12786
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10742 11744 10950
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 11900 9178 11928 11834
rect 12452 11286 12480 13518
rect 12728 12782 12756 15302
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12544 11218 12572 12038
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12820 9926 12848 20284
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19922 13400 20538
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13464 19786 13492 20402
rect 13556 20369 13584 24958
rect 13728 24268 13780 24274
rect 13728 24210 13780 24216
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13648 23254 13676 23734
rect 13636 23248 13688 23254
rect 13636 23190 13688 23196
rect 13740 22094 13768 24210
rect 13832 23848 13860 26200
rect 14094 24848 14150 24857
rect 14094 24783 14150 24792
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13832 23820 13952 23848
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13832 23526 13860 23666
rect 13820 23520 13872 23526
rect 13818 23488 13820 23497
rect 13872 23488 13874 23497
rect 13818 23423 13874 23432
rect 13924 23186 13952 23820
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22710 13860 23054
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13648 22066 13768 22094
rect 14016 22094 14044 24006
rect 14108 23866 14136 24783
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14200 22234 14228 26200
rect 14372 25084 14424 25090
rect 14372 25026 14424 25032
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14292 22098 14320 23054
rect 14016 22066 14228 22094
rect 13648 21865 13676 22066
rect 13728 21888 13780 21894
rect 13634 21856 13690 21865
rect 13728 21830 13780 21836
rect 13634 21791 13690 21800
rect 13636 21344 13688 21350
rect 13634 21312 13636 21321
rect 13688 21312 13690 21321
rect 13634 21247 13690 21256
rect 13542 20360 13598 20369
rect 13542 20295 13598 20304
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19530 13216 19654
rect 13188 19502 13308 19530
rect 13174 19408 13230 19417
rect 13174 19343 13230 19352
rect 13188 19174 13216 19343
rect 13280 19334 13308 19502
rect 13464 19446 13492 19722
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13556 19334 13584 19722
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13280 19306 13584 19334
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13542 19136 13598 19145
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18766 13400 19110
rect 13542 19071 13598 19080
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18222 12940 18566
rect 13280 18358 13308 18634
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17134 13032 17546
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13372 17082 13400 18158
rect 13464 17882 13492 18634
rect 13556 18426 13584 19071
rect 13648 18970 13676 19654
rect 13740 19310 13768 21830
rect 14200 21690 14228 22066
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14108 20874 14136 21626
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14200 21146 14228 21354
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 14292 20618 14320 22034
rect 14384 21729 14412 25026
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14370 21720 14426 21729
rect 14370 21655 14426 21664
rect 14476 21622 14504 24346
rect 14568 23497 14596 26200
rect 14936 25945 14964 26200
rect 14922 25936 14978 25945
rect 14922 25871 14978 25880
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14648 23520 14700 23526
rect 14554 23488 14610 23497
rect 14648 23462 14700 23468
rect 14554 23423 14610 23432
rect 14660 23032 14688 23462
rect 14568 23004 14688 23032
rect 14568 22710 14596 23004
rect 14646 22944 14702 22953
rect 14646 22879 14702 22888
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14568 21962 14596 22646
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14568 21554 14596 21898
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14200 20602 14320 20618
rect 14188 20596 14320 20602
rect 14240 20590 14320 20596
rect 14188 20538 14240 20544
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13832 19514 13860 20470
rect 13924 19910 14320 19938
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13636 18964 13688 18970
rect 13688 18924 13768 18952
rect 13636 18906 13688 18912
rect 13740 18698 13768 18924
rect 13832 18834 13860 19450
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13636 18692 13688 18698
rect 13636 18634 13688 18640
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13556 17270 13584 18226
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13648 17202 13676 18634
rect 13740 17338 13768 18634
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13832 17134 13860 18362
rect 13820 17128 13872 17134
rect 13372 17054 13492 17082
rect 13820 17070 13872 17076
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13372 16833 13400 16934
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 12238 13400 15506
rect 13464 12850 13492 17054
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13556 15910 13584 17002
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13726 15872 13782 15881
rect 13556 14414 13584 15846
rect 13726 15807 13782 15816
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 15162 13676 15302
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13648 14006 13676 14826
rect 13740 14822 13768 15807
rect 13924 15502 13952 19910
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14016 19378 14044 19790
rect 14200 19689 14228 19790
rect 14292 19718 14320 19910
rect 14280 19712 14332 19718
rect 14186 19680 14242 19689
rect 14280 19654 14332 19660
rect 14186 19615 14242 19624
rect 14384 19530 14412 21286
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14200 19502 14412 19530
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 14016 18426 14044 19178
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 16658 14044 17478
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14108 17134 14136 17274
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16794 14136 16934
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13832 14550 13860 15098
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13832 14278 13860 14486
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13634 13832 13690 13841
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13556 12617 13584 13806
rect 13634 13767 13690 13776
rect 13542 12608 13598 12617
rect 13542 12543 13598 12552
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11830 13124 12038
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 13556 11694 13584 12543
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13648 10810 13676 13767
rect 13832 13394 13860 14214
rect 14016 13530 14044 16390
rect 14200 15994 14228 19502
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14370 19408 14426 19417
rect 14292 18970 14320 19382
rect 14370 19343 14426 19352
rect 14384 19009 14412 19343
rect 14370 19000 14426 19009
rect 14280 18964 14332 18970
rect 14370 18935 14426 18944
rect 14280 18906 14332 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14292 18426 14320 18770
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14278 17776 14334 17785
rect 14278 17711 14280 17720
rect 14332 17711 14334 17720
rect 14280 17682 14332 17688
rect 14108 15966 14228 15994
rect 14108 14482 14136 15966
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15026 14228 15846
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14200 14074 14228 14962
rect 14292 14482 14320 15506
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14292 14006 14320 14418
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 12442 13768 13194
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11694 13768 12174
rect 13832 11898 13860 12922
rect 14016 12238 14044 13466
rect 14292 13394 14320 13942
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12986 14320 13330
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13726 11520 13782 11529
rect 13726 11455 13782 11464
rect 13740 11150 13768 11455
rect 14384 11286 14412 18935
rect 14476 17814 14504 20878
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 20369 14596 20742
rect 14554 20360 14610 20369
rect 14554 20295 14610 20304
rect 14568 19514 14596 20295
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14568 17678 14596 18906
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14660 17320 14688 22879
rect 14752 19514 14780 24550
rect 15304 24410 15332 26200
rect 15382 24440 15438 24449
rect 15292 24404 15344 24410
rect 15382 24375 15438 24384
rect 15292 24346 15344 24352
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 14832 23044 14884 23050
rect 14832 22986 14884 22992
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14752 17542 14780 19110
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14568 17292 14688 17320
rect 14568 16697 14596 17292
rect 14738 17232 14794 17241
rect 14648 17196 14700 17202
rect 14738 17167 14794 17176
rect 14648 17138 14700 17144
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14476 12170 14504 16458
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14568 15910 14596 15982
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14568 15162 14596 15370
rect 14660 15366 14688 17138
rect 14752 16969 14780 17167
rect 14738 16960 14794 16969
rect 14738 16895 14794 16904
rect 14752 16114 14780 16895
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14482 14596 14758
rect 14646 14648 14702 14657
rect 14646 14583 14702 14592
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14554 14376 14610 14385
rect 14554 14311 14610 14320
rect 14568 14278 14596 14311
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14568 14006 14596 14214
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14554 11384 14610 11393
rect 14554 11319 14610 11328
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 13728 11144 13780 11150
rect 14568 11121 14596 11319
rect 13728 11086 13780 11092
rect 14554 11112 14610 11121
rect 14554 11047 14610 11056
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 13832 8906 13860 10746
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 10266 14504 10542
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14660 10062 14688 14583
rect 14844 10266 14872 22986
rect 14936 22234 14964 24006
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 15028 22386 15056 23734
rect 15120 22506 15148 24006
rect 15212 23662 15240 24142
rect 15396 24041 15424 24375
rect 15382 24032 15438 24041
rect 15382 23967 15438 23976
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 15304 23186 15332 23666
rect 15384 23656 15436 23662
rect 15476 23656 15528 23662
rect 15384 23598 15436 23604
rect 15474 23624 15476 23633
rect 15528 23624 15530 23633
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15396 22778 15424 23598
rect 15474 23559 15530 23568
rect 15672 23497 15700 26200
rect 15752 23520 15804 23526
rect 15658 23488 15714 23497
rect 15752 23462 15804 23468
rect 15658 23423 15714 23432
rect 15764 23050 15792 23462
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15028 22358 15148 22386
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 20890 14964 21490
rect 15028 21078 15056 22170
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 14936 20862 15056 20890
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14936 19174 14964 20742
rect 15028 20330 15056 20862
rect 15120 20398 15148 22358
rect 15212 20641 15240 22442
rect 15752 22092 15804 22098
rect 15672 22052 15752 22080
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15476 21480 15528 21486
rect 15568 21480 15620 21486
rect 15476 21422 15528 21428
rect 15566 21448 15568 21457
rect 15620 21448 15622 21457
rect 15198 20632 15254 20641
rect 15198 20567 15254 20576
rect 15304 20398 15332 21422
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15292 20392 15344 20398
rect 15292 20334 15344 20340
rect 15016 20324 15068 20330
rect 15016 20266 15068 20272
rect 15396 19802 15424 21354
rect 15488 20874 15516 21422
rect 15566 21383 15622 21392
rect 15672 21026 15700 22052
rect 15752 22034 15804 22040
rect 15752 21616 15804 21622
rect 15752 21558 15804 21564
rect 15764 21418 15792 21558
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15672 20998 15792 21026
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 20058 15516 20198
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15028 19774 15424 19802
rect 15028 19242 15056 19774
rect 15396 19718 15424 19774
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15120 19334 15148 19654
rect 15120 19306 15332 19334
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15016 18760 15068 18766
rect 14936 18720 15016 18748
rect 14936 18426 14964 18720
rect 15016 18702 15068 18708
rect 15304 18578 15332 19306
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15396 18902 15424 19110
rect 15488 18902 15516 19654
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15212 18550 15332 18578
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 14936 17746 14964 18362
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15028 18057 15056 18090
rect 15108 18080 15160 18086
rect 15014 18048 15070 18057
rect 15212 18068 15240 18550
rect 15396 18426 15424 18838
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15160 18040 15240 18068
rect 15108 18022 15160 18028
rect 15014 17983 15070 17992
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14936 16658 14964 17682
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 15028 16522 15056 17478
rect 15212 17338 15240 17546
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 15434 15056 16458
rect 15304 16182 15332 18362
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15106 16008 15162 16017
rect 15106 15943 15162 15952
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15028 15094 15056 15370
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15028 14385 15056 15030
rect 15014 14376 15070 14385
rect 15014 14311 15016 14320
rect 15068 14311 15070 14320
rect 15016 14282 15068 14288
rect 15028 13258 15056 14282
rect 15120 14056 15148 15943
rect 15396 14890 15424 18226
rect 15488 18222 15516 18838
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17338 15516 18022
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15474 17232 15530 17241
rect 15474 17167 15530 17176
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15212 14385 15240 14758
rect 15198 14376 15254 14385
rect 15198 14311 15254 14320
rect 15120 14028 15240 14056
rect 15212 13920 15240 14028
rect 15292 13932 15344 13938
rect 15212 13892 15292 13920
rect 15292 13874 15344 13880
rect 15290 13832 15346 13841
rect 15290 13767 15346 13776
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12850 15056 13194
rect 15212 13190 15240 13466
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 11830 15056 12786
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15028 11200 15056 11766
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14936 11172 15056 11200
rect 14936 11014 14964 11172
rect 15014 11112 15070 11121
rect 15014 11047 15070 11056
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10810 14964 10950
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 9722 14688 9998
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 15028 9450 15056 11047
rect 15120 10248 15148 11630
rect 15304 11286 15332 13767
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 12918 15424 13670
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15488 12764 15516 17167
rect 15580 16561 15608 20742
rect 15672 16833 15700 20878
rect 15764 19990 15792 20998
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15764 18630 15792 19178
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15856 17490 15884 26302
rect 16026 26200 16082 26302
rect 16394 26200 16450 27000
rect 16762 26200 16818 27000
rect 17130 26200 17186 27000
rect 17498 26200 17554 27000
rect 17866 26330 17922 27000
rect 18234 26330 18290 27000
rect 17788 26302 17922 26330
rect 16408 24682 16436 26200
rect 16776 25401 16804 26200
rect 17144 25673 17172 26200
rect 17130 25664 17186 25673
rect 17130 25599 17186 25608
rect 16762 25392 16818 25401
rect 16762 25327 16818 25336
rect 16396 24676 16448 24682
rect 16396 24618 16448 24624
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15764 17462 15884 17490
rect 15658 16824 15714 16833
rect 15658 16759 15714 16768
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15566 16552 15622 16561
rect 15566 16487 15622 16496
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15580 13530 15608 15943
rect 15672 14113 15700 16662
rect 15658 14104 15714 14113
rect 15658 14039 15714 14048
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 12850 15608 13126
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15396 12736 15516 12764
rect 15396 11286 15424 12736
rect 15764 12714 15792 17462
rect 15842 17368 15898 17377
rect 15842 17303 15844 17312
rect 15896 17303 15898 17312
rect 15844 17274 15896 17280
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15474 12336 15530 12345
rect 15474 12271 15476 12280
rect 15528 12271 15530 12280
rect 15476 12242 15528 12248
rect 15474 12200 15530 12209
rect 15474 12135 15476 12144
rect 15528 12135 15530 12144
rect 15476 12106 15528 12112
rect 15488 11801 15516 12106
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15580 10538 15608 12582
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15200 10260 15252 10266
rect 15120 10220 15200 10248
rect 15200 10202 15252 10208
rect 15290 10160 15346 10169
rect 15290 10095 15346 10104
rect 15304 10062 15332 10095
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15304 9722 15332 9998
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15660 9648 15712 9654
rect 15658 9616 15660 9625
rect 15712 9616 15714 9625
rect 15658 9551 15714 9560
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15856 9178 15884 16050
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6840 2650 6868 8842
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 15948 4826 15976 22646
rect 16040 22166 16068 23666
rect 16210 23624 16266 23633
rect 16210 23559 16266 23568
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16040 20097 16068 21898
rect 16132 21010 16160 22578
rect 16224 21962 16252 23559
rect 16316 22710 16344 24006
rect 16500 23730 16528 24006
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16488 23248 16540 23254
rect 16486 23216 16488 23225
rect 16540 23216 16542 23225
rect 16486 23151 16542 23160
rect 16776 22982 16804 24142
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16684 22817 16712 22918
rect 16670 22808 16726 22817
rect 16670 22743 16726 22752
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 16776 22574 16804 22918
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16396 22432 16448 22438
rect 16396 22374 16448 22380
rect 16302 22128 16358 22137
rect 16302 22063 16358 22072
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16316 21554 16344 22063
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16408 21400 16436 22374
rect 16486 22128 16542 22137
rect 16868 22098 16896 24142
rect 17130 23896 17186 23905
rect 17130 23831 17186 23840
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 17052 23322 17080 23462
rect 17040 23316 17092 23322
rect 17040 23258 17092 23264
rect 16946 23216 17002 23225
rect 16946 23151 17002 23160
rect 16960 22953 16988 23151
rect 17144 23118 17172 23831
rect 17408 23724 17460 23730
rect 17408 23666 17460 23672
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17040 22976 17092 22982
rect 16946 22944 17002 22953
rect 17040 22918 17092 22924
rect 16946 22879 17002 22888
rect 16486 22063 16542 22072
rect 16856 22092 16908 22098
rect 16500 22030 16528 22063
rect 16856 22034 16908 22040
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16580 22024 16632 22030
rect 17052 21978 17080 22918
rect 17132 22704 17184 22710
rect 17130 22672 17132 22681
rect 17184 22672 17186 22681
rect 17130 22607 17186 22616
rect 17130 22400 17186 22409
rect 17130 22335 17186 22344
rect 16580 21966 16632 21972
rect 16224 21372 16436 21400
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16224 20874 16252 21372
rect 16592 21350 16620 21966
rect 16684 21950 17080 21978
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16486 21176 16542 21185
rect 16486 21111 16542 21120
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16026 20088 16082 20097
rect 16026 20023 16082 20032
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19310 16068 19790
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 16794 16068 19246
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 14618 16068 15982
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16040 13870 16068 13942
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16040 11150 16068 13466
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16132 6662 16160 20402
rect 16224 19174 16252 20810
rect 16500 20777 16528 21111
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 16486 20768 16542 20777
rect 16486 20703 16542 20712
rect 16302 20632 16358 20641
rect 16302 20567 16358 20576
rect 16488 20596 16540 20602
rect 16316 20534 16344 20567
rect 16488 20538 16540 20544
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19718 16344 19790
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16408 19446 16436 20266
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16408 19242 16436 19382
rect 16500 19378 16528 20538
rect 16592 20369 16620 20946
rect 16578 20360 16634 20369
rect 16578 20295 16634 20304
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16212 18692 16264 18698
rect 16408 18680 16436 19178
rect 16578 19136 16634 19145
rect 16578 19071 16634 19080
rect 16264 18652 16436 18680
rect 16212 18634 16264 18640
rect 16224 18086 16252 18634
rect 16592 18358 16620 19071
rect 16580 18352 16632 18358
rect 16486 18320 16542 18329
rect 16580 18294 16632 18300
rect 16486 18255 16542 18264
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17542 16252 18022
rect 16316 17814 16344 18090
rect 16500 17814 16528 18255
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16684 17762 16712 21950
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 21078 16804 21286
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 18834 16804 19654
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16764 18080 16816 18086
rect 16762 18048 16764 18057
rect 16816 18048 16818 18057
rect 16762 17983 16818 17992
rect 16580 17740 16632 17746
rect 16684 17734 16804 17762
rect 16580 17682 16632 17688
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16212 17128 16264 17134
rect 16500 17105 16528 17546
rect 16212 17070 16264 17076
rect 16486 17096 16542 17105
rect 16224 16454 16252 17070
rect 16304 17060 16356 17066
rect 16486 17031 16542 17040
rect 16304 17002 16356 17008
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16224 15366 16252 15846
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15094 16252 15302
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16224 14074 16252 15030
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16224 7274 16252 13806
rect 16316 12481 16344 17002
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16408 14249 16436 16118
rect 16592 15026 16620 17682
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16394 14240 16450 14249
rect 16394 14175 16450 14184
rect 16500 13394 16528 14418
rect 16592 14278 16620 14962
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16488 13388 16540 13394
rect 16540 13348 16620 13376
rect 16488 13330 16540 13336
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16302 12472 16358 12481
rect 16302 12407 16358 12416
rect 16500 12170 16528 12854
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16316 11286 16344 12106
rect 16500 11898 16528 12106
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16486 11656 16542 11665
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16408 10130 16436 11630
rect 16592 11626 16620 13348
rect 16486 11591 16488 11600
rect 16540 11591 16542 11600
rect 16580 11620 16632 11626
rect 16488 11562 16540 11568
rect 16580 11562 16632 11568
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16500 10062 16528 10474
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 8945 16344 9522
rect 16302 8936 16358 8945
rect 16302 8871 16358 8880
rect 16592 8566 16620 10950
rect 16684 10810 16712 17614
rect 16776 16726 16804 17734
rect 16868 17513 16896 21830
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16960 19174 16988 21354
rect 17052 20806 17080 21490
rect 17040 20800 17092 20806
rect 17038 20768 17040 20777
rect 17092 20768 17094 20777
rect 17038 20703 17094 20712
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 17542 16988 19110
rect 17052 18766 17080 19178
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17052 17542 17080 18566
rect 17144 18034 17172 22335
rect 17236 20534 17264 23462
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17328 21486 17356 22986
rect 17420 21486 17448 23666
rect 17512 23254 17540 26200
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17500 23248 17552 23254
rect 17500 23190 17552 23196
rect 17604 23118 17632 23802
rect 17696 23322 17724 24006
rect 17788 23322 17816 26302
rect 17866 26200 17922 26302
rect 17972 26302 18290 26330
rect 17972 26246 18000 26302
rect 17960 26240 18012 26246
rect 18234 26200 18290 26302
rect 18602 26200 18658 27000
rect 18970 26200 19026 27000
rect 19338 26200 19394 27000
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 17960 26182 18012 26188
rect 18616 25537 18644 26200
rect 18984 25809 19012 26200
rect 19352 26081 19380 26200
rect 19628 26160 19656 26250
rect 19706 26200 19762 27000
rect 20074 26330 20130 27000
rect 19812 26302 20130 26330
rect 19720 26160 19748 26200
rect 19812 26178 19840 26302
rect 20074 26200 20130 26302
rect 20166 26344 20222 26353
rect 20442 26330 20498 27000
rect 20810 26330 20866 27000
rect 20222 26302 20498 26330
rect 20166 26279 20222 26288
rect 20442 26200 20498 26302
rect 20732 26302 20866 26330
rect 20732 26217 20760 26302
rect 20718 26208 20774 26217
rect 19628 26132 19748 26160
rect 19800 26172 19852 26178
rect 20810 26200 20866 26302
rect 21178 26200 21234 27000
rect 21270 26752 21326 26761
rect 21546 26738 21602 27000
rect 21326 26710 21602 26738
rect 21270 26687 21326 26696
rect 21546 26200 21602 26710
rect 21914 26200 21970 27000
rect 22282 26200 22338 27000
rect 22376 26376 22428 26382
rect 22650 26330 22706 27000
rect 23018 26330 23074 27000
rect 22428 26324 22706 26330
rect 22376 26318 22706 26324
rect 22388 26302 22706 26318
rect 22650 26200 22706 26302
rect 22756 26302 23074 26330
rect 20718 26143 20774 26152
rect 19800 26114 19852 26120
rect 19338 26072 19394 26081
rect 19338 26007 19394 26016
rect 18970 25800 19026 25809
rect 18970 25735 19026 25744
rect 18602 25528 18658 25537
rect 18602 25463 18658 25472
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17866 23352 17922 23361
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17776 23316 17828 23322
rect 17866 23287 17922 23296
rect 17776 23258 17828 23264
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17512 22094 17540 23054
rect 17592 22976 17644 22982
rect 17592 22918 17644 22924
rect 17604 22438 17632 22918
rect 17696 22710 17724 23258
rect 17880 23186 17908 23287
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17684 22704 17736 22710
rect 17684 22646 17736 22652
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17696 22234 17724 22646
rect 17788 22438 17816 23122
rect 17972 23118 18000 23598
rect 18340 23322 18368 24210
rect 18420 23792 18472 23798
rect 18420 23734 18472 23740
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 17960 23112 18012 23118
rect 17880 23060 17960 23066
rect 17880 23054 18012 23060
rect 17880 23038 18000 23054
rect 18340 23050 18368 23258
rect 18328 23044 18380 23050
rect 17880 22778 17908 23038
rect 18328 22986 18380 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17512 22066 17632 22094
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17512 21486 17540 21898
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17408 21480 17460 21486
rect 17500 21480 17552 21486
rect 17408 21422 17460 21428
rect 17498 21448 17500 21457
rect 17552 21448 17554 21457
rect 17224 20528 17276 20534
rect 17224 20470 17276 20476
rect 17420 20380 17448 21422
rect 17498 21383 17554 21392
rect 17604 21146 17632 22066
rect 17972 21894 18000 22714
rect 18326 22536 18382 22545
rect 18432 22506 18460 23734
rect 18616 23322 18644 25230
rect 20720 25084 20772 25090
rect 20720 25026 20772 25032
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18708 23050 18736 24210
rect 18800 24177 18828 24210
rect 19628 24206 19656 24346
rect 19524 24200 19576 24206
rect 18786 24168 18842 24177
rect 19524 24142 19576 24148
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 18786 24103 18842 24112
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18326 22471 18382 22480
rect 18420 22500 18472 22506
rect 18234 22128 18290 22137
rect 18234 22063 18236 22072
rect 18288 22063 18290 22072
rect 18340 22094 18368 22471
rect 18420 22442 18472 22448
rect 18340 22066 18460 22094
rect 18236 22034 18288 22040
rect 17684 21888 17736 21894
rect 17960 21888 18012 21894
rect 17684 21830 17736 21836
rect 17880 21848 17960 21876
rect 17696 21690 17724 21830
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17880 21434 17908 21848
rect 17960 21830 18012 21836
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18432 21486 18460 22066
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18708 21690 18736 22034
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 17788 21406 17908 21434
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18604 21412 18656 21418
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17696 20618 17724 21014
rect 17788 20777 17816 21406
rect 18604 21354 18656 21360
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17774 20768 17830 20777
rect 17774 20703 17830 20712
rect 17696 20590 17816 20618
rect 17236 20352 17448 20380
rect 17236 18902 17264 20352
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17328 18426 17356 19246
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 18193 17264 18226
rect 17222 18184 17278 18193
rect 17222 18119 17278 18128
rect 17144 18006 17356 18034
rect 17328 17814 17356 18006
rect 17420 17921 17448 19654
rect 17604 19334 17632 19926
rect 17604 19306 17724 19334
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17406 17912 17462 17921
rect 17406 17847 17462 17856
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 16948 17536 17000 17542
rect 16854 17504 16910 17513
rect 16948 17478 17000 17484
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16854 17439 16910 17448
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16776 15978 16804 16526
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16776 15638 16804 15914
rect 16868 15706 16896 16934
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14822 16804 14962
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14618 16804 14758
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13258 16804 13670
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16868 12850 16896 15506
rect 16960 13841 16988 17138
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17038 15736 17094 15745
rect 17038 15671 17094 15680
rect 17052 15473 17080 15671
rect 17038 15464 17094 15473
rect 17038 15399 17094 15408
rect 17144 14822 17172 16526
rect 17236 15570 17264 17274
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17224 15428 17276 15434
rect 17328 15416 17356 16458
rect 17276 15388 17356 15416
rect 17224 15370 17276 15376
rect 17236 15094 17264 15370
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 17236 14346 17264 15030
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17236 14074 17264 14282
rect 17512 14074 17540 18022
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 16946 13832 17002 13841
rect 16946 13767 17002 13776
rect 17040 13796 17092 13802
rect 17040 13738 17092 13744
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12434 16896 12786
rect 16776 12406 16896 12434
rect 16946 12472 17002 12481
rect 16946 12407 17002 12416
rect 16776 12306 16804 12406
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16960 11778 16988 12407
rect 16868 11750 16988 11778
rect 16762 11248 16818 11257
rect 16762 11183 16818 11192
rect 16776 11150 16804 11183
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16868 10810 16896 11750
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16960 11150 16988 11630
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16868 10674 16896 10746
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16684 9926 16712 9998
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16960 9722 16988 10406
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 17052 9586 17080 13738
rect 17236 13258 17264 14010
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12918 17264 13194
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12776 17276 12782
rect 17276 12736 17356 12764
rect 17224 12718 17276 12724
rect 17144 10810 17172 12718
rect 17328 12434 17356 12736
rect 17236 12406 17356 12434
rect 17236 11286 17264 12406
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17328 10674 17356 12038
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17132 10464 17184 10470
rect 17130 10432 17132 10441
rect 17184 10432 17186 10441
rect 17130 10367 17186 10376
rect 17144 10062 17172 10367
rect 17222 10296 17278 10305
rect 17222 10231 17224 10240
rect 17276 10231 17278 10240
rect 17224 10202 17276 10208
rect 17420 10130 17448 13874
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17512 13530 17540 13738
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17498 13424 17554 13433
rect 17498 13359 17554 13368
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16868 6390 16896 9318
rect 17512 7954 17540 13359
rect 17604 12102 17632 18770
rect 17696 17542 17724 19306
rect 17788 18698 17816 20590
rect 17880 19310 17908 21286
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18340 21010 18368 21082
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18432 19990 18460 21014
rect 18616 20942 18644 21354
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18708 20602 18736 20946
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18708 20505 18736 20538
rect 18694 20496 18750 20505
rect 18694 20431 18750 20440
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18156 19718 18184 19926
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18432 19417 18460 19790
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18418 19408 18474 19417
rect 18418 19343 18474 19352
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17866 19000 17922 19009
rect 17866 18935 17922 18944
rect 17880 18766 17908 18935
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17788 18290 17816 18634
rect 18328 18624 18380 18630
rect 18380 18584 18460 18612
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17202 17724 17478
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 12782 17724 17138
rect 17788 17066 17816 17614
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17202 18368 17682
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17776 17060 17828 17066
rect 17776 17002 17828 17008
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17880 16794 17908 16934
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17880 16522 17908 16730
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17788 12889 17816 14418
rect 17880 14074 17908 14894
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18432 14090 18460 18584
rect 18524 18222 18552 19654
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18524 15881 18552 18158
rect 18510 15872 18566 15881
rect 18510 15807 18566 15816
rect 18616 14618 18644 18158
rect 18708 16697 18736 18226
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18604 14612 18656 14618
rect 18656 14572 18736 14600
rect 18604 14554 18656 14560
rect 17868 14068 17920 14074
rect 18432 14062 18644 14090
rect 17868 14010 17920 14016
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17774 12880 17830 12889
rect 17774 12815 17830 12824
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17880 12481 17908 13806
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18234 12880 18290 12889
rect 18234 12815 18290 12824
rect 17866 12472 17922 12481
rect 17866 12407 17922 12416
rect 18248 12374 18276 12815
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17696 11082 17724 12242
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11830 17908 12106
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 18340 11286 18368 13330
rect 18432 12986 18460 13942
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18340 10606 18368 11018
rect 18432 10674 18460 12650
rect 18524 12238 18552 13670
rect 18616 12986 18644 14062
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18432 10266 18460 10474
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 17604 9926 17632 10202
rect 18326 10160 18382 10169
rect 18326 10095 18382 10104
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17880 7546 17908 8366
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18340 7546 18368 10095
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18432 7478 18460 8774
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 17236 6254 17264 6802
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 18524 5778 18552 12038
rect 18616 9654 18644 12786
rect 18708 11218 18736 14572
rect 18800 13394 18828 24006
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18984 22778 19012 22918
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18984 22030 19012 22374
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 19076 21894 19104 22170
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18892 18222 18920 19654
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18892 15473 18920 18158
rect 19076 18154 19104 21490
rect 19168 18698 19196 24006
rect 19432 23520 19484 23526
rect 19430 23488 19432 23497
rect 19484 23488 19486 23497
rect 19430 23423 19486 23432
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19430 23080 19486 23089
rect 19248 22500 19300 22506
rect 19248 22442 19300 22448
rect 19260 22409 19288 22442
rect 19246 22400 19302 22409
rect 19246 22335 19302 22344
rect 19352 22094 19380 23054
rect 19430 23015 19486 23024
rect 19444 22982 19472 23015
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19536 22778 19564 24142
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19812 23050 19840 23122
rect 19800 23044 19852 23050
rect 19800 22986 19852 22992
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19892 22704 19944 22710
rect 19892 22646 19944 22652
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19352 22066 19656 22094
rect 19352 21350 19380 22066
rect 19628 22030 19656 22066
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20392 19300 20398
rect 19352 20380 19380 20878
rect 19300 20352 19380 20380
rect 19248 20334 19300 20340
rect 19260 18766 19288 20334
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19514 19472 19654
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19340 19168 19392 19174
rect 19338 19136 19340 19145
rect 19432 19168 19484 19174
rect 19392 19136 19394 19145
rect 19432 19110 19484 19116
rect 19338 19071 19394 19080
rect 19444 18902 19472 19110
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18760 19300 18766
rect 19352 18737 19380 18770
rect 19248 18702 19300 18708
rect 19338 18728 19394 18737
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18984 17105 19012 17546
rect 18970 17096 19026 17105
rect 18970 17031 19026 17040
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16590 19012 16934
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18878 15464 18934 15473
rect 18878 15399 18934 15408
rect 18984 15162 19012 16050
rect 19076 16046 19104 18090
rect 19260 17746 19288 18702
rect 19338 18663 19394 18672
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19248 16992 19300 16998
rect 19168 16952 19248 16980
rect 19168 16794 19196 16952
rect 19248 16934 19300 16940
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18892 14414 18920 14758
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18786 13152 18842 13161
rect 18786 13087 18842 13096
rect 18800 12617 18828 13087
rect 18786 12608 18842 12617
rect 18786 12543 18842 12552
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18786 11112 18842 11121
rect 18786 11047 18842 11056
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18800 9450 18828 11047
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18786 9208 18842 9217
rect 18786 9143 18842 9152
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18708 7410 18736 9046
rect 18800 8838 18828 9143
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18892 8430 18920 11494
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18984 4078 19012 15098
rect 19076 14414 19104 15982
rect 19168 15706 19196 16594
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 16046 19288 16526
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19352 15609 19380 18090
rect 19444 16522 19472 18634
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19338 15600 19394 15609
rect 19338 15535 19394 15544
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19076 14006 19104 14350
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19076 12102 19104 12582
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19076 10810 19104 11630
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19062 10568 19118 10577
rect 19062 10503 19064 10512
rect 19116 10503 19118 10512
rect 19064 10474 19116 10480
rect 19168 10418 19196 15302
rect 19340 14952 19392 14958
rect 19392 14912 19472 14940
rect 19340 14894 19392 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14550 19288 14826
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19260 13734 19288 14486
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19076 10390 19196 10418
rect 19076 8430 19104 10390
rect 19154 9208 19210 9217
rect 19154 9143 19156 9152
rect 19208 9143 19210 9152
rect 19156 9114 19208 9120
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19260 6798 19288 12718
rect 19352 10538 19380 14214
rect 19444 14074 19472 14912
rect 19536 14618 19564 21966
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21729 19656 21830
rect 19614 21720 19670 21729
rect 19614 21655 19670 21664
rect 19720 21486 19748 22578
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19628 18902 19656 21422
rect 19720 21010 19748 21422
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19706 20904 19762 20913
rect 19706 20839 19708 20848
rect 19760 20839 19762 20848
rect 19708 20810 19760 20816
rect 19904 20777 19932 22646
rect 19996 22234 20024 24754
rect 20732 24410 20760 25026
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20074 24304 20130 24313
rect 20074 24239 20130 24248
rect 20088 24206 20116 24239
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20088 23089 20116 24142
rect 20824 23866 20852 25434
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20916 23798 20944 24074
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20720 23520 20772 23526
rect 20824 23497 20852 23598
rect 20720 23462 20772 23468
rect 20810 23488 20866 23497
rect 20074 23080 20130 23089
rect 20074 23015 20130 23024
rect 20732 22574 20760 23462
rect 20810 23423 20866 23432
rect 20916 23186 20944 23734
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20916 22778 20944 23122
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19890 20768 19946 20777
rect 19890 20703 19946 20712
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19720 19786 19748 20198
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19628 16266 19656 17478
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 16658 19748 17002
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19628 16238 19748 16266
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19444 12306 19472 14010
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11898 19472 12038
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11150 19472 11834
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19430 9752 19486 9761
rect 19430 9687 19486 9696
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 9081 19380 9318
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19444 8974 19472 9687
rect 19432 8968 19484 8974
rect 19352 8928 19432 8956
rect 19352 7342 19380 8928
rect 19432 8910 19484 8916
rect 19430 8120 19486 8129
rect 19430 8055 19432 8064
rect 19484 8055 19486 8064
rect 19432 8026 19484 8032
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6458 19288 6734
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19536 5710 19564 12582
rect 19628 10266 19656 16050
rect 19720 13410 19748 16238
rect 19812 14482 19840 18022
rect 19904 15502 19932 18158
rect 19996 15570 20024 21286
rect 20364 21010 20392 22442
rect 20732 22438 20760 22510
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20534 22264 20590 22273
rect 20534 22199 20590 22208
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20602 20208 20810
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20180 20058 20208 20538
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19982 15464 20038 15473
rect 19982 15399 20038 15408
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 13841 19840 14214
rect 19798 13832 19854 13841
rect 19798 13767 19854 13776
rect 19720 13382 19840 13410
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 11830 19748 13262
rect 19812 12986 19840 13382
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19798 12336 19854 12345
rect 19798 12271 19854 12280
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19720 10674 19748 10950
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19628 8974 19656 9658
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19720 7410 19748 10474
rect 19812 9450 19840 12271
rect 19904 11121 19932 15302
rect 19996 13977 20024 15399
rect 19982 13968 20038 13977
rect 19982 13903 20038 13912
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19996 12986 20024 13194
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19996 11286 20024 12106
rect 20088 12102 20116 17682
rect 20180 17270 20208 19246
rect 20272 17649 20300 20334
rect 20364 19145 20392 20946
rect 20548 20058 20576 22199
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20720 21888 20772 21894
rect 20718 21856 20720 21865
rect 20772 21856 20774 21865
rect 20718 21791 20774 21800
rect 21100 21690 21128 21898
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20626 21176 20682 21185
rect 20626 21111 20682 21120
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20350 19136 20406 19145
rect 20350 19071 20406 19080
rect 20640 18698 20668 21111
rect 20732 21078 20760 21354
rect 20824 21321 20852 21490
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 20810 21312 20866 21321
rect 20810 21247 20866 21256
rect 20810 21176 20866 21185
rect 20810 21111 20812 21120
rect 20864 21111 20866 21120
rect 20812 21082 20864 21088
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 19922 20852 20334
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20258 17640 20314 17649
rect 20258 17575 20314 17584
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20272 16402 20300 17138
rect 20352 16448 20404 16454
rect 20272 16396 20352 16402
rect 20272 16390 20404 16396
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20272 16374 20392 16390
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20180 13530 20208 15982
rect 20272 15570 20300 16374
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 20272 11218 20300 14418
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 19984 11144 20036 11150
rect 19890 11112 19946 11121
rect 19984 11086 20036 11092
rect 19890 11047 19946 11056
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19996 8906 20024 11086
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19798 8664 19854 8673
rect 19798 8599 19800 8608
rect 19852 8599 19854 8608
rect 19800 8570 19852 8576
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 20088 3058 20116 11018
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20180 9722 20208 10406
rect 20272 10062 20300 10406
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20364 9994 20392 14486
rect 20456 13433 20484 16390
rect 20548 16046 20576 18566
rect 20732 18290 20760 19246
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20640 17202 20668 17614
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20732 16114 20760 18226
rect 20824 18154 20852 19654
rect 20916 19553 20944 21422
rect 21008 19689 21036 21490
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20994 19680 21050 19689
rect 20994 19615 21050 19624
rect 20902 19544 20958 19553
rect 20902 19479 20958 19488
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20824 16590 20852 16934
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20548 15638 20576 15846
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20640 15337 20668 15846
rect 20626 15328 20682 15337
rect 20626 15263 20682 15272
rect 20534 15192 20590 15201
rect 20534 15127 20590 15136
rect 20442 13424 20498 13433
rect 20442 13359 20498 13368
rect 20548 12850 20576 15127
rect 20720 15020 20772 15026
rect 20824 15008 20852 16526
rect 20772 14980 20852 15008
rect 20720 14962 20772 14968
rect 20732 14618 20760 14962
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14074 20852 14350
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20916 13920 20944 19382
rect 21100 19009 21128 20878
rect 21192 20777 21220 26200
rect 21730 25256 21786 25265
rect 21730 25191 21786 25200
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21560 22778 21588 23258
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21376 22094 21404 22374
rect 21376 22066 21496 22094
rect 21284 21978 21312 22034
rect 21376 21978 21404 22066
rect 21284 21950 21404 21978
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21468 21434 21496 22066
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21652 21690 21680 21966
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21272 20800 21324 20806
rect 21178 20768 21234 20777
rect 21272 20742 21324 20748
rect 21178 20703 21234 20712
rect 21284 19718 21312 20742
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21086 19000 21142 19009
rect 21086 18935 21142 18944
rect 21192 18290 21220 19246
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20824 13892 20944 13920
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20536 12708 20588 12714
rect 20536 12650 20588 12656
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11898 20484 12106
rect 20548 12102 20576 12650
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20442 11248 20498 11257
rect 20442 11183 20498 11192
rect 20352 9988 20404 9994
rect 20352 9930 20404 9936
rect 20350 9888 20406 9897
rect 20350 9823 20406 9832
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20364 9586 20392 9823
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20180 8838 20208 8978
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8090 20208 8774
rect 20456 8498 20484 11183
rect 20548 11150 20576 12038
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20534 9616 20590 9625
rect 20534 9551 20590 9560
rect 20548 9450 20576 9551
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20272 6458 20300 8434
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20456 6322 20484 8298
rect 20640 7886 20668 12786
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20732 7410 20760 13670
rect 20824 11218 20852 13892
rect 21008 12782 21036 17546
rect 21100 14074 21128 18022
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21008 12345 21036 12378
rect 20994 12336 21050 12345
rect 20994 12271 21050 12280
rect 21100 12238 21128 13767
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21192 11778 21220 15982
rect 21284 15570 21312 19450
rect 21376 17116 21404 21422
rect 21468 21406 21680 21434
rect 21548 21344 21600 21350
rect 21454 21312 21510 21321
rect 21548 21286 21600 21292
rect 21454 21247 21510 21256
rect 21468 20466 21496 21247
rect 21560 20602 21588 21286
rect 21652 20913 21680 21406
rect 21638 20904 21694 20913
rect 21638 20839 21694 20848
rect 21652 20618 21680 20839
rect 21744 20777 21772 25191
rect 21822 22808 21878 22817
rect 21822 22743 21878 22752
rect 21730 20768 21786 20777
rect 21730 20703 21786 20712
rect 21548 20596 21600 20602
rect 21652 20590 21772 20618
rect 21548 20538 21600 20544
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21468 19961 21496 19994
rect 21454 19952 21510 19961
rect 21454 19887 21510 19896
rect 21456 19780 21508 19786
rect 21560 19768 21588 20198
rect 21508 19740 21588 19768
rect 21456 19722 21508 19728
rect 21468 18204 21496 19722
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21560 18358 21588 19178
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21468 18176 21588 18204
rect 21456 17128 21508 17134
rect 21376 17088 21456 17116
rect 21456 17070 21508 17076
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21376 15570 21404 16390
rect 21468 15570 21496 17070
rect 21560 16017 21588 18176
rect 21546 16008 21602 16017
rect 21652 15978 21680 19654
rect 21744 19242 21772 20590
rect 21836 19417 21864 22743
rect 21928 22234 21956 26200
rect 22296 24954 22324 26200
rect 22560 25424 22612 25430
rect 22560 25366 22612 25372
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22468 24880 22520 24886
rect 22098 24848 22154 24857
rect 22468 24822 22520 24828
rect 22098 24783 22154 24792
rect 22112 24342 22140 24783
rect 22282 24712 22338 24721
rect 22282 24647 22338 24656
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22020 23322 22048 23734
rect 22112 23633 22140 24006
rect 22204 23746 22232 24142
rect 22296 23866 22324 24647
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 24138 22416 24550
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22204 23718 22324 23746
rect 22296 23662 22324 23718
rect 22284 23656 22336 23662
rect 22098 23624 22154 23633
rect 22284 23598 22336 23604
rect 22098 23559 22154 23568
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 22020 22030 22048 23258
rect 22296 23186 22324 23598
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22388 23066 22416 24074
rect 22296 23038 22416 23066
rect 22296 22710 22324 23038
rect 22480 22930 22508 24822
rect 22388 22902 22508 22930
rect 22284 22704 22336 22710
rect 22112 22664 22284 22692
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 21185 21956 21286
rect 21914 21176 21970 21185
rect 21914 21111 21970 21120
rect 22020 21078 22048 21830
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21928 20058 21956 20946
rect 22006 20904 22062 20913
rect 22006 20839 22062 20848
rect 22020 20806 22048 20839
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21822 19408 21878 19417
rect 21822 19343 21878 19352
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21744 17610 21772 18702
rect 22020 18358 22048 20538
rect 22112 20534 22140 22664
rect 22284 22646 22336 22652
rect 22284 22500 22336 22506
rect 22284 22442 22336 22448
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22112 19514 22140 20470
rect 22204 19961 22232 21626
rect 22296 20330 22324 22442
rect 22388 20913 22416 22902
rect 22468 22568 22520 22574
rect 22468 22510 22520 22516
rect 22480 22137 22508 22510
rect 22466 22128 22522 22137
rect 22466 22063 22522 22072
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22374 20904 22430 20913
rect 22480 20874 22508 21830
rect 22572 20942 22600 25366
rect 22756 25129 22784 26302
rect 23018 26200 23074 26302
rect 23386 26200 23442 27000
rect 24490 26200 24546 27000
rect 24858 26200 24914 27000
rect 25226 26200 25282 27000
rect 25778 26480 25834 26489
rect 25778 26415 25834 26424
rect 22742 25120 22798 25129
rect 22742 25055 22798 25064
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22848 23866 22876 24210
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21146 22692 21830
rect 22756 21690 22784 22918
rect 23308 22574 23336 23122
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22374 20839 22430 20848
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22190 19952 22246 19961
rect 22190 19887 22246 19896
rect 22388 19718 22416 20402
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22112 19174 22140 19450
rect 22480 19417 22508 19450
rect 22466 19408 22522 19417
rect 22466 19343 22522 19352
rect 22284 19304 22336 19310
rect 22572 19258 22600 20266
rect 22756 20233 22784 21354
rect 22848 21010 22876 22374
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 21554 23336 22510
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22836 21004 22888 21010
rect 22836 20946 22888 20952
rect 22940 20641 22968 21082
rect 22926 20632 22982 20641
rect 22926 20567 22982 20576
rect 23308 20466 23336 21490
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22742 20224 22798 20233
rect 22742 20159 22798 20168
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22284 19246 22336 19252
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21744 17270 21772 17546
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21744 16998 21772 17206
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21546 15943 21602 15952
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21100 11750 21220 11778
rect 21100 11558 21128 11750
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20810 11112 20866 11121
rect 20810 11047 20866 11056
rect 20824 8974 20852 11047
rect 21008 10130 21036 11154
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 21100 10010 21128 11494
rect 21192 11286 21220 11630
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21008 9982 21128 10010
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20810 8800 20866 8809
rect 20810 8735 20866 8744
rect 20824 8634 20852 8735
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20916 8090 20944 9590
rect 21008 9353 21036 9982
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 20994 9344 21050 9353
rect 20994 9279 21050 9288
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 7744 20864 7750
rect 21008 7732 21036 8842
rect 21100 7750 21128 9590
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21192 9489 21220 9522
rect 21178 9480 21234 9489
rect 21178 9415 21234 9424
rect 20864 7704 21036 7732
rect 21088 7744 21140 7750
rect 20812 7686 20864 7692
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6798 20668 7142
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20916 6458 20944 7704
rect 21088 7686 21140 7692
rect 21192 6662 21220 9415
rect 21284 8634 21312 15370
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21376 14074 21404 14282
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21468 12782 21496 13942
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21376 12628 21404 12718
rect 21376 12600 21496 12628
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21376 10130 21404 12242
rect 21468 10674 21496 12600
rect 21560 10792 21588 15302
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21652 13870 21680 14282
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21652 13530 21680 13806
rect 21744 13734 21772 16118
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21836 14822 21864 15370
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21928 13920 21956 18090
rect 22020 15094 22048 18294
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17746 22232 18022
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22098 17096 22154 17105
rect 22098 17031 22154 17040
rect 22112 16046 22140 17031
rect 22296 16794 22324 19246
rect 22480 19230 22600 19258
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22098 15192 22154 15201
rect 22098 15127 22154 15136
rect 22112 15094 22140 15127
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22020 14414 22048 15030
rect 22204 14793 22232 15982
rect 22296 15026 22324 16594
rect 22388 15910 22416 18566
rect 22480 17678 22508 19230
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18442 22600 19110
rect 22664 18630 22692 19314
rect 22756 19174 22784 19722
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22572 18414 22692 18442
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22480 17270 22508 17614
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22572 17202 22600 18022
rect 22664 17542 22692 18414
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22190 14784 22246 14793
rect 22190 14719 22246 14728
rect 22296 14618 22324 14962
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21836 13892 21956 13920
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21640 13252 21692 13258
rect 21640 13194 21692 13200
rect 21652 12646 21680 13194
rect 21836 13161 21864 13892
rect 22192 13864 22244 13870
rect 21928 13812 22192 13818
rect 22296 13818 22324 14554
rect 22244 13812 22324 13818
rect 21928 13790 22324 13812
rect 21928 13394 21956 13790
rect 22098 13696 22154 13705
rect 22098 13631 22154 13640
rect 22006 13424 22062 13433
rect 21916 13388 21968 13394
rect 22006 13359 22062 13368
rect 21916 13330 21968 13336
rect 21822 13152 21878 13161
rect 21822 13087 21878 13096
rect 21928 12850 21956 13330
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21652 11830 21680 12582
rect 21824 12368 21876 12374
rect 21822 12336 21824 12345
rect 21876 12336 21878 12345
rect 21928 12306 21956 12786
rect 21822 12271 21878 12280
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 21640 11824 21692 11830
rect 21640 11766 21692 11772
rect 21652 11558 21680 11766
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21652 11286 21680 11494
rect 21730 11384 21786 11393
rect 21730 11319 21786 11328
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21744 11150 21772 11319
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21836 11082 21864 11562
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21560 10764 21864 10792
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21560 9926 21588 10610
rect 21640 9988 21692 9994
rect 21640 9930 21692 9936
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21362 9752 21418 9761
rect 21362 9687 21418 9696
rect 21376 8956 21404 9687
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21454 9344 21510 9353
rect 21454 9279 21510 9288
rect 21468 9058 21496 9279
rect 21560 9178 21588 9522
rect 21652 9178 21680 9930
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21468 9030 21588 9058
rect 21560 8974 21588 9030
rect 21548 8968 21600 8974
rect 21376 8928 21496 8956
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21376 8362 21404 8570
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21284 6458 21312 6734
rect 21468 6730 21496 8928
rect 21548 8910 21600 8916
rect 21744 6730 21772 9454
rect 21836 9217 21864 10764
rect 21822 9208 21878 9217
rect 21822 9143 21878 9152
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21836 6390 21864 6666
rect 21824 6384 21876 6390
rect 21824 6326 21876 6332
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 19444 2650 19472 2926
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 6920 2440 6972 2446
rect 6748 2388 6920 2394
rect 6748 2382 6972 2388
rect 6748 2366 6960 2382
rect 6748 800 6776 2366
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 4014
rect 21928 3534 21956 11018
rect 22020 10538 22048 13359
rect 22112 12646 22140 13631
rect 22282 13560 22338 13569
rect 22282 13495 22338 13504
rect 22296 13161 22324 13495
rect 22282 13152 22338 13161
rect 22282 13087 22338 13096
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22112 11354 22140 11834
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22008 9648 22060 9654
rect 22112 9602 22140 9658
rect 22060 9596 22140 9602
rect 22008 9590 22140 9596
rect 22020 9574 22140 9590
rect 22098 9480 22154 9489
rect 22008 9444 22060 9450
rect 22098 9415 22100 9424
rect 22008 9386 22060 9392
rect 22152 9415 22154 9424
rect 22100 9386 22152 9392
rect 22020 9353 22048 9386
rect 22006 9344 22062 9353
rect 22006 9279 22062 9288
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22112 7886 22140 8570
rect 22204 8022 22232 11698
rect 22296 10810 22324 12718
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 4146 22140 6598
rect 22204 6322 22232 7686
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22296 5386 22324 10610
rect 22388 10606 22416 15846
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22480 10282 22508 17070
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22572 15960 22600 17002
rect 22652 16992 22704 16998
rect 22650 16960 22652 16969
rect 22704 16960 22706 16969
rect 22650 16895 22706 16904
rect 22650 16552 22706 16561
rect 22650 16487 22652 16496
rect 22704 16487 22706 16496
rect 22652 16458 22704 16464
rect 22652 15972 22704 15978
rect 22572 15932 22652 15960
rect 22652 15914 22704 15920
rect 22756 15858 22784 18770
rect 22664 15830 22784 15858
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22572 15162 22600 15302
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22558 15056 22614 15065
rect 22558 14991 22614 15000
rect 22572 14113 22600 14991
rect 22558 14104 22614 14113
rect 22558 14039 22614 14048
rect 22558 13832 22614 13841
rect 22558 13767 22614 13776
rect 22572 13138 22600 13767
rect 22664 13394 22692 15830
rect 22848 15042 22876 20402
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19922 23336 20402
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19378 23336 19858
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23032 18601 23060 18634
rect 23018 18592 23074 18601
rect 23018 18527 23074 18536
rect 23308 18426 23336 19314
rect 23400 19281 23428 26200
rect 23756 25560 23808 25566
rect 23756 25502 23808 25508
rect 23480 25016 23532 25022
rect 23480 24958 23532 24964
rect 23492 22710 23520 24958
rect 23570 24304 23626 24313
rect 23570 24239 23626 24248
rect 23664 24268 23716 24274
rect 23584 23066 23612 24239
rect 23664 24210 23716 24216
rect 23676 23730 23704 24210
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23676 23322 23704 23666
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23676 23186 23704 23258
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23584 23038 23704 23066
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23492 21049 23520 22102
rect 23478 21040 23534 21049
rect 23478 20975 23534 20984
rect 23584 20806 23612 22918
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23676 19922 23704 23038
rect 23768 22098 23796 25502
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23860 22030 23888 25298
rect 24400 25220 24452 25226
rect 24400 25162 24452 25168
rect 24216 25152 24268 25158
rect 24216 25094 24268 25100
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 24044 23225 24072 23462
rect 24030 23216 24086 23225
rect 24030 23151 24032 23160
rect 24084 23151 24086 23160
rect 24032 23122 24084 23128
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23952 22094 23980 22918
rect 24136 22166 24164 24006
rect 24124 22160 24176 22166
rect 24124 22102 24176 22108
rect 23952 22066 24072 22094
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23386 19272 23442 19281
rect 23386 19207 23442 19216
rect 23386 19136 23442 19145
rect 23386 19071 23442 19080
rect 23400 18970 23428 19071
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23400 18426 23428 18566
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23308 18086 23336 18362
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23386 17912 23442 17921
rect 23386 17847 23388 17856
rect 23440 17847 23442 17856
rect 23388 17818 23440 17824
rect 22928 17808 22980 17814
rect 22926 17776 22928 17785
rect 23480 17808 23532 17814
rect 22980 17776 22982 17785
rect 22926 17711 22982 17720
rect 23400 17756 23480 17762
rect 23400 17750 23532 17756
rect 23400 17734 23520 17750
rect 22926 17640 22982 17649
rect 22926 17575 22928 17584
rect 22980 17575 22982 17584
rect 22928 17546 22980 17552
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23216 17377 23244 17478
rect 23202 17368 23258 17377
rect 23202 17303 23258 17312
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22940 17134 22968 17206
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23124 16114 23152 16730
rect 23308 16697 23336 17478
rect 23400 16998 23428 17734
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 17542 23520 17614
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23386 16824 23442 16833
rect 23386 16759 23442 16768
rect 23294 16688 23350 16697
rect 23294 16623 23350 16632
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23400 15994 23428 16759
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23308 15966 23428 15994
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 23032 15162 23060 15574
rect 23308 15434 23336 15966
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23400 15337 23428 15846
rect 23492 15638 23520 16050
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23492 15201 23520 15370
rect 23478 15192 23534 15201
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23296 15156 23348 15162
rect 23478 15127 23534 15136
rect 23296 15098 23348 15104
rect 22756 15014 22876 15042
rect 22756 14498 22784 15014
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22848 14618 22876 14826
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22756 14470 23244 14498
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 23216 14226 23244 14470
rect 23308 14385 23336 15098
rect 23386 14648 23442 14657
rect 23386 14583 23442 14592
rect 23400 14550 23428 14583
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23584 14482 23612 19654
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23676 18737 23704 19246
rect 23662 18728 23718 18737
rect 23662 18663 23718 18672
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23294 14376 23350 14385
rect 23676 14362 23704 18566
rect 23768 17746 23796 21830
rect 24044 20890 24072 22066
rect 24044 20862 24164 20890
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23860 16250 23888 20198
rect 23952 19514 23980 20742
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24044 18698 24072 20742
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24044 16538 24072 18158
rect 24136 16561 24164 20862
rect 24228 20398 24256 25094
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17270 24256 17478
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24228 16590 24256 17206
rect 24216 16584 24268 16590
rect 23952 16510 24072 16538
rect 24122 16552 24178 16561
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23768 15366 23796 15642
rect 23846 15464 23902 15473
rect 23846 15399 23902 15408
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 15094 23796 15302
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23294 14311 23350 14320
rect 23492 14334 23704 14362
rect 23386 14240 23442 14249
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22572 13110 22692 13138
rect 22558 13016 22614 13025
rect 22558 12951 22614 12960
rect 22572 12918 22600 12951
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22664 12730 22692 13110
rect 22572 12702 22692 12730
rect 22572 10674 22600 12702
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22664 12102 22692 12582
rect 22848 12434 22876 14214
rect 23216 14198 23336 14226
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 22940 13734 22968 13903
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22928 13388 22980 13394
rect 22980 13348 23060 13376
rect 22928 13330 22980 13336
rect 23032 12646 23060 13348
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 12442 23336 14198
rect 23386 14175 23442 14184
rect 23400 14006 23428 14175
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23296 12436 23348 12442
rect 22848 12406 22968 12434
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22388 10266 22508 10282
rect 22376 10260 22508 10266
rect 22428 10254 22508 10260
rect 22376 10202 22428 10208
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22388 7886 22416 9318
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22480 6866 22508 9522
rect 22572 8838 22600 10406
rect 22664 9994 22692 11290
rect 22756 11150 22784 11630
rect 22940 11540 22968 12406
rect 23296 12378 23348 12384
rect 23400 12186 23428 12650
rect 22848 11512 22968 11540
rect 23308 12158 23428 12186
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22664 9722 22692 9930
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22848 9042 22876 11512
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 10470 23336 12158
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11082 23428 12038
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23216 9926 23244 10134
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9466 23244 9862
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23216 9438 23336 9466
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22664 7546 22692 8910
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 22204 5358 22324 5386
rect 22204 4622 22232 5358
rect 22282 5264 22338 5273
rect 22282 5199 22284 5208
rect 22336 5199 22338 5208
rect 22284 5170 22336 5176
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 1170 22048 3402
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22112 2009 22140 2586
rect 22098 2000 22154 2009
rect 22098 1935 22154 1944
rect 22204 1601 22232 4014
rect 22756 3602 22784 5578
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22296 3058 22324 3334
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23308 2582 23336 9438
rect 23400 7818 23428 9930
rect 23492 9654 23520 14334
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23584 9330 23612 14214
rect 23768 13682 23796 14758
rect 23492 9302 23612 9330
rect 23676 13654 23796 13682
rect 23492 7954 23520 9302
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 7812 23440 7818
rect 23388 7754 23440 7760
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23492 6186 23520 7346
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23400 4622 23428 5782
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 23676 4146 23704 13654
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23768 12782 23796 13330
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 8974 23796 12718
rect 23860 12714 23888 15399
rect 23952 13530 23980 16510
rect 24216 16526 24268 16532
rect 24122 16487 24178 16496
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 16046 24072 16390
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 24044 15502 24072 15982
rect 24228 15706 24256 16526
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24032 15496 24084 15502
rect 24320 15450 24348 22714
rect 24412 21593 24440 25162
rect 24504 23089 24532 26200
rect 25594 26072 25650 26081
rect 25594 26007 25650 26016
rect 24766 25664 24822 25673
rect 24766 25599 24822 25608
rect 24780 24614 24808 25599
rect 24950 25256 25006 25265
rect 24950 25191 25006 25200
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24780 23798 24808 24550
rect 24964 24206 24992 25191
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24964 24070 24992 24142
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 24768 23792 24820 23798
rect 24768 23734 24820 23740
rect 24490 23080 24546 23089
rect 24490 23015 24546 23024
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24780 22574 24808 22986
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24398 21584 24454 21593
rect 24780 21554 24808 22510
rect 24398 21519 24454 21528
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24780 21350 24808 21490
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24032 15438 24084 15444
rect 24136 15422 24348 15450
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 24044 14346 24072 15302
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 24136 13682 24164 15422
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24320 14958 24348 15302
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24216 14340 24268 14346
rect 24216 14282 24268 14288
rect 24228 13938 24256 14282
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24044 13654 24164 13682
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 23952 12850 23980 13466
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23848 12708 23900 12714
rect 23848 12650 23900 12656
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23860 11354 23888 12106
rect 23952 12102 23980 12582
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23768 5234 23796 7482
rect 23860 6322 23888 9590
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23952 3058 23980 9862
rect 24044 9518 24072 13654
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24136 12238 24164 13466
rect 24228 13462 24256 13874
rect 24412 13530 24440 17070
rect 24504 14958 24532 19858
rect 24596 18057 24624 20742
rect 24780 20534 24808 21286
rect 24872 21010 24900 24006
rect 24952 23588 25004 23594
rect 24952 23530 25004 23536
rect 24964 21690 24992 23530
rect 25136 23520 25188 23526
rect 25136 23462 25188 23468
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 24964 21457 24992 21626
rect 24950 21448 25006 21457
rect 24950 21383 25006 21392
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24768 20528 24820 20534
rect 24820 20488 24992 20516
rect 24768 20470 24820 20476
rect 24858 19952 24914 19961
rect 24858 19887 24860 19896
rect 24912 19887 24914 19896
rect 24860 19858 24912 19864
rect 24964 19854 24992 20488
rect 25056 20058 25084 22918
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24858 19544 24914 19553
rect 24858 19479 24914 19488
rect 24872 19334 24900 19479
rect 24964 19446 24992 19790
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24780 19306 24900 19334
rect 24674 19000 24730 19009
rect 24674 18935 24730 18944
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24596 17338 24624 17614
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24492 14952 24544 14958
rect 24544 14900 24624 14906
rect 24492 14894 24624 14900
rect 24504 14878 24624 14894
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24504 13870 24532 14418
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24216 13456 24268 13462
rect 24268 13416 24348 13444
rect 24216 13398 24268 13404
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24124 12232 24176 12238
rect 24124 12174 24176 12180
rect 24032 9512 24084 9518
rect 24032 9454 24084 9460
rect 24228 8362 24256 13126
rect 24320 12850 24348 13416
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12170 24348 12786
rect 24308 12164 24360 12170
rect 24308 12106 24360 12112
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24504 7886 24532 13806
rect 24596 11150 24624 14878
rect 24688 14074 24716 18935
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24780 12288 24808 19306
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24964 18329 24992 18566
rect 24950 18320 25006 18329
rect 24950 18255 25006 18264
rect 25056 16697 25084 19654
rect 25148 18698 25176 23462
rect 25412 22500 25464 22506
rect 25412 22442 25464 22448
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25240 19514 25268 22034
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25240 18358 25268 19314
rect 25332 18970 25360 22374
rect 25424 21010 25452 22442
rect 25412 21004 25464 21010
rect 25412 20946 25464 20952
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 19786 25452 20742
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25516 19310 25544 24006
rect 25608 22030 25636 26007
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 20806 25636 21966
rect 25792 21962 25820 26415
rect 25962 24440 26018 24449
rect 25962 24375 26018 24384
rect 25870 22672 25926 22681
rect 25870 22607 25926 22616
rect 25780 21956 25832 21962
rect 25780 21898 25832 21904
rect 25792 21690 25820 21898
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25596 20052 25648 20058
rect 25596 19994 25648 20000
rect 25504 19304 25556 19310
rect 25504 19246 25556 19252
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25504 18896 25556 18902
rect 25504 18838 25556 18844
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25240 17270 25268 18294
rect 25228 17264 25280 17270
rect 25228 17206 25280 17212
rect 25042 16688 25098 16697
rect 25042 16623 25098 16632
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24952 14000 25004 14006
rect 24950 13968 24952 13977
rect 25004 13968 25006 13977
rect 24950 13903 25006 13912
rect 24952 13796 25004 13802
rect 24952 13738 25004 13744
rect 24688 12260 24808 12288
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24688 10849 24716 12260
rect 24766 12200 24822 12209
rect 24964 12186 24992 13738
rect 25056 13161 25084 14010
rect 25042 13152 25098 13161
rect 25042 13087 25098 13096
rect 25148 12986 25176 16594
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25240 16182 25268 16390
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25134 12608 25190 12617
rect 25134 12543 25190 12552
rect 24964 12158 25084 12186
rect 24766 12135 24822 12144
rect 24674 10840 24730 10849
rect 24674 10775 24730 10784
rect 24780 10606 24808 12135
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24858 11384 24914 11393
rect 25056 11354 25084 12158
rect 25148 11830 25176 12543
rect 25240 12322 25268 14758
rect 25332 13190 25360 18566
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25424 17338 25452 18362
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25424 13705 25452 17138
rect 25410 13696 25466 13705
rect 25410 13631 25466 13640
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25332 12442 25360 12922
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25240 12294 25360 12322
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 24858 11319 24914 11328
rect 25044 11348 25096 11354
rect 24872 11218 24900 11319
rect 25044 11290 25096 11296
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 25134 10976 25190 10985
rect 25134 10911 25190 10920
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24768 10600 24820 10606
rect 24872 10577 24900 10678
rect 24768 10542 24820 10548
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 24766 10160 24822 10169
rect 24766 10095 24822 10104
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24490 6896 24546 6905
rect 24490 6831 24492 6840
rect 24544 6831 24546 6840
rect 24492 6802 24544 6808
rect 24596 5370 24624 9862
rect 24780 8430 24808 10095
rect 25148 9654 25176 10911
rect 25136 9648 25188 9654
rect 25136 9590 25188 9596
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24872 9042 24900 9279
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 24950 8528 25006 8537
rect 24950 8463 24952 8472
rect 25004 8463 25006 8472
rect 24952 8434 25004 8440
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24858 8120 24914 8129
rect 24858 8055 24914 8064
rect 24872 7954 24900 8055
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24674 6896 24730 6905
rect 24674 6831 24676 6840
rect 24728 6831 24730 6840
rect 24676 6802 24728 6808
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 25148 7478 25176 8871
rect 25240 8090 25268 12174
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24950 6896 25006 6905
rect 24950 6831 25006 6840
rect 24964 6798 24992 6831
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 25056 5710 25084 7142
rect 25332 6882 25360 12294
rect 25424 9178 25452 13262
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25410 7984 25466 7993
rect 25410 7919 25466 7928
rect 25148 6854 25360 6882
rect 25044 5704 25096 5710
rect 24950 5672 25006 5681
rect 25044 5646 25096 5652
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24860 5296 24912 5302
rect 24766 5264 24822 5273
rect 24860 5238 24912 5244
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23296 2576 23348 2582
rect 23296 2518 23348 2524
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 22190 1592 22246 1601
rect 22190 1527 22246 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2450
rect 24596 2446 24624 4966
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24688 3534 24716 4422
rect 24780 4078 24808 5199
rect 24872 4865 24900 5238
rect 24858 4856 24914 4865
rect 24858 4791 24914 4800
rect 25148 4690 25176 6854
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25240 6186 25268 6734
rect 25320 6724 25372 6730
rect 25320 6666 25372 6672
rect 25228 6180 25280 6186
rect 25228 6122 25280 6128
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25134 4040 25190 4049
rect 24952 4004 25004 4010
rect 25134 3975 25190 3984
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24952 3460 25004 3466
rect 24952 3402 25004 3408
rect 24964 3233 24992 3402
rect 24950 3224 25006 3233
rect 24950 3159 25006 3168
rect 25148 3126 25176 3975
rect 25240 3738 25268 6122
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 25332 3194 25360 6666
rect 25424 5846 25452 7919
rect 25516 6458 25544 18838
rect 25608 14074 25636 19994
rect 25700 19825 25728 20198
rect 25686 19816 25742 19825
rect 25686 19751 25742 19760
rect 25700 18834 25728 19751
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25700 13870 25728 18770
rect 25792 18426 25820 21626
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25778 17368 25834 17377
rect 25778 17303 25834 17312
rect 25792 16454 25820 17303
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25412 5840 25464 5846
rect 25412 5782 25464 5788
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25516 4457 25544 4490
rect 25502 4448 25558 4457
rect 25502 4383 25558 4392
rect 25608 3942 25636 13806
rect 25686 13696 25742 13705
rect 25686 13631 25742 13640
rect 25700 12753 25728 13631
rect 25686 12744 25742 12753
rect 25686 12679 25742 12688
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 5914 25728 12582
rect 25792 10062 25820 15506
rect 25884 14006 25912 22607
rect 25976 22522 26004 24375
rect 26054 23624 26110 23633
rect 26110 23582 26464 23610
rect 26054 23559 26110 23568
rect 26054 23216 26110 23225
rect 26110 23174 26372 23202
rect 26054 23151 26110 23160
rect 25976 22494 26280 22522
rect 26054 22400 26110 22409
rect 26054 22335 26110 22344
rect 25962 20360 26018 20369
rect 25962 20295 26018 20304
rect 25976 16538 26004 20295
rect 26068 20058 26096 22335
rect 26252 22094 26280 22494
rect 26160 22066 26280 22094
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 26054 19952 26110 19961
rect 26054 19887 26110 19896
rect 26068 19378 26096 19887
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 26068 17202 26096 18906
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26160 16658 26188 22066
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 25976 16510 26188 16538
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25872 14000 25924 14006
rect 25872 13942 25924 13948
rect 25976 13938 26004 16390
rect 26056 16380 26108 16386
rect 26056 16322 26108 16328
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25872 13864 25924 13870
rect 25924 13812 26004 13818
rect 25872 13806 26004 13812
rect 25884 13790 26004 13806
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25700 4826 25728 5850
rect 25884 5778 25912 13194
rect 25976 11665 26004 13790
rect 25962 11656 26018 11665
rect 25962 11591 26018 11600
rect 25964 9240 26016 9246
rect 25962 9208 25964 9217
rect 26016 9208 26018 9217
rect 25962 9143 26018 9152
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25688 4820 25740 4826
rect 25688 4762 25740 4768
rect 25976 4758 26004 9143
rect 26068 9081 26096 16322
rect 26160 14550 26188 16510
rect 26148 14544 26200 14550
rect 26148 14486 26200 14492
rect 26252 11898 26280 19314
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26054 9072 26110 9081
rect 26054 9007 26110 9016
rect 26344 8906 26372 23174
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 26436 8022 26464 23582
rect 26792 23044 26844 23050
rect 26792 22986 26844 22992
rect 26804 22094 26832 22986
rect 26884 22228 26936 22234
rect 26884 22170 26936 22176
rect 26712 22066 26832 22094
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26528 10538 26556 19450
rect 26516 10532 26568 10538
rect 26516 10474 26568 10480
rect 26620 9246 26648 21830
rect 26712 18154 26740 22066
rect 26792 21004 26844 21010
rect 26792 20946 26844 20952
rect 26700 18148 26752 18154
rect 26700 18090 26752 18096
rect 26700 17060 26752 17066
rect 26700 17002 26752 17008
rect 26608 9240 26660 9246
rect 26608 9182 26660 9188
rect 26712 8634 26740 17002
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 26424 8016 26476 8022
rect 26424 7958 26476 7964
rect 26804 5846 26832 20946
rect 26896 9450 26924 22170
rect 26884 9444 26936 9450
rect 26884 9386 26936 9392
rect 26792 5840 26844 5846
rect 26792 5782 26844 5788
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25136 3120 25188 3126
rect 25136 3062 25188 3068
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24950 2408 25006 2417
rect 24950 2343 24952 2352
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 25056 785 25084 2926
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 1490 24792 1546 24848
rect 1582 23044 1638 23080
rect 1582 23024 1584 23044
rect 1584 23024 1636 23044
rect 1636 23024 1638 23044
rect 2134 26152 2190 26208
rect 2042 23840 2098 23896
rect 2134 18808 2190 18864
rect 1858 16108 1914 16144
rect 1858 16088 1860 16108
rect 1860 16088 1912 16108
rect 1912 16088 1914 16108
rect 2502 26152 2558 26208
rect 2042 16496 2098 16552
rect 2318 14456 2374 14512
rect 2318 13932 2374 13968
rect 2318 13912 2320 13932
rect 2320 13912 2372 13932
rect 2372 13912 2374 13932
rect 2134 13388 2190 13424
rect 2134 13368 2136 13388
rect 2136 13368 2188 13388
rect 2188 13368 2190 13388
rect 3146 25880 3202 25936
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2962 24112 3018 24168
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2778 17040 2834 17096
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3514 21256 3570 21312
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 3974 23568 4030 23624
rect 3698 21936 3754 21992
rect 3698 20712 3754 20768
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2778 15020 2834 15056
rect 2778 15000 2780 15020
rect 2780 15000 2832 15020
rect 2832 15000 2834 15020
rect 3974 22616 4030 22672
rect 3882 19352 3938 19408
rect 3790 15156 3846 15192
rect 3790 15136 3792 15156
rect 3792 15136 3844 15156
rect 3844 15136 3846 15156
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2134 12844 2190 12880
rect 2134 12824 2136 12844
rect 2136 12824 2188 12844
rect 2188 12824 2190 12844
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 3514 12280 3570 12336
rect 1950 11600 2006 11656
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 4434 23568 4490 23624
rect 4342 23160 4398 23216
rect 4158 22072 4214 22128
rect 4250 21936 4306 21992
rect 4342 18284 4398 18320
rect 4342 18264 4344 18284
rect 4344 18264 4396 18284
rect 4396 18264 4398 18284
rect 4802 22480 4858 22536
rect 4526 21936 4582 21992
rect 4526 19488 4582 19544
rect 4802 21120 4858 21176
rect 4894 19896 4950 19952
rect 5446 26832 5502 26888
rect 4342 14728 4398 14784
rect 4894 15680 4950 15736
rect 5262 18672 5318 18728
rect 5170 18264 5226 18320
rect 5446 19080 5502 19136
rect 5446 15816 5502 15872
rect 5814 25472 5870 25528
rect 5722 21800 5778 21856
rect 6090 21936 6146 21992
rect 5630 16632 5686 16688
rect 5538 14456 5594 14512
rect 5446 13232 5502 13288
rect 5354 12688 5410 12744
rect 3974 10648 4030 10704
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 1766 9560 1822 9616
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 5906 17040 5962 17096
rect 6734 22616 6790 22672
rect 7010 25064 7066 25120
rect 7010 21800 7066 21856
rect 6826 20460 6882 20496
rect 6826 20440 6828 20460
rect 6828 20440 6880 20460
rect 6880 20440 6882 20460
rect 6550 19780 6606 19816
rect 6550 19760 6552 19780
rect 6552 19760 6604 19780
rect 6604 19760 6606 19780
rect 6182 17620 6184 17640
rect 6184 17620 6236 17640
rect 6236 17620 6238 17640
rect 6182 17584 6238 17620
rect 6366 16224 6422 16280
rect 6918 17212 6920 17232
rect 6920 17212 6972 17232
rect 6972 17212 6974 17232
rect 6918 17176 6974 17212
rect 6734 15000 6790 15056
rect 5814 11192 5870 11248
rect 5630 11056 5686 11112
rect 4986 7928 5042 7984
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 6366 13504 6422 13560
rect 6550 12824 6606 12880
rect 7930 25608 7986 25664
rect 7930 25200 7986 25256
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7470 20848 7526 20904
rect 7470 20032 7526 20088
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 8574 24928 8630 24984
rect 9218 25200 9274 25256
rect 9126 23432 9182 23488
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8298 21528 8354 21584
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 8390 20576 8446 20632
rect 7838 20304 7894 20360
rect 7746 20168 7802 20224
rect 7286 19488 7342 19544
rect 7194 15544 7250 15600
rect 7470 17992 7526 18048
rect 8114 19896 8170 19952
rect 8298 19896 8354 19952
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7654 18400 7710 18456
rect 7562 17720 7618 17776
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8390 18400 8446 18456
rect 8206 18148 8262 18184
rect 8206 18128 8208 18148
rect 8208 18128 8260 18148
rect 8260 18128 8262 18148
rect 8666 20712 8722 20768
rect 9126 22208 9182 22264
rect 8298 17992 8354 18048
rect 8298 17856 8354 17912
rect 7286 14320 7342 14376
rect 7010 12144 7066 12200
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8482 17448 8538 17504
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8206 15564 8262 15600
rect 8206 15544 8208 15564
rect 8208 15544 8260 15564
rect 8260 15544 8262 15564
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 8390 15136 8446 15192
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7838 13932 7894 13968
rect 7838 13912 7840 13932
rect 7840 13912 7892 13932
rect 7892 13912 7894 13932
rect 7930 13776 7986 13832
rect 8666 17312 8722 17368
rect 8666 16496 8722 16552
rect 8758 14864 8814 14920
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 8298 12416 8354 12472
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7378 11736 7434 11792
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 8942 19624 8998 19680
rect 9034 18400 9090 18456
rect 9402 20984 9458 21040
rect 9402 20576 9458 20632
rect 9310 20168 9366 20224
rect 9310 19624 9366 19680
rect 9402 19252 9404 19272
rect 9404 19252 9456 19272
rect 9456 19252 9458 19272
rect 9402 19216 9458 19252
rect 9126 15952 9182 16008
rect 9678 23840 9734 23896
rect 9770 23724 9826 23760
rect 9770 23704 9772 23724
rect 9772 23704 9824 23724
rect 9824 23704 9826 23724
rect 9862 23568 9918 23624
rect 10230 23568 10286 23624
rect 10046 23432 10102 23488
rect 9586 20168 9642 20224
rect 9678 16788 9734 16824
rect 9678 16768 9680 16788
rect 9680 16768 9732 16788
rect 9732 16768 9734 16788
rect 9770 15408 9826 15464
rect 10322 17176 10378 17232
rect 11150 22344 11206 22400
rect 10966 19080 11022 19136
rect 11058 17176 11114 17232
rect 9678 13912 9734 13968
rect 9678 13776 9734 13832
rect 9586 13504 9642 13560
rect 9678 13096 9734 13152
rect 9586 12824 9642 12880
rect 9218 12144 9274 12200
rect 10138 14184 10194 14240
rect 12070 23296 12126 23352
rect 11150 16224 11206 16280
rect 11518 19624 11574 19680
rect 11426 18944 11482 19000
rect 11426 18672 11482 18728
rect 11242 15272 11298 15328
rect 11518 16768 11574 16824
rect 12438 23160 12494 23216
rect 12162 22208 12218 22264
rect 12070 20032 12126 20088
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13266 23160 13322 23216
rect 12806 22888 12862 22944
rect 12714 22344 12770 22400
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12530 20304 12586 20360
rect 12530 20032 12586 20088
rect 11794 15680 11850 15736
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12530 16632 12586 16688
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 14094 24792 14150 24848
rect 13818 23468 13820 23488
rect 13820 23468 13872 23488
rect 13872 23468 13874 23488
rect 13818 23432 13874 23468
rect 13634 21800 13690 21856
rect 13634 21292 13636 21312
rect 13636 21292 13688 21312
rect 13688 21292 13690 21312
rect 13634 21256 13690 21292
rect 13542 20304 13598 20360
rect 13174 19352 13230 19408
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13542 19080 13598 19136
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 14370 21664 14426 21720
rect 14922 25880 14978 25936
rect 14554 23432 14610 23488
rect 14646 22888 14702 22944
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13358 16768 13414 16824
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13726 15816 13782 15872
rect 14186 19624 14242 19680
rect 13634 13776 13690 13832
rect 13542 12552 13598 12608
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 14370 19352 14426 19408
rect 14370 18944 14426 19000
rect 14278 17740 14334 17776
rect 14278 17720 14280 17740
rect 14280 17720 14332 17740
rect 14332 17720 14334 17740
rect 13726 11464 13782 11520
rect 14554 20304 14610 20360
rect 15382 24384 15438 24440
rect 14738 17176 14794 17232
rect 14554 16632 14610 16688
rect 14738 16904 14794 16960
rect 14646 14592 14702 14648
rect 14554 14320 14610 14376
rect 14554 11328 14610 11384
rect 14554 11056 14610 11112
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 15382 23976 15438 24032
rect 15474 23604 15476 23624
rect 15476 23604 15528 23624
rect 15528 23604 15530 23624
rect 15474 23568 15530 23604
rect 15658 23432 15714 23488
rect 15566 21428 15568 21448
rect 15568 21428 15620 21448
rect 15620 21428 15622 21448
rect 15198 20576 15254 20632
rect 15566 21392 15622 21428
rect 15014 17992 15070 18048
rect 15106 15952 15162 16008
rect 15014 14340 15070 14376
rect 15014 14320 15016 14340
rect 15016 14320 15068 14340
rect 15068 14320 15070 14340
rect 15474 17176 15530 17232
rect 15198 14320 15254 14376
rect 15290 13776 15346 13832
rect 15014 11056 15070 11112
rect 17130 25608 17186 25664
rect 16762 25336 16818 25392
rect 15658 16768 15714 16824
rect 15566 16496 15622 16552
rect 15566 15952 15622 16008
rect 15658 14048 15714 14104
rect 15842 17332 15898 17368
rect 15842 17312 15844 17332
rect 15844 17312 15896 17332
rect 15896 17312 15898 17332
rect 15474 12300 15530 12336
rect 15474 12280 15476 12300
rect 15476 12280 15528 12300
rect 15528 12280 15530 12300
rect 15474 12164 15530 12200
rect 15474 12144 15476 12164
rect 15476 12144 15528 12164
rect 15528 12144 15530 12164
rect 15474 11736 15530 11792
rect 15290 10104 15346 10160
rect 15658 9596 15660 9616
rect 15660 9596 15712 9616
rect 15712 9596 15714 9616
rect 15658 9560 15714 9596
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 16210 23568 16266 23624
rect 16486 23196 16488 23216
rect 16488 23196 16540 23216
rect 16540 23196 16542 23216
rect 16486 23160 16542 23196
rect 16670 22752 16726 22808
rect 16302 22072 16358 22128
rect 16486 22072 16542 22128
rect 17130 23840 17186 23896
rect 16946 23160 17002 23216
rect 16946 22888 17002 22944
rect 17130 22652 17132 22672
rect 17132 22652 17184 22672
rect 17184 22652 17186 22672
rect 17130 22616 17186 22652
rect 17130 22344 17186 22400
rect 16486 21120 16542 21176
rect 16026 20032 16082 20088
rect 16486 20712 16542 20768
rect 16302 20576 16358 20632
rect 16578 20304 16634 20360
rect 16578 19080 16634 19136
rect 16486 18264 16542 18320
rect 16762 18028 16764 18048
rect 16764 18028 16816 18048
rect 16816 18028 16818 18048
rect 16762 17992 16818 18028
rect 16486 17040 16542 17096
rect 16394 14184 16450 14240
rect 16302 12416 16358 12472
rect 16486 11620 16542 11656
rect 16486 11600 16488 11620
rect 16488 11600 16540 11620
rect 16540 11600 16542 11620
rect 16302 8880 16358 8936
rect 17038 20748 17040 20768
rect 17040 20748 17092 20768
rect 17092 20748 17094 20768
rect 17038 20712 17094 20748
rect 20166 26288 20222 26344
rect 20718 26152 20774 26208
rect 21270 26696 21326 26752
rect 19338 26016 19394 26072
rect 18970 25744 19026 25800
rect 18602 25472 18658 25528
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17866 23296 17922 23352
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17498 21428 17500 21448
rect 17500 21428 17552 21448
rect 17552 21428 17554 21448
rect 17498 21392 17554 21428
rect 18326 22480 18382 22536
rect 18786 24112 18842 24168
rect 18234 22092 18290 22128
rect 18234 22072 18236 22092
rect 18236 22072 18288 22092
rect 18288 22072 18290 22092
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17774 20712 17830 20768
rect 17222 18128 17278 18184
rect 17406 17856 17462 17912
rect 16854 17448 16910 17504
rect 17038 15680 17094 15736
rect 17038 15408 17094 15464
rect 16946 13776 17002 13832
rect 16946 12416 17002 12472
rect 16762 11192 16818 11248
rect 17130 10412 17132 10432
rect 17132 10412 17184 10432
rect 17184 10412 17186 10432
rect 17130 10376 17186 10412
rect 17222 10260 17278 10296
rect 17222 10240 17224 10260
rect 17224 10240 17276 10260
rect 17276 10240 17278 10260
rect 17498 13368 17554 13424
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18694 20440 18750 20496
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18418 19352 18474 19408
rect 17866 18944 17922 19000
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18510 15816 18566 15872
rect 18694 16632 18750 16688
rect 17774 12824 17830 12880
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18234 12824 18290 12880
rect 17866 12416 17922 12472
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18326 10104 18382 10160
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 19430 23468 19432 23488
rect 19432 23468 19484 23488
rect 19484 23468 19486 23488
rect 19430 23432 19486 23468
rect 19246 22344 19302 22400
rect 19430 23024 19486 23080
rect 19338 19116 19340 19136
rect 19340 19116 19392 19136
rect 19392 19116 19394 19136
rect 19338 19080 19394 19116
rect 18970 17040 19026 17096
rect 18878 15408 18934 15464
rect 19338 18672 19394 18728
rect 18786 13096 18842 13152
rect 18786 12552 18842 12608
rect 18786 11056 18842 11112
rect 18786 9152 18842 9208
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19338 15544 19394 15600
rect 19062 10532 19118 10568
rect 19062 10512 19064 10532
rect 19064 10512 19116 10532
rect 19116 10512 19118 10532
rect 19154 9172 19210 9208
rect 19154 9152 19156 9172
rect 19156 9152 19208 9172
rect 19208 9152 19210 9172
rect 19614 21664 19670 21720
rect 19706 20868 19762 20904
rect 19706 20848 19708 20868
rect 19708 20848 19760 20868
rect 19760 20848 19762 20868
rect 20074 24248 20130 24304
rect 20074 23024 20130 23080
rect 20810 23432 20866 23488
rect 19890 20712 19946 20768
rect 19430 9696 19486 9752
rect 19338 9016 19394 9072
rect 19430 8084 19486 8120
rect 19430 8064 19432 8084
rect 19432 8064 19484 8084
rect 19484 8064 19486 8084
rect 20534 22208 20590 22264
rect 19982 15408 20038 15464
rect 19798 13776 19854 13832
rect 19798 12280 19854 12336
rect 19982 13912 20038 13968
rect 20718 21836 20720 21856
rect 20720 21836 20772 21856
rect 20772 21836 20774 21856
rect 20718 21800 20774 21836
rect 20626 21120 20682 21176
rect 20350 19080 20406 19136
rect 20810 21256 20866 21312
rect 20810 21140 20866 21176
rect 20810 21120 20812 21140
rect 20812 21120 20864 21140
rect 20864 21120 20866 21140
rect 20258 17584 20314 17640
rect 19890 11056 19946 11112
rect 19798 8628 19854 8664
rect 19798 8608 19800 8628
rect 19800 8608 19852 8628
rect 19852 8608 19854 8628
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 20994 19624 21050 19680
rect 20902 19488 20958 19544
rect 20626 15272 20682 15328
rect 20534 15136 20590 15192
rect 20442 13368 20498 13424
rect 21730 25200 21786 25256
rect 21178 20712 21234 20768
rect 21086 18944 21142 19000
rect 20442 11192 20498 11248
rect 20350 9832 20406 9888
rect 20534 9560 20590 9616
rect 21086 13776 21142 13832
rect 20994 12280 21050 12336
rect 21454 21256 21510 21312
rect 21638 20848 21694 20904
rect 21822 22752 21878 22808
rect 21730 20712 21786 20768
rect 21454 19896 21510 19952
rect 21546 15952 21602 16008
rect 22098 24792 22154 24848
rect 22282 24656 22338 24712
rect 22098 23568 22154 23624
rect 21914 21120 21970 21176
rect 22006 20848 22062 20904
rect 21822 19352 21878 19408
rect 22466 22072 22522 22128
rect 22374 20848 22430 20904
rect 25778 26424 25834 26480
rect 22742 25064 22798 25120
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22190 19896 22246 19952
rect 22466 19352 22522 19408
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22926 20576 22982 20632
rect 22742 20168 22798 20224
rect 20810 11056 20866 11112
rect 20810 8744 20866 8800
rect 20994 9288 21050 9344
rect 21178 9424 21234 9480
rect 22098 17040 22154 17096
rect 22098 15136 22154 15192
rect 22190 14728 22246 14784
rect 22098 13640 22154 13696
rect 22006 13368 22062 13424
rect 21822 13096 21878 13152
rect 21822 12316 21824 12336
rect 21824 12316 21876 12336
rect 21876 12316 21878 12336
rect 21822 12280 21878 12316
rect 21730 11328 21786 11384
rect 21362 9696 21418 9752
rect 21454 9288 21510 9344
rect 21822 9152 21878 9208
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22282 13504 22338 13560
rect 22282 13096 22338 13152
rect 22098 9444 22154 9480
rect 22098 9424 22100 9444
rect 22100 9424 22152 9444
rect 22152 9424 22154 9444
rect 22006 9288 22062 9344
rect 22650 16940 22652 16960
rect 22652 16940 22704 16960
rect 22704 16940 22706 16960
rect 22650 16904 22706 16940
rect 22650 16516 22706 16552
rect 22650 16496 22652 16516
rect 22652 16496 22704 16516
rect 22704 16496 22706 16516
rect 22558 15000 22614 15056
rect 22558 14048 22614 14104
rect 22558 13776 22614 13832
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 23018 18536 23074 18592
rect 23570 24248 23626 24304
rect 23478 20984 23534 21040
rect 24030 23180 24086 23216
rect 24030 23160 24032 23180
rect 24032 23160 24084 23180
rect 24084 23160 24086 23180
rect 23386 19216 23442 19272
rect 23386 19080 23442 19136
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17876 23442 17912
rect 23386 17856 23388 17876
rect 23388 17856 23440 17876
rect 23440 17856 23442 17876
rect 22926 17756 22928 17776
rect 22928 17756 22980 17776
rect 22980 17756 22982 17776
rect 22926 17720 22982 17756
rect 22926 17604 22982 17640
rect 22926 17584 22928 17604
rect 22928 17584 22980 17604
rect 22980 17584 22982 17604
rect 23202 17312 23258 17368
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 23386 16768 23442 16824
rect 23294 16632 23350 16688
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 23386 15272 23442 15328
rect 23478 15136 23534 15192
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 23386 14592 23442 14648
rect 23662 18672 23718 18728
rect 23294 14320 23350 14376
rect 23846 15408 23902 15464
rect 22558 12960 22614 13016
rect 22926 13912 22982 13968
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 23386 14184 23442 14240
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22282 5228 22338 5264
rect 22282 5208 22284 5228
rect 22284 5208 22336 5228
rect 22336 5208 22338 5228
rect 22098 1944 22154 2000
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24122 16496 24178 16552
rect 25594 26016 25650 26072
rect 24766 25608 24822 25664
rect 24950 25200 25006 25256
rect 24490 23024 24546 23080
rect 24398 21528 24454 21584
rect 24950 21392 25006 21448
rect 24858 19916 24914 19952
rect 24858 19896 24860 19916
rect 24860 19896 24912 19916
rect 24912 19896 24914 19916
rect 24858 19488 24914 19544
rect 24674 18944 24730 19000
rect 24582 17992 24638 18048
rect 24950 18264 25006 18320
rect 25962 24384 26018 24440
rect 25870 22616 25926 22672
rect 25042 16632 25098 16688
rect 24950 13948 24952 13968
rect 24952 13948 25004 13968
rect 25004 13948 25006 13968
rect 24950 13912 25006 13948
rect 24766 12144 24822 12200
rect 25042 13096 25098 13152
rect 25134 12552 25190 12608
rect 24674 10784 24730 10840
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24858 11328 24914 11384
rect 25410 13640 25466 13696
rect 25134 10920 25190 10976
rect 24858 10512 24914 10568
rect 24766 10104 24822 10160
rect 24490 6860 24546 6896
rect 24490 6840 24492 6860
rect 24492 6840 24544 6860
rect 24544 6840 24546 6860
rect 24858 9288 24914 9344
rect 25134 8880 25190 8936
rect 24950 8492 25006 8528
rect 24950 8472 24952 8492
rect 24952 8472 25004 8492
rect 25004 8472 25006 8492
rect 24858 8064 24914 8120
rect 24766 7656 24822 7712
rect 24674 6860 24730 6896
rect 24674 6840 24676 6860
rect 24676 6840 24728 6860
rect 24728 6840 24730 6860
rect 24674 6432 24730 6488
rect 24858 7248 24914 7304
rect 24950 6840 25006 6896
rect 24858 6024 24914 6080
rect 25410 7928 25466 7984
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24766 5208 24822 5264
rect 22190 1536 22246 1592
rect 22098 1128 22154 1184
rect 24858 4800 24914 4856
rect 25134 3984 25190 4040
rect 24950 3576 25006 3632
rect 24950 3168 25006 3224
rect 25686 19760 25742 19816
rect 25778 17312 25834 17368
rect 25502 4392 25558 4448
rect 25686 13640 25742 13696
rect 25686 12688 25742 12744
rect 26054 23568 26110 23624
rect 26054 23160 26110 23216
rect 26054 22344 26110 22400
rect 25962 20304 26018 20360
rect 26054 19896 26110 19952
rect 25962 11600 26018 11656
rect 25962 9188 25964 9208
rect 25964 9188 26016 9208
rect 26016 9188 26018 9208
rect 25962 9152 26018 9188
rect 26054 9016 26110 9072
rect 24858 2760 24914 2816
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 5441 26890 5507 26893
rect 16614 26890 16620 26892
rect 5441 26888 16620 26890
rect 5441 26832 5446 26888
rect 5502 26832 16620 26888
rect 5441 26830 16620 26832
rect 5441 26827 5507 26830
rect 16614 26828 16620 26830
rect 16684 26828 16690 26892
rect 10174 26692 10180 26756
rect 10244 26754 10250 26756
rect 21265 26754 21331 26757
rect 10244 26752 21331 26754
rect 10244 26696 21270 26752
rect 21326 26696 21331 26752
rect 10244 26694 21331 26696
rect 10244 26692 10250 26694
rect 21265 26691 21331 26694
rect 15326 26618 15332 26620
rect 2270 26558 15332 26618
rect 2129 26210 2195 26213
rect 2270 26210 2330 26558
rect 15326 26556 15332 26558
rect 15396 26556 15402 26620
rect 21398 26482 21404 26484
rect 2129 26208 2330 26210
rect 2129 26152 2134 26208
rect 2190 26152 2330 26208
rect 2129 26150 2330 26152
rect 2454 26422 21404 26482
rect 2454 26213 2514 26422
rect 21398 26420 21404 26422
rect 21468 26420 21474 26484
rect 25773 26482 25839 26485
rect 26200 26482 27000 26512
rect 25773 26480 27000 26482
rect 25773 26424 25778 26480
rect 25834 26424 27000 26480
rect 25773 26422 27000 26424
rect 25773 26419 25839 26422
rect 26200 26392 27000 26422
rect 2630 26284 2636 26348
rect 2700 26346 2706 26348
rect 20161 26346 20227 26349
rect 2700 26344 20227 26346
rect 2700 26288 20166 26344
rect 20222 26288 20227 26344
rect 2700 26286 20227 26288
rect 2700 26284 2706 26286
rect 20161 26283 20227 26286
rect 2454 26208 2563 26213
rect 2454 26152 2502 26208
rect 2558 26152 2563 26208
rect 2454 26150 2563 26152
rect 2129 26147 2195 26150
rect 2497 26147 2563 26150
rect 5390 26148 5396 26212
rect 5460 26210 5466 26212
rect 20713 26210 20779 26213
rect 5460 26208 20779 26210
rect 5460 26152 20718 26208
rect 20774 26152 20779 26208
rect 5460 26150 20779 26152
rect 5460 26148 5466 26150
rect 20713 26147 20779 26150
rect 5574 26012 5580 26076
rect 5644 26074 5650 26076
rect 19333 26074 19399 26077
rect 5644 26072 19399 26074
rect 5644 26016 19338 26072
rect 19394 26016 19399 26072
rect 5644 26014 19399 26016
rect 5644 26012 5650 26014
rect 19333 26011 19399 26014
rect 25589 26074 25655 26077
rect 26200 26074 27000 26104
rect 25589 26072 27000 26074
rect 25589 26016 25594 26072
rect 25650 26016 27000 26072
rect 25589 26014 27000 26016
rect 25589 26011 25655 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 3141 25938 3207 25941
rect 14917 25938 14983 25941
rect 0 25936 3207 25938
rect 0 25880 3146 25936
rect 3202 25880 3207 25936
rect 0 25878 3207 25880
rect 0 25848 800 25878
rect 3141 25875 3207 25878
rect 7606 25936 14983 25938
rect 7606 25880 14922 25936
rect 14978 25880 14983 25936
rect 7606 25878 14983 25880
rect 2262 25740 2268 25804
rect 2332 25802 2338 25804
rect 7606 25802 7666 25878
rect 14917 25875 14983 25878
rect 18965 25802 19031 25805
rect 2332 25742 7666 25802
rect 7790 25800 19031 25802
rect 7790 25744 18970 25800
rect 19026 25744 19031 25800
rect 7790 25742 19031 25744
rect 2332 25740 2338 25742
rect 6494 25604 6500 25668
rect 6564 25666 6570 25668
rect 7790 25666 7850 25742
rect 18965 25739 19031 25742
rect 6564 25606 7850 25666
rect 7925 25666 7991 25669
rect 17125 25666 17191 25669
rect 7925 25664 17191 25666
rect 7925 25608 7930 25664
rect 7986 25608 17130 25664
rect 17186 25608 17191 25664
rect 7925 25606 17191 25608
rect 6564 25604 6570 25606
rect 7925 25603 7991 25606
rect 17125 25603 17191 25606
rect 24761 25666 24827 25669
rect 26200 25666 27000 25696
rect 24761 25664 27000 25666
rect 24761 25608 24766 25664
rect 24822 25608 27000 25664
rect 24761 25606 27000 25608
rect 24761 25603 24827 25606
rect 26200 25576 27000 25606
rect 5809 25530 5875 25533
rect 18597 25530 18663 25533
rect 5809 25528 18663 25530
rect 5809 25472 5814 25528
rect 5870 25472 18602 25528
rect 18658 25472 18663 25528
rect 5809 25470 18663 25472
rect 5809 25467 5875 25470
rect 18597 25467 18663 25470
rect 7598 25332 7604 25396
rect 7668 25394 7674 25396
rect 16757 25394 16823 25397
rect 7668 25392 16823 25394
rect 7668 25336 16762 25392
rect 16818 25336 16823 25392
rect 7668 25334 16823 25336
rect 7668 25332 7674 25334
rect 16757 25331 16823 25334
rect 4654 25196 4660 25260
rect 4724 25258 4730 25260
rect 7925 25258 7991 25261
rect 4724 25256 7991 25258
rect 4724 25200 7930 25256
rect 7986 25200 7991 25256
rect 4724 25198 7991 25200
rect 4724 25196 4730 25198
rect 7925 25195 7991 25198
rect 9213 25258 9279 25261
rect 21725 25258 21791 25261
rect 9213 25256 21791 25258
rect 9213 25200 9218 25256
rect 9274 25200 21730 25256
rect 21786 25200 21791 25256
rect 9213 25198 21791 25200
rect 9213 25195 9279 25198
rect 21725 25195 21791 25198
rect 24945 25258 25011 25261
rect 26200 25258 27000 25288
rect 24945 25256 27000 25258
rect 24945 25200 24950 25256
rect 25006 25200 27000 25256
rect 24945 25198 27000 25200
rect 24945 25195 25011 25198
rect 26200 25168 27000 25198
rect 7005 25122 7071 25125
rect 22737 25122 22803 25125
rect 7005 25120 22803 25122
rect 7005 25064 7010 25120
rect 7066 25064 22742 25120
rect 22798 25064 22803 25120
rect 7005 25062 22803 25064
rect 7005 25059 7071 25062
rect 22737 25059 22803 25062
rect 8569 24986 8635 24989
rect 16430 24986 16436 24988
rect 8569 24984 16436 24986
rect 8569 24928 8574 24984
rect 8630 24928 16436 24984
rect 8569 24926 16436 24928
rect 8569 24923 8635 24926
rect 16430 24924 16436 24926
rect 16500 24924 16506 24988
rect 0 24850 800 24880
rect 1485 24850 1551 24853
rect 0 24848 1551 24850
rect 0 24792 1490 24848
rect 1546 24792 1551 24848
rect 0 24790 1551 24792
rect 0 24760 800 24790
rect 1485 24787 1551 24790
rect 5942 24788 5948 24852
rect 6012 24850 6018 24852
rect 14089 24850 14155 24853
rect 6012 24848 14155 24850
rect 6012 24792 14094 24848
rect 14150 24792 14155 24848
rect 6012 24790 14155 24792
rect 6012 24788 6018 24790
rect 14089 24787 14155 24790
rect 22093 24850 22159 24853
rect 26200 24850 27000 24880
rect 22093 24848 27000 24850
rect 22093 24792 22098 24848
rect 22154 24792 27000 24848
rect 22093 24790 27000 24792
rect 22093 24787 22159 24790
rect 26200 24760 27000 24790
rect 7782 24652 7788 24716
rect 7852 24714 7858 24716
rect 22277 24714 22343 24717
rect 7852 24712 22343 24714
rect 7852 24656 22282 24712
rect 22338 24656 22343 24712
rect 7852 24654 22343 24656
rect 7852 24652 7858 24654
rect 22277 24651 22343 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 15377 24442 15443 24445
rect 18454 24442 18460 24444
rect 15377 24440 18460 24442
rect 15377 24384 15382 24440
rect 15438 24384 18460 24440
rect 15377 24382 18460 24384
rect 15377 24379 15443 24382
rect 18454 24380 18460 24382
rect 18524 24380 18530 24444
rect 25957 24442 26023 24445
rect 26200 24442 27000 24472
rect 22050 24382 22754 24442
rect 11646 24244 11652 24308
rect 11716 24306 11722 24308
rect 20069 24306 20135 24309
rect 11716 24304 20135 24306
rect 11716 24248 20074 24304
rect 20130 24248 20135 24304
rect 11716 24246 20135 24248
rect 11716 24244 11722 24246
rect 20069 24243 20135 24246
rect 2957 24170 3023 24173
rect 2957 24168 8402 24170
rect 2957 24112 2962 24168
rect 3018 24112 8402 24168
rect 2957 24110 8402 24112
rect 2957 24107 3023 24110
rect 8342 24034 8402 24110
rect 8518 24108 8524 24172
rect 8588 24170 8594 24172
rect 18781 24170 18847 24173
rect 8588 24168 18847 24170
rect 8588 24112 18786 24168
rect 18842 24112 18847 24168
rect 8588 24110 18847 24112
rect 8588 24108 8594 24110
rect 18781 24107 18847 24110
rect 15377 24034 15443 24037
rect 8342 24032 15443 24034
rect 8342 23976 15382 24032
rect 15438 23976 15443 24032
rect 8342 23974 15443 23976
rect 15377 23971 15443 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 2037 23898 2103 23901
rect 9673 23898 9739 23901
rect 17125 23898 17191 23901
rect 2037 23896 3250 23898
rect 2037 23840 2042 23896
rect 2098 23840 3250 23896
rect 2037 23838 3250 23840
rect 2037 23835 2103 23838
rect 0 23762 800 23792
rect 3190 23762 3250 23838
rect 9673 23896 17191 23898
rect 9673 23840 9678 23896
rect 9734 23840 17130 23896
rect 17186 23840 17191 23896
rect 9673 23838 17191 23840
rect 9673 23835 9739 23838
rect 17125 23835 17191 23838
rect 9765 23762 9831 23765
rect 22050 23762 22110 24382
rect 22694 24306 22754 24382
rect 25957 24440 27000 24442
rect 25957 24384 25962 24440
rect 26018 24384 27000 24440
rect 25957 24382 27000 24384
rect 25957 24379 26023 24382
rect 26200 24352 27000 24382
rect 23565 24306 23631 24309
rect 22694 24304 23631 24306
rect 22694 24248 23570 24304
rect 23626 24248 23631 24304
rect 22694 24246 23631 24248
rect 23565 24243 23631 24246
rect 23974 23972 23980 24036
rect 24044 24034 24050 24036
rect 26200 24034 27000 24064
rect 24044 23974 27000 24034
rect 24044 23972 24050 23974
rect 26200 23944 27000 23974
rect 0 23702 2790 23762
rect 3190 23760 9831 23762
rect 3190 23704 9770 23760
rect 9826 23704 9831 23760
rect 3190 23702 9831 23704
rect 0 23672 800 23702
rect 2730 23626 2790 23702
rect 9765 23699 9831 23702
rect 12574 23702 22110 23762
rect 3969 23626 4035 23629
rect 2730 23624 4035 23626
rect 2730 23568 3974 23624
rect 4030 23568 4035 23624
rect 2730 23566 4035 23568
rect 3969 23563 4035 23566
rect 4429 23626 4495 23629
rect 9857 23626 9923 23629
rect 4429 23624 9923 23626
rect 4429 23568 4434 23624
rect 4490 23568 9862 23624
rect 9918 23568 9923 23624
rect 4429 23566 9923 23568
rect 4429 23563 4495 23566
rect 9857 23563 9923 23566
rect 10225 23626 10291 23629
rect 12574 23626 12634 23702
rect 10225 23624 12634 23626
rect 10225 23568 10230 23624
rect 10286 23568 12634 23624
rect 10225 23566 12634 23568
rect 12758 23566 13554 23626
rect 10225 23563 10291 23566
rect 5758 23428 5764 23492
rect 5828 23490 5834 23492
rect 9121 23490 9187 23493
rect 10041 23492 10107 23493
rect 9990 23490 9996 23492
rect 5828 23488 9187 23490
rect 5828 23432 9126 23488
rect 9182 23432 9187 23488
rect 5828 23430 9187 23432
rect 9950 23430 9996 23490
rect 10060 23488 10107 23492
rect 10102 23432 10107 23488
rect 5828 23428 5834 23430
rect 9121 23427 9187 23430
rect 9990 23428 9996 23430
rect 10060 23428 10107 23432
rect 10041 23427 10107 23428
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12065 23354 12131 23357
rect 12758 23354 12818 23566
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 12065 23352 12818 23354
rect 12065 23296 12070 23352
rect 12126 23296 12818 23352
rect 12065 23294 12818 23296
rect 13494 23354 13554 23566
rect 14958 23564 14964 23628
rect 15028 23626 15034 23628
rect 15469 23626 15535 23629
rect 15028 23624 15535 23626
rect 15028 23568 15474 23624
rect 15530 23568 15535 23624
rect 15028 23566 15535 23568
rect 15028 23564 15034 23566
rect 15469 23563 15535 23566
rect 16205 23626 16271 23629
rect 22093 23626 22159 23629
rect 16205 23624 22159 23626
rect 16205 23568 16210 23624
rect 16266 23568 22098 23624
rect 22154 23568 22159 23624
rect 16205 23566 22159 23568
rect 16205 23563 16271 23566
rect 22093 23563 22159 23566
rect 26049 23626 26115 23629
rect 26200 23626 27000 23656
rect 26049 23624 27000 23626
rect 26049 23568 26054 23624
rect 26110 23568 27000 23624
rect 26049 23566 27000 23568
rect 26049 23563 26115 23566
rect 26200 23536 27000 23566
rect 13813 23492 13879 23493
rect 13813 23490 13860 23492
rect 13768 23488 13860 23490
rect 13768 23432 13818 23488
rect 13768 23430 13860 23432
rect 13813 23428 13860 23430
rect 13924 23428 13930 23492
rect 14038 23428 14044 23492
rect 14108 23490 14114 23492
rect 14549 23490 14615 23493
rect 14108 23488 14615 23490
rect 14108 23432 14554 23488
rect 14610 23432 14615 23488
rect 14108 23430 14615 23432
rect 14108 23428 14114 23430
rect 13813 23427 13879 23428
rect 14549 23427 14615 23430
rect 15142 23428 15148 23492
rect 15212 23490 15218 23492
rect 15653 23490 15719 23493
rect 15212 23488 15719 23490
rect 15212 23432 15658 23488
rect 15714 23432 15719 23488
rect 15212 23430 15719 23432
rect 15212 23428 15218 23430
rect 15653 23427 15719 23430
rect 16062 23428 16068 23492
rect 16132 23490 16138 23492
rect 19425 23490 19491 23493
rect 16132 23488 19491 23490
rect 16132 23432 19430 23488
rect 19486 23432 19491 23488
rect 16132 23430 19491 23432
rect 16132 23428 16138 23430
rect 19425 23427 19491 23430
rect 19558 23428 19564 23492
rect 19628 23490 19634 23492
rect 20805 23490 20871 23493
rect 19628 23488 20871 23490
rect 19628 23432 20810 23488
rect 20866 23432 20871 23488
rect 19628 23430 20871 23432
rect 19628 23428 19634 23430
rect 20805 23427 20871 23430
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 17861 23354 17927 23357
rect 13494 23352 17927 23354
rect 13494 23296 17866 23352
rect 17922 23296 17927 23352
rect 13494 23294 17927 23296
rect 12065 23291 12131 23294
rect 17861 23291 17927 23294
rect 4337 23218 4403 23221
rect 12433 23218 12499 23221
rect 4337 23216 12499 23218
rect 4337 23160 4342 23216
rect 4398 23160 12438 23216
rect 12494 23160 12499 23216
rect 4337 23158 12499 23160
rect 4337 23155 4403 23158
rect 12433 23155 12499 23158
rect 12750 23156 12756 23220
rect 12820 23218 12826 23220
rect 13261 23218 13327 23221
rect 12820 23216 13327 23218
rect 12820 23160 13266 23216
rect 13322 23160 13327 23216
rect 12820 23158 13327 23160
rect 12820 23156 12826 23158
rect 13261 23155 13327 23158
rect 13670 23156 13676 23220
rect 13740 23218 13746 23220
rect 16481 23218 16547 23221
rect 13740 23216 16547 23218
rect 13740 23160 16486 23216
rect 16542 23160 16547 23216
rect 13740 23158 16547 23160
rect 13740 23156 13746 23158
rect 16481 23155 16547 23158
rect 16941 23218 17007 23221
rect 24025 23218 24091 23221
rect 16941 23216 24091 23218
rect 16941 23160 16946 23216
rect 17002 23160 24030 23216
rect 24086 23160 24091 23216
rect 16941 23158 24091 23160
rect 16941 23155 17007 23158
rect 24025 23155 24091 23158
rect 26049 23218 26115 23221
rect 26200 23218 27000 23248
rect 26049 23216 27000 23218
rect 26049 23160 26054 23216
rect 26110 23160 27000 23216
rect 26049 23158 27000 23160
rect 26049 23155 26115 23158
rect 26200 23128 27000 23158
rect 1577 23082 1643 23085
rect 19425 23082 19491 23085
rect 1577 23080 19491 23082
rect 1577 23024 1582 23080
rect 1638 23024 19430 23080
rect 19486 23024 19491 23080
rect 1577 23022 19491 23024
rect 1577 23019 1643 23022
rect 19425 23019 19491 23022
rect 20069 23082 20135 23085
rect 24485 23082 24551 23085
rect 20069 23080 24551 23082
rect 20069 23024 20074 23080
rect 20130 23024 24490 23080
rect 24546 23024 24551 23080
rect 20069 23022 24551 23024
rect 20069 23019 20135 23022
rect 24485 23019 24551 23022
rect 9254 22884 9260 22948
rect 9324 22946 9330 22948
rect 12801 22946 12867 22949
rect 9324 22944 12867 22946
rect 9324 22888 12806 22944
rect 12862 22888 12867 22944
rect 9324 22886 12867 22888
rect 9324 22884 9330 22886
rect 12801 22883 12867 22886
rect 14641 22946 14707 22949
rect 16941 22946 17007 22949
rect 14641 22944 17007 22946
rect 14641 22888 14646 22944
rect 14702 22888 16946 22944
rect 17002 22888 17007 22944
rect 14641 22886 17007 22888
rect 14641 22883 14707 22886
rect 16941 22883 17007 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 16665 22810 16731 22813
rect 21817 22810 21883 22813
rect 26200 22810 27000 22840
rect 16665 22808 17786 22810
rect 16665 22752 16670 22808
rect 16726 22752 17786 22808
rect 16665 22750 17786 22752
rect 16665 22747 16731 22750
rect 0 22674 800 22704
rect 3969 22674 4035 22677
rect 0 22672 4035 22674
rect 0 22616 3974 22672
rect 4030 22616 4035 22672
rect 0 22614 4035 22616
rect 0 22584 800 22614
rect 3969 22611 4035 22614
rect 6729 22674 6795 22677
rect 17125 22674 17191 22677
rect 6729 22672 17191 22674
rect 6729 22616 6734 22672
rect 6790 22616 17130 22672
rect 17186 22616 17191 22672
rect 6729 22614 17191 22616
rect 17726 22674 17786 22750
rect 21817 22808 27000 22810
rect 21817 22752 21822 22808
rect 21878 22752 27000 22808
rect 21817 22750 27000 22752
rect 21817 22747 21883 22750
rect 26200 22720 27000 22750
rect 25865 22674 25931 22677
rect 17726 22672 25931 22674
rect 17726 22616 25870 22672
rect 25926 22616 25931 22672
rect 17726 22614 25931 22616
rect 6729 22611 6795 22614
rect 17125 22611 17191 22614
rect 25865 22611 25931 22614
rect 4797 22538 4863 22541
rect 18321 22538 18387 22541
rect 4797 22536 18387 22538
rect 4797 22480 4802 22536
rect 4858 22480 18326 22536
rect 18382 22480 18387 22536
rect 4797 22478 18387 22480
rect 4797 22475 4863 22478
rect 18321 22475 18387 22478
rect 11145 22402 11211 22405
rect 12709 22402 12775 22405
rect 11145 22400 12775 22402
rect 11145 22344 11150 22400
rect 11206 22344 12714 22400
rect 12770 22344 12775 22400
rect 11145 22342 12775 22344
rect 11145 22339 11211 22342
rect 12709 22339 12775 22342
rect 16614 22340 16620 22404
rect 16684 22402 16690 22404
rect 17125 22402 17191 22405
rect 16684 22400 17191 22402
rect 16684 22344 17130 22400
rect 17186 22344 17191 22400
rect 16684 22342 17191 22344
rect 16684 22340 16690 22342
rect 17125 22339 17191 22342
rect 18638 22340 18644 22404
rect 18708 22402 18714 22404
rect 19241 22402 19307 22405
rect 18708 22400 19307 22402
rect 18708 22344 19246 22400
rect 19302 22344 19307 22400
rect 18708 22342 19307 22344
rect 18708 22340 18714 22342
rect 19241 22339 19307 22342
rect 26049 22402 26115 22405
rect 26200 22402 27000 22432
rect 26049 22400 27000 22402
rect 26049 22344 26054 22400
rect 26110 22344 27000 22400
rect 26049 22342 27000 22344
rect 26049 22339 26115 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 26200 22312 27000 22342
rect 22946 22271 23262 22272
rect 9121 22266 9187 22269
rect 12157 22266 12223 22269
rect 9121 22264 12223 22266
rect 9121 22208 9126 22264
rect 9182 22208 12162 22264
rect 12218 22208 12223 22264
rect 9121 22206 12223 22208
rect 9121 22203 9187 22206
rect 12157 22203 12223 22206
rect 16430 22204 16436 22268
rect 16500 22266 16506 22268
rect 20529 22266 20595 22269
rect 16500 22264 20595 22266
rect 16500 22208 20534 22264
rect 20590 22208 20595 22264
rect 16500 22206 20595 22208
rect 16500 22204 16506 22206
rect 20529 22203 20595 22206
rect 4153 22130 4219 22133
rect 16297 22130 16363 22133
rect 4153 22128 16363 22130
rect 4153 22072 4158 22128
rect 4214 22072 16302 22128
rect 16358 22072 16363 22128
rect 4153 22070 16363 22072
rect 4153 22067 4219 22070
rect 16297 22067 16363 22070
rect 16481 22130 16547 22133
rect 18229 22130 18295 22133
rect 16481 22128 18295 22130
rect 16481 22072 16486 22128
rect 16542 22072 18234 22128
rect 18290 22072 18295 22128
rect 16481 22070 18295 22072
rect 16481 22067 16547 22070
rect 18229 22067 18295 22070
rect 21950 22068 21956 22132
rect 22020 22130 22026 22132
rect 22461 22130 22527 22133
rect 22020 22128 22527 22130
rect 22020 22072 22466 22128
rect 22522 22072 22527 22128
rect 22020 22070 22527 22072
rect 22020 22068 22026 22070
rect 22461 22067 22527 22070
rect 3693 21994 3759 21997
rect 4245 21994 4311 21997
rect 4521 21994 4587 21997
rect 3693 21992 3802 21994
rect 3693 21936 3698 21992
rect 3754 21936 3802 21992
rect 3693 21931 3802 21936
rect 4245 21992 4587 21994
rect 4245 21936 4250 21992
rect 4306 21936 4526 21992
rect 4582 21936 4587 21992
rect 4245 21934 4587 21936
rect 4245 21931 4311 21934
rect 4521 21931 4587 21934
rect 6085 21994 6151 21997
rect 26200 21994 27000 22024
rect 6085 21992 18476 21994
rect 6085 21936 6090 21992
rect 6146 21936 18476 21992
rect 6085 21934 18476 21936
rect 6085 21931 6151 21934
rect 3742 21450 3802 21931
rect 5717 21858 5783 21861
rect 7005 21858 7071 21861
rect 5717 21856 7071 21858
rect 5717 21800 5722 21856
rect 5778 21800 7010 21856
rect 7066 21800 7071 21856
rect 5717 21798 7071 21800
rect 5717 21795 5783 21798
rect 7005 21795 7071 21798
rect 9806 21796 9812 21860
rect 9876 21858 9882 21860
rect 13629 21858 13695 21861
rect 9876 21856 13695 21858
rect 9876 21800 13634 21856
rect 13690 21800 13695 21856
rect 9876 21798 13695 21800
rect 18416 21858 18476 21934
rect 22050 21934 27000 21994
rect 20713 21858 20779 21861
rect 18416 21856 20779 21858
rect 18416 21800 20718 21856
rect 20774 21800 20779 21856
rect 18416 21798 20779 21800
rect 9876 21796 9882 21798
rect 13629 21795 13695 21798
rect 20713 21795 20779 21798
rect 21398 21796 21404 21860
rect 21468 21858 21474 21860
rect 22050 21858 22110 21934
rect 26200 21904 27000 21934
rect 21468 21798 22110 21858
rect 21468 21796 21474 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 11462 21660 11468 21724
rect 11532 21722 11538 21724
rect 14365 21722 14431 21725
rect 11532 21720 14431 21722
rect 11532 21664 14370 21720
rect 14426 21664 14431 21720
rect 11532 21662 14431 21664
rect 11532 21660 11538 21662
rect 14365 21659 14431 21662
rect 18454 21660 18460 21724
rect 18524 21722 18530 21724
rect 19609 21722 19675 21725
rect 18524 21720 19675 21722
rect 18524 21664 19614 21720
rect 19670 21664 19675 21720
rect 18524 21662 19675 21664
rect 18524 21660 18530 21662
rect 19609 21659 19675 21662
rect 8293 21586 8359 21589
rect 13486 21586 13492 21588
rect 8293 21584 13492 21586
rect 8293 21528 8298 21584
rect 8354 21528 13492 21584
rect 8293 21526 13492 21528
rect 8293 21523 8359 21526
rect 13486 21524 13492 21526
rect 13556 21586 13562 21588
rect 24393 21586 24459 21589
rect 26200 21586 27000 21616
rect 13556 21526 17786 21586
rect 13556 21524 13562 21526
rect 15561 21450 15627 21453
rect 17493 21452 17559 21453
rect 16062 21450 16068 21452
rect 3742 21448 16068 21450
rect 3742 21392 15566 21448
rect 15622 21392 16068 21448
rect 3742 21390 16068 21392
rect 3509 21314 3575 21317
rect 3742 21314 3802 21390
rect 15561 21387 15627 21390
rect 16062 21388 16068 21390
rect 16132 21388 16138 21452
rect 17493 21450 17540 21452
rect 17448 21448 17540 21450
rect 17448 21392 17498 21448
rect 17448 21390 17540 21392
rect 17493 21388 17540 21390
rect 17604 21388 17610 21452
rect 17726 21450 17786 21526
rect 24393 21584 27000 21586
rect 24393 21528 24398 21584
rect 24454 21528 27000 21584
rect 24393 21526 27000 21528
rect 24393 21523 24459 21526
rect 26200 21496 27000 21526
rect 24945 21450 25011 21453
rect 17726 21448 25011 21450
rect 17726 21392 24950 21448
rect 25006 21392 25011 21448
rect 17726 21390 25011 21392
rect 17493 21387 17559 21388
rect 24945 21387 25011 21390
rect 3509 21312 3802 21314
rect 3509 21256 3514 21312
rect 3570 21256 3802 21312
rect 3509 21254 3802 21256
rect 13629 21314 13695 21317
rect 20805 21314 20871 21317
rect 21449 21314 21515 21317
rect 13629 21312 21515 21314
rect 13629 21256 13634 21312
rect 13690 21256 20810 21312
rect 20866 21256 21454 21312
rect 21510 21256 21515 21312
rect 13629 21254 21515 21256
rect 3509 21251 3575 21254
rect 13629 21251 13695 21254
rect 20805 21251 20871 21254
rect 21449 21251 21515 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 4797 21178 4863 21181
rect 16481 21178 16547 21181
rect 20621 21178 20687 21181
rect 4797 21176 12450 21178
rect 4797 21120 4802 21176
rect 4858 21120 12450 21176
rect 4797 21118 12450 21120
rect 4797 21115 4863 21118
rect 9397 21042 9463 21045
rect 9622 21042 9628 21044
rect 9397 21040 9628 21042
rect 9397 20984 9402 21040
rect 9458 20984 9628 21040
rect 9397 20982 9628 20984
rect 9397 20979 9463 20982
rect 9622 20980 9628 20982
rect 9692 20980 9698 21044
rect 12390 21042 12450 21118
rect 16481 21176 20687 21178
rect 16481 21120 16486 21176
rect 16542 21120 20626 21176
rect 20682 21120 20687 21176
rect 16481 21118 20687 21120
rect 16481 21115 16547 21118
rect 20621 21115 20687 21118
rect 20805 21178 20871 21181
rect 21909 21178 21975 21181
rect 26200 21178 27000 21208
rect 20805 21176 21975 21178
rect 20805 21120 20810 21176
rect 20866 21120 21914 21176
rect 21970 21120 21975 21176
rect 20805 21118 21975 21120
rect 20805 21115 20871 21118
rect 21909 21115 21975 21118
rect 23614 21118 27000 21178
rect 23473 21042 23539 21045
rect 12390 21040 23539 21042
rect 12390 20984 23478 21040
rect 23534 20984 23539 21040
rect 12390 20982 23539 20984
rect 23473 20979 23539 20982
rect 7465 20906 7531 20909
rect 19701 20906 19767 20909
rect 7465 20904 19767 20906
rect 7465 20848 7470 20904
rect 7526 20848 19706 20904
rect 19762 20848 19767 20904
rect 7465 20846 19767 20848
rect 7465 20843 7531 20846
rect 19701 20843 19767 20846
rect 21633 20906 21699 20909
rect 22001 20906 22067 20909
rect 21633 20904 22067 20906
rect 21633 20848 21638 20904
rect 21694 20848 22006 20904
rect 22062 20848 22067 20904
rect 21633 20846 22067 20848
rect 21633 20843 21699 20846
rect 22001 20843 22067 20846
rect 22369 20906 22435 20909
rect 23614 20906 23674 21118
rect 26200 21088 27000 21118
rect 22369 20904 23674 20906
rect 22369 20848 22374 20904
rect 22430 20848 23674 20904
rect 22369 20846 23674 20848
rect 22369 20843 22435 20846
rect 3693 20770 3759 20773
rect 5758 20770 5764 20772
rect 3693 20768 5764 20770
rect 3693 20712 3698 20768
rect 3754 20712 5764 20768
rect 3693 20710 5764 20712
rect 3693 20707 3759 20710
rect 5758 20708 5764 20710
rect 5828 20708 5834 20772
rect 8661 20770 8727 20773
rect 16481 20770 16547 20773
rect 8661 20768 16547 20770
rect 8661 20712 8666 20768
rect 8722 20712 16486 20768
rect 16542 20712 16547 20768
rect 8661 20710 16547 20712
rect 8661 20707 8727 20710
rect 16481 20707 16547 20710
rect 16614 20708 16620 20772
rect 16684 20770 16690 20772
rect 17033 20770 17099 20773
rect 16684 20768 17099 20770
rect 16684 20712 17038 20768
rect 17094 20712 17099 20768
rect 16684 20710 17099 20712
rect 16684 20708 16690 20710
rect 17033 20707 17099 20710
rect 17166 20708 17172 20772
rect 17236 20770 17242 20772
rect 17769 20770 17835 20773
rect 19885 20772 19951 20773
rect 21173 20772 21239 20773
rect 19885 20770 19932 20772
rect 17236 20768 17835 20770
rect 17236 20712 17774 20768
rect 17830 20712 17835 20768
rect 17236 20710 17835 20712
rect 19840 20768 19932 20770
rect 19840 20712 19890 20768
rect 19840 20710 19932 20712
rect 17236 20708 17242 20710
rect 17769 20707 17835 20710
rect 19885 20708 19932 20710
rect 19996 20708 20002 20772
rect 21173 20770 21220 20772
rect 21128 20768 21220 20770
rect 21128 20712 21178 20768
rect 21128 20710 21220 20712
rect 21173 20708 21220 20710
rect 21284 20708 21290 20772
rect 21725 20770 21791 20773
rect 26200 20770 27000 20800
rect 21725 20768 27000 20770
rect 21725 20712 21730 20768
rect 21786 20712 27000 20768
rect 21725 20710 27000 20712
rect 19885 20707 19951 20708
rect 21173 20707 21239 20708
rect 21725 20707 21791 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 26200 20680 27000 20710
rect 17946 20639 18262 20640
rect 8385 20634 8451 20637
rect 9397 20634 9463 20637
rect 8385 20632 9463 20634
rect 8385 20576 8390 20632
rect 8446 20576 9402 20632
rect 9458 20576 9463 20632
rect 8385 20574 9463 20576
rect 8385 20571 8451 20574
rect 9397 20571 9463 20574
rect 12566 20572 12572 20636
rect 12636 20634 12642 20636
rect 15193 20634 15259 20637
rect 12636 20632 15259 20634
rect 12636 20576 15198 20632
rect 15254 20576 15259 20632
rect 12636 20574 15259 20576
rect 12636 20572 12642 20574
rect 15193 20571 15259 20574
rect 15326 20572 15332 20636
rect 15396 20634 15402 20636
rect 16297 20634 16363 20637
rect 15396 20632 16363 20634
rect 15396 20576 16302 20632
rect 16358 20576 16363 20632
rect 15396 20574 16363 20576
rect 15396 20572 15402 20574
rect 16297 20571 16363 20574
rect 22502 20572 22508 20636
rect 22572 20634 22578 20636
rect 22921 20634 22987 20637
rect 22572 20632 22987 20634
rect 22572 20576 22926 20632
rect 22982 20576 22987 20632
rect 22572 20574 22987 20576
rect 22572 20572 22578 20574
rect 22921 20571 22987 20574
rect 6821 20498 6887 20501
rect 18689 20498 18755 20501
rect 6821 20496 18755 20498
rect 6821 20440 6826 20496
rect 6882 20440 18694 20496
rect 18750 20440 18755 20496
rect 6821 20438 18755 20440
rect 6821 20435 6887 20438
rect 18689 20435 18755 20438
rect 7833 20362 7899 20365
rect 12525 20362 12591 20365
rect 13537 20362 13603 20365
rect 7833 20360 12591 20362
rect 7833 20304 7838 20360
rect 7894 20304 12530 20360
rect 12586 20304 12591 20360
rect 7833 20302 12591 20304
rect 7833 20299 7899 20302
rect 12525 20299 12591 20302
rect 12804 20360 13603 20362
rect 12804 20304 13542 20360
rect 13598 20304 13603 20360
rect 12804 20302 13603 20304
rect 7741 20226 7807 20229
rect 9305 20226 9371 20229
rect 7741 20224 9371 20226
rect 7741 20168 7746 20224
rect 7802 20168 9310 20224
rect 9366 20168 9371 20224
rect 7741 20166 9371 20168
rect 7741 20163 7807 20166
rect 9305 20163 9371 20166
rect 9581 20226 9647 20229
rect 12804 20226 12864 20302
rect 13537 20299 13603 20302
rect 14549 20362 14615 20365
rect 16573 20362 16639 20365
rect 14549 20360 16639 20362
rect 14549 20304 14554 20360
rect 14610 20304 16578 20360
rect 16634 20304 16639 20360
rect 14549 20302 16639 20304
rect 14549 20299 14615 20302
rect 16573 20299 16639 20302
rect 25957 20362 26023 20365
rect 26200 20362 27000 20392
rect 25957 20360 27000 20362
rect 25957 20304 25962 20360
rect 26018 20304 27000 20360
rect 25957 20302 27000 20304
rect 25957 20299 26023 20302
rect 26200 20272 27000 20302
rect 9581 20224 12864 20226
rect 9581 20168 9586 20224
rect 9642 20168 12864 20224
rect 9581 20166 12864 20168
rect 9581 20163 9647 20166
rect 15510 20164 15516 20228
rect 15580 20226 15586 20228
rect 15580 20166 16314 20226
rect 15580 20164 15586 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 7465 20090 7531 20093
rect 12065 20090 12131 20093
rect 7465 20088 12131 20090
rect 7465 20032 7470 20088
rect 7526 20032 12070 20088
rect 12126 20032 12131 20088
rect 7465 20030 12131 20032
rect 7465 20027 7531 20030
rect 12065 20027 12131 20030
rect 12525 20090 12591 20093
rect 12525 20088 12864 20090
rect 12525 20032 12530 20088
rect 12586 20032 12864 20088
rect 12525 20030 12864 20032
rect 12525 20027 12591 20030
rect 4889 19954 4955 19957
rect 8109 19954 8175 19957
rect 4889 19952 8175 19954
rect 4889 19896 4894 19952
rect 4950 19896 8114 19952
rect 8170 19896 8175 19952
rect 4889 19894 8175 19896
rect 4889 19891 4955 19894
rect 8109 19891 8175 19894
rect 8293 19954 8359 19957
rect 12566 19954 12572 19956
rect 8293 19952 12572 19954
rect 8293 19896 8298 19952
rect 8354 19896 12572 19952
rect 8293 19894 12572 19896
rect 8293 19891 8359 19894
rect 12566 19892 12572 19894
rect 12636 19892 12642 19956
rect 12804 19954 12864 20030
rect 15694 20028 15700 20092
rect 15764 20090 15770 20092
rect 16021 20090 16087 20093
rect 15764 20088 16087 20090
rect 15764 20032 16026 20088
rect 16082 20032 16087 20088
rect 15764 20030 16087 20032
rect 16254 20090 16314 20166
rect 16798 20164 16804 20228
rect 16868 20226 16874 20228
rect 22737 20226 22803 20229
rect 16868 20224 22803 20226
rect 16868 20168 22742 20224
rect 22798 20168 22803 20224
rect 16868 20166 22803 20168
rect 16868 20164 16874 20166
rect 22737 20163 22803 20166
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 16254 20030 22110 20090
rect 15764 20028 15770 20030
rect 16021 20027 16087 20030
rect 21449 19954 21515 19957
rect 12804 19952 21515 19954
rect 12804 19896 21454 19952
rect 21510 19896 21515 19952
rect 12804 19894 21515 19896
rect 22050 19954 22110 20030
rect 22185 19954 22251 19957
rect 24853 19954 24919 19957
rect 22050 19952 24919 19954
rect 22050 19896 22190 19952
rect 22246 19896 24858 19952
rect 24914 19896 24919 19952
rect 22050 19894 24919 19896
rect 21449 19891 21515 19894
rect 22185 19891 22251 19894
rect 24853 19891 24919 19894
rect 26049 19954 26115 19957
rect 26200 19954 27000 19984
rect 26049 19952 27000 19954
rect 26049 19896 26054 19952
rect 26110 19896 27000 19952
rect 26049 19894 27000 19896
rect 26049 19891 26115 19894
rect 26200 19864 27000 19894
rect 6545 19818 6611 19821
rect 25681 19818 25747 19821
rect 6545 19816 25747 19818
rect 6545 19760 6550 19816
rect 6606 19760 25686 19816
rect 25742 19760 25747 19816
rect 6545 19758 25747 19760
rect 6545 19755 6611 19758
rect 25681 19755 25747 19758
rect 8937 19682 9003 19685
rect 9305 19682 9371 19685
rect 8937 19680 9371 19682
rect 8937 19624 8942 19680
rect 8998 19624 9310 19680
rect 9366 19624 9371 19680
rect 8937 19622 9371 19624
rect 8937 19619 9003 19622
rect 9305 19619 9371 19622
rect 11513 19682 11579 19685
rect 14181 19682 14247 19685
rect 11513 19680 14247 19682
rect 11513 19624 11518 19680
rect 11574 19624 14186 19680
rect 14242 19624 14247 19680
rect 11513 19622 14247 19624
rect 11513 19619 11579 19622
rect 14181 19619 14247 19622
rect 20110 19620 20116 19684
rect 20180 19682 20186 19684
rect 20989 19682 21055 19685
rect 20180 19680 21055 19682
rect 20180 19624 20994 19680
rect 21050 19624 21055 19680
rect 20180 19622 21055 19624
rect 20180 19620 20186 19622
rect 20989 19619 21055 19622
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 4521 19546 4587 19549
rect 7281 19546 7347 19549
rect 15694 19546 15700 19548
rect 4521 19544 7347 19546
rect 4521 19488 4526 19544
rect 4582 19488 7286 19544
rect 7342 19488 7347 19544
rect 4521 19486 7347 19488
rect 4521 19483 4587 19486
rect 7281 19483 7347 19486
rect 12390 19486 15700 19546
rect 3877 19410 3943 19413
rect 12390 19410 12450 19486
rect 15694 19484 15700 19486
rect 15764 19484 15770 19548
rect 20662 19484 20668 19548
rect 20732 19546 20738 19548
rect 20897 19546 20963 19549
rect 20732 19544 20963 19546
rect 20732 19488 20902 19544
rect 20958 19488 20963 19544
rect 20732 19486 20963 19488
rect 20732 19484 20738 19486
rect 20897 19483 20963 19486
rect 24853 19546 24919 19549
rect 26200 19546 27000 19576
rect 24853 19544 27000 19546
rect 24853 19488 24858 19544
rect 24914 19488 27000 19544
rect 24853 19486 27000 19488
rect 24853 19483 24919 19486
rect 26200 19456 27000 19486
rect 3877 19408 12450 19410
rect 3877 19352 3882 19408
rect 3938 19352 12450 19408
rect 3877 19350 12450 19352
rect 13169 19410 13235 19413
rect 14365 19410 14431 19413
rect 13169 19408 14431 19410
rect 13169 19352 13174 19408
rect 13230 19352 14370 19408
rect 14426 19352 14431 19408
rect 13169 19350 14431 19352
rect 3877 19347 3943 19350
rect 13169 19347 13235 19350
rect 14365 19347 14431 19350
rect 14774 19348 14780 19412
rect 14844 19410 14850 19412
rect 18413 19410 18479 19413
rect 14844 19408 18479 19410
rect 14844 19352 18418 19408
rect 18474 19352 18479 19408
rect 14844 19350 18479 19352
rect 14844 19348 14850 19350
rect 18413 19347 18479 19350
rect 20846 19348 20852 19412
rect 20916 19410 20922 19412
rect 21817 19410 21883 19413
rect 20916 19408 21883 19410
rect 20916 19352 21822 19408
rect 21878 19352 21883 19408
rect 20916 19350 21883 19352
rect 20916 19348 20922 19350
rect 21817 19347 21883 19350
rect 22318 19348 22324 19412
rect 22388 19410 22394 19412
rect 22461 19410 22527 19413
rect 22388 19408 22527 19410
rect 22388 19352 22466 19408
rect 22522 19352 22527 19408
rect 22388 19350 22527 19352
rect 22388 19348 22394 19350
rect 22461 19347 22527 19350
rect 9397 19274 9463 19277
rect 9397 19272 20178 19274
rect 9397 19216 9402 19272
rect 9458 19216 20178 19272
rect 9397 19214 20178 19216
rect 9397 19211 9463 19214
rect 5441 19138 5507 19141
rect 10961 19138 11027 19141
rect 5441 19136 11027 19138
rect 5441 19080 5446 19136
rect 5502 19080 10966 19136
rect 11022 19080 11027 19136
rect 5441 19078 11027 19080
rect 5441 19075 5507 19078
rect 10961 19075 11027 19078
rect 13537 19138 13603 19141
rect 16573 19138 16639 19141
rect 13537 19136 16639 19138
rect 13537 19080 13542 19136
rect 13598 19080 16578 19136
rect 16634 19080 16639 19136
rect 13537 19078 16639 19080
rect 13537 19075 13603 19078
rect 16573 19075 16639 19078
rect 18454 19076 18460 19140
rect 18524 19138 18530 19140
rect 19333 19138 19399 19141
rect 18524 19136 19399 19138
rect 18524 19080 19338 19136
rect 19394 19080 19399 19136
rect 18524 19078 19399 19080
rect 20118 19138 20178 19214
rect 20294 19212 20300 19276
rect 20364 19274 20370 19276
rect 23381 19274 23447 19277
rect 20364 19272 23447 19274
rect 20364 19216 23386 19272
rect 23442 19216 23447 19272
rect 20364 19214 23447 19216
rect 20364 19212 20370 19214
rect 23381 19211 23447 19214
rect 20345 19138 20411 19141
rect 20118 19136 20411 19138
rect 20118 19080 20350 19136
rect 20406 19080 20411 19136
rect 20118 19078 20411 19080
rect 18524 19076 18530 19078
rect 19333 19075 19399 19078
rect 20345 19075 20411 19078
rect 23381 19138 23447 19141
rect 26200 19138 27000 19168
rect 23381 19136 27000 19138
rect 23381 19080 23386 19136
rect 23442 19080 27000 19136
rect 23381 19078 27000 19080
rect 23381 19075 23447 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 26200 19048 27000 19078
rect 22946 19007 23262 19008
rect 10910 18940 10916 19004
rect 10980 19002 10986 19004
rect 11421 19002 11487 19005
rect 10980 19000 11487 19002
rect 10980 18944 11426 19000
rect 11482 18944 11487 19000
rect 10980 18942 11487 18944
rect 10980 18940 10986 18942
rect 11421 18939 11487 18942
rect 14365 19002 14431 19005
rect 17861 19002 17927 19005
rect 14365 19000 17927 19002
rect 14365 18944 14370 19000
rect 14426 18944 17866 19000
rect 17922 18944 17927 19000
rect 14365 18942 17927 18944
rect 14365 18939 14431 18942
rect 17861 18939 17927 18942
rect 18822 18940 18828 19004
rect 18892 19002 18898 19004
rect 21081 19002 21147 19005
rect 18892 19000 21147 19002
rect 18892 18944 21086 19000
rect 21142 18944 21147 19000
rect 18892 18942 21147 18944
rect 18892 18940 18898 18942
rect 21081 18939 21147 18942
rect 24669 19002 24735 19005
rect 24669 19000 25330 19002
rect 24669 18944 24674 19000
rect 24730 18944 25330 19000
rect 24669 18942 25330 18944
rect 24669 18939 24735 18942
rect 2129 18866 2195 18869
rect 2129 18864 25146 18866
rect 2129 18808 2134 18864
rect 2190 18808 25146 18864
rect 2129 18806 25146 18808
rect 2129 18803 2195 18806
rect 5257 18730 5323 18733
rect 9254 18730 9260 18732
rect 5257 18728 9260 18730
rect 5257 18672 5262 18728
rect 5318 18672 9260 18728
rect 5257 18670 9260 18672
rect 5257 18667 5323 18670
rect 9254 18668 9260 18670
rect 9324 18668 9330 18732
rect 11421 18730 11487 18733
rect 19333 18730 19399 18733
rect 11421 18728 19399 18730
rect 11421 18672 11426 18728
rect 11482 18672 19338 18728
rect 19394 18672 19399 18728
rect 11421 18670 19399 18672
rect 11421 18667 11487 18670
rect 19333 18667 19399 18670
rect 23422 18668 23428 18732
rect 23492 18730 23498 18732
rect 23657 18730 23723 18733
rect 23492 18728 23723 18730
rect 23492 18672 23662 18728
rect 23718 18672 23723 18728
rect 23492 18670 23723 18672
rect 23492 18668 23498 18670
rect 23657 18667 23723 18670
rect 11094 18532 11100 18596
rect 11164 18594 11170 18596
rect 15142 18594 15148 18596
rect 11164 18534 15148 18594
rect 11164 18532 11170 18534
rect 15142 18532 15148 18534
rect 15212 18532 15218 18596
rect 22134 18532 22140 18596
rect 22204 18594 22210 18596
rect 23013 18594 23079 18597
rect 22204 18592 23079 18594
rect 22204 18536 23018 18592
rect 23074 18536 23079 18592
rect 22204 18534 23079 18536
rect 22204 18532 22210 18534
rect 23013 18531 23079 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 7649 18458 7715 18461
rect 7782 18458 7788 18460
rect 7649 18456 7788 18458
rect 7649 18400 7654 18456
rect 7710 18400 7788 18456
rect 7649 18398 7788 18400
rect 7649 18395 7715 18398
rect 7782 18396 7788 18398
rect 7852 18396 7858 18460
rect 8385 18458 8451 18461
rect 9029 18458 9095 18461
rect 8385 18456 17234 18458
rect 8385 18400 8390 18456
rect 8446 18400 9034 18456
rect 9090 18400 17234 18456
rect 8385 18398 17234 18400
rect 8385 18395 8451 18398
rect 9029 18395 9095 18398
rect 4337 18322 4403 18325
rect 5165 18322 5231 18325
rect 16481 18322 16547 18325
rect 4337 18320 16547 18322
rect 4337 18264 4342 18320
rect 4398 18264 5170 18320
rect 5226 18264 16486 18320
rect 16542 18264 16547 18320
rect 4337 18262 16547 18264
rect 17174 18322 17234 18398
rect 24945 18322 25011 18325
rect 17174 18320 25011 18322
rect 17174 18264 24950 18320
rect 25006 18264 25011 18320
rect 17174 18262 25011 18264
rect 25086 18322 25146 18806
rect 25270 18730 25330 18942
rect 26200 18730 27000 18760
rect 25270 18670 27000 18730
rect 26200 18640 27000 18670
rect 26200 18322 27000 18352
rect 25086 18262 27000 18322
rect 4337 18259 4403 18262
rect 5165 18259 5231 18262
rect 16481 18259 16547 18262
rect 24945 18259 25011 18262
rect 26200 18232 27000 18262
rect 8201 18186 8267 18189
rect 17217 18186 17283 18189
rect 8201 18184 17283 18186
rect 8201 18128 8206 18184
rect 8262 18128 17222 18184
rect 17278 18128 17283 18184
rect 8201 18126 17283 18128
rect 8201 18123 8267 18126
rect 17217 18123 17283 18126
rect 3366 17988 3372 18052
rect 3436 18050 3442 18052
rect 5942 18050 5948 18052
rect 3436 17990 5948 18050
rect 3436 17988 3442 17990
rect 5942 17988 5948 17990
rect 6012 17988 6018 18052
rect 7465 18050 7531 18053
rect 7598 18050 7604 18052
rect 7465 18048 7604 18050
rect 7465 17992 7470 18048
rect 7526 17992 7604 18048
rect 7465 17990 7604 17992
rect 7465 17987 7531 17990
rect 7598 17988 7604 17990
rect 7668 17988 7674 18052
rect 8293 18050 8359 18053
rect 11462 18050 11468 18052
rect 8293 18048 11468 18050
rect 8293 17992 8298 18048
rect 8354 17992 11468 18048
rect 8293 17990 11468 17992
rect 8293 17987 8359 17990
rect 11462 17988 11468 17990
rect 11532 17988 11538 18052
rect 15009 18050 15075 18053
rect 16757 18050 16823 18053
rect 15009 18048 16823 18050
rect 15009 17992 15014 18048
rect 15070 17992 16762 18048
rect 16818 17992 16823 18048
rect 15009 17990 16823 17992
rect 15009 17987 15075 17990
rect 16757 17987 16823 17990
rect 23606 17988 23612 18052
rect 23676 18050 23682 18052
rect 24577 18050 24643 18053
rect 23676 18048 24643 18050
rect 23676 17992 24582 18048
rect 24638 17992 24643 18048
rect 23676 17990 24643 17992
rect 23676 17988 23682 17990
rect 24577 17987 24643 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 8293 17914 8359 17917
rect 8518 17914 8524 17916
rect 8293 17912 8524 17914
rect 8293 17856 8298 17912
rect 8354 17856 8524 17912
rect 8293 17854 8524 17856
rect 8293 17851 8359 17854
rect 8518 17852 8524 17854
rect 8588 17852 8594 17916
rect 17401 17914 17467 17917
rect 14046 17912 17467 17914
rect 14046 17856 17406 17912
rect 17462 17856 17467 17912
rect 14046 17854 17467 17856
rect 7557 17778 7623 17781
rect 14046 17778 14106 17854
rect 17401 17851 17467 17854
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 7557 17776 14106 17778
rect 7557 17720 7562 17776
rect 7618 17720 14106 17776
rect 7557 17718 14106 17720
rect 14273 17778 14339 17781
rect 22921 17778 22987 17781
rect 14273 17776 22987 17778
rect 14273 17720 14278 17776
rect 14334 17720 22926 17776
rect 22982 17720 22987 17776
rect 14273 17718 22987 17720
rect 7557 17715 7623 17718
rect 14273 17715 14339 17718
rect 22921 17715 22987 17718
rect 6177 17642 6243 17645
rect 20253 17642 20319 17645
rect 22921 17642 22987 17645
rect 6177 17640 18476 17642
rect 6177 17584 6182 17640
rect 6238 17584 18476 17640
rect 6177 17582 18476 17584
rect 6177 17579 6243 17582
rect 8477 17506 8543 17509
rect 16849 17506 16915 17509
rect 8477 17504 16915 17506
rect 8477 17448 8482 17504
rect 8538 17448 16854 17504
rect 16910 17448 16915 17504
rect 8477 17446 16915 17448
rect 18416 17506 18476 17582
rect 20253 17640 22987 17642
rect 20253 17584 20258 17640
rect 20314 17584 22926 17640
rect 22982 17584 22987 17640
rect 20253 17582 22987 17584
rect 20253 17579 20319 17582
rect 22921 17579 22987 17582
rect 26200 17506 27000 17536
rect 18416 17446 27000 17506
rect 8477 17443 8543 17446
rect 16849 17443 16915 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 26200 17416 27000 17446
rect 17946 17375 18262 17376
rect 8661 17370 8727 17373
rect 15837 17370 15903 17373
rect 8661 17368 15903 17370
rect 8661 17312 8666 17368
rect 8722 17312 15842 17368
rect 15898 17312 15903 17368
rect 8661 17310 15903 17312
rect 8661 17307 8727 17310
rect 15837 17307 15903 17310
rect 23197 17370 23263 17373
rect 25773 17370 25839 17373
rect 23197 17368 25839 17370
rect 23197 17312 23202 17368
rect 23258 17312 25778 17368
rect 25834 17312 25839 17368
rect 23197 17310 25839 17312
rect 23197 17307 23263 17310
rect 25773 17307 25839 17310
rect 6913 17234 6979 17237
rect 10317 17234 10383 17237
rect 6913 17232 10383 17234
rect 6913 17176 6918 17232
rect 6974 17176 10322 17232
rect 10378 17176 10383 17232
rect 6913 17174 10383 17176
rect 6913 17171 6979 17174
rect 10317 17171 10383 17174
rect 11053 17234 11119 17237
rect 14733 17234 14799 17237
rect 11053 17232 14799 17234
rect 11053 17176 11058 17232
rect 11114 17176 14738 17232
rect 14794 17176 14799 17232
rect 11053 17174 14799 17176
rect 11053 17171 11119 17174
rect 14733 17171 14799 17174
rect 15469 17234 15535 17237
rect 15469 17232 16682 17234
rect 15469 17176 15474 17232
rect 15530 17176 16682 17232
rect 15469 17174 16682 17176
rect 15469 17171 15535 17174
rect 2773 17098 2839 17101
rect 5901 17098 5967 17101
rect 16481 17098 16547 17101
rect 2773 17096 3434 17098
rect 2773 17040 2778 17096
rect 2834 17040 3434 17096
rect 2773 17038 3434 17040
rect 2773 17035 2839 17038
rect 3374 16962 3434 17038
rect 5901 17096 16547 17098
rect 5901 17040 5906 17096
rect 5962 17040 16486 17096
rect 16542 17040 16547 17096
rect 5901 17038 16547 17040
rect 16622 17098 16682 17174
rect 16982 17172 16988 17236
rect 17052 17234 17058 17236
rect 22318 17234 22324 17236
rect 17052 17174 22324 17234
rect 17052 17172 17058 17174
rect 22318 17172 22324 17174
rect 22388 17172 22394 17236
rect 18965 17098 19031 17101
rect 16622 17096 19031 17098
rect 16622 17040 18970 17096
rect 19026 17040 19031 17096
rect 16622 17038 19031 17040
rect 5901 17035 5967 17038
rect 16481 17035 16547 17038
rect 18965 17035 19031 17038
rect 22093 17098 22159 17101
rect 26200 17098 27000 17128
rect 22093 17096 27000 17098
rect 22093 17040 22098 17096
rect 22154 17040 27000 17096
rect 22093 17038 27000 17040
rect 22093 17035 22159 17038
rect 26200 17008 27000 17038
rect 11646 16962 11652 16964
rect 3374 16902 11652 16962
rect 11646 16900 11652 16902
rect 11716 16900 11722 16964
rect 14733 16962 14799 16965
rect 22645 16962 22711 16965
rect 14733 16960 22711 16962
rect 14733 16904 14738 16960
rect 14794 16904 22650 16960
rect 22706 16904 22711 16960
rect 14733 16902 22711 16904
rect 14733 16899 14799 16902
rect 22645 16899 22711 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 9673 16826 9739 16829
rect 11513 16828 11579 16829
rect 10174 16826 10180 16828
rect 9673 16824 10180 16826
rect 9673 16768 9678 16824
rect 9734 16768 10180 16824
rect 9673 16766 10180 16768
rect 9673 16763 9739 16766
rect 10174 16764 10180 16766
rect 10244 16764 10250 16828
rect 11462 16826 11468 16828
rect 11422 16766 11468 16826
rect 11532 16824 11579 16828
rect 11574 16768 11579 16824
rect 11462 16764 11468 16766
rect 11532 16764 11579 16768
rect 11513 16763 11579 16764
rect 13353 16826 13419 16829
rect 15653 16826 15719 16829
rect 15878 16826 15884 16828
rect 13353 16824 14796 16826
rect 13353 16768 13358 16824
rect 13414 16768 14796 16824
rect 13353 16766 14796 16768
rect 13353 16763 13419 16766
rect 5625 16690 5691 16693
rect 12525 16690 12591 16693
rect 14549 16690 14615 16693
rect 5625 16688 14615 16690
rect 5625 16632 5630 16688
rect 5686 16632 12530 16688
rect 12586 16632 14554 16688
rect 14610 16632 14615 16688
rect 5625 16630 14615 16632
rect 14736 16690 14796 16766
rect 15653 16824 15884 16826
rect 15653 16768 15658 16824
rect 15714 16768 15884 16824
rect 15653 16766 15884 16768
rect 15653 16763 15719 16766
rect 15878 16764 15884 16766
rect 15948 16764 15954 16828
rect 23381 16826 23447 16829
rect 23381 16824 25330 16826
rect 23381 16768 23386 16824
rect 23442 16768 25330 16824
rect 23381 16766 25330 16768
rect 23381 16763 23447 16766
rect 18689 16690 18755 16693
rect 14736 16688 18755 16690
rect 14736 16632 18694 16688
rect 18750 16632 18755 16688
rect 14736 16630 18755 16632
rect 5625 16627 5691 16630
rect 12525 16627 12591 16630
rect 14549 16627 14615 16630
rect 18689 16627 18755 16630
rect 22686 16628 22692 16692
rect 22756 16690 22762 16692
rect 23289 16690 23355 16693
rect 22756 16688 23355 16690
rect 22756 16632 23294 16688
rect 23350 16632 23355 16688
rect 22756 16630 23355 16632
rect 22756 16628 22762 16630
rect 23289 16627 23355 16630
rect 24526 16628 24532 16692
rect 24596 16690 24602 16692
rect 25037 16690 25103 16693
rect 24596 16688 25103 16690
rect 24596 16632 25042 16688
rect 25098 16632 25103 16688
rect 24596 16630 25103 16632
rect 25270 16690 25330 16766
rect 26200 16690 27000 16720
rect 25270 16630 27000 16690
rect 24596 16628 24602 16630
rect 25037 16627 25103 16630
rect 26200 16600 27000 16630
rect 2037 16554 2103 16557
rect 8661 16554 8727 16557
rect 15561 16554 15627 16557
rect 2037 16552 8402 16554
rect 2037 16496 2042 16552
rect 2098 16496 8402 16552
rect 2037 16494 8402 16496
rect 2037 16491 2103 16494
rect 8342 16418 8402 16494
rect 8661 16552 15627 16554
rect 8661 16496 8666 16552
rect 8722 16496 15566 16552
rect 15622 16496 15627 16552
rect 8661 16494 15627 16496
rect 8661 16491 8727 16494
rect 15561 16491 15627 16494
rect 22645 16554 22711 16557
rect 24117 16554 24183 16557
rect 22645 16552 24183 16554
rect 22645 16496 22650 16552
rect 22706 16496 24122 16552
rect 24178 16496 24183 16552
rect 22645 16494 24183 16496
rect 22645 16491 22711 16494
rect 24117 16491 24183 16494
rect 16430 16418 16436 16420
rect 8342 16358 16436 16418
rect 16430 16356 16436 16358
rect 16500 16356 16506 16420
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 6361 16282 6427 16285
rect 6494 16282 6500 16284
rect 6361 16280 6500 16282
rect 6361 16224 6366 16280
rect 6422 16224 6500 16280
rect 6361 16222 6500 16224
rect 6361 16219 6427 16222
rect 6494 16220 6500 16222
rect 6564 16220 6570 16284
rect 11145 16282 11211 16285
rect 26200 16282 27000 16312
rect 11145 16280 17234 16282
rect 11145 16224 11150 16280
rect 11206 16224 17234 16280
rect 11145 16222 17234 16224
rect 11145 16219 11211 16222
rect 1853 16146 1919 16149
rect 16982 16146 16988 16148
rect 1853 16144 16988 16146
rect 1853 16088 1858 16144
rect 1914 16088 16988 16144
rect 1853 16086 16988 16088
rect 1853 16083 1919 16086
rect 16982 16084 16988 16086
rect 17052 16084 17058 16148
rect 17174 16146 17234 16222
rect 22050 16222 27000 16282
rect 22050 16146 22110 16222
rect 26200 16192 27000 16222
rect 17174 16086 22110 16146
rect 9121 16010 9187 16013
rect 15101 16010 15167 16013
rect 9121 16008 15167 16010
rect 9121 15952 9126 16008
rect 9182 15952 15106 16008
rect 15162 15952 15167 16008
rect 9121 15950 15167 15952
rect 9121 15947 9187 15950
rect 15101 15947 15167 15950
rect 15561 16010 15627 16013
rect 21541 16010 21607 16013
rect 15561 16008 21607 16010
rect 15561 15952 15566 16008
rect 15622 15952 21546 16008
rect 21602 15952 21607 16008
rect 15561 15950 21607 15952
rect 15561 15947 15627 15950
rect 21541 15947 21607 15950
rect 5441 15874 5507 15877
rect 10910 15874 10916 15876
rect 5441 15872 10916 15874
rect 5441 15816 5446 15872
rect 5502 15816 10916 15872
rect 5441 15814 10916 15816
rect 5441 15811 5507 15814
rect 10910 15812 10916 15814
rect 10980 15812 10986 15876
rect 13721 15874 13787 15877
rect 18505 15874 18571 15877
rect 26200 15874 27000 15904
rect 13721 15872 18571 15874
rect 13721 15816 13726 15872
rect 13782 15816 18510 15872
rect 18566 15816 18571 15872
rect 13721 15814 18571 15816
rect 13721 15811 13787 15814
rect 18505 15811 18571 15814
rect 24166 15814 27000 15874
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 4889 15738 4955 15741
rect 11789 15738 11855 15741
rect 4889 15736 11855 15738
rect 4889 15680 4894 15736
rect 4950 15680 11794 15736
rect 11850 15680 11855 15736
rect 4889 15678 11855 15680
rect 4889 15675 4955 15678
rect 11789 15675 11855 15678
rect 17033 15738 17099 15741
rect 18822 15738 18828 15740
rect 17033 15736 18828 15738
rect 17033 15680 17038 15736
rect 17094 15680 18828 15736
rect 17033 15678 18828 15680
rect 17033 15675 17099 15678
rect 18822 15676 18828 15678
rect 18892 15676 18898 15740
rect 5390 15540 5396 15604
rect 5460 15602 5466 15604
rect 7189 15602 7255 15605
rect 5460 15600 7255 15602
rect 5460 15544 7194 15600
rect 7250 15544 7255 15600
rect 5460 15542 7255 15544
rect 5460 15540 5466 15542
rect 7189 15539 7255 15542
rect 8201 15602 8267 15605
rect 19333 15602 19399 15605
rect 8201 15600 19399 15602
rect 8201 15544 8206 15600
rect 8262 15544 19338 15600
rect 19394 15544 19399 15600
rect 8201 15542 19399 15544
rect 8201 15539 8267 15542
rect 19333 15539 19399 15542
rect 21398 15540 21404 15604
rect 21468 15602 21474 15604
rect 24166 15602 24226 15814
rect 26200 15784 27000 15814
rect 21468 15542 24226 15602
rect 21468 15540 21474 15542
rect 9765 15466 9831 15469
rect 17033 15466 17099 15469
rect 18873 15466 18939 15469
rect 9765 15464 17099 15466
rect 9765 15408 9770 15464
rect 9826 15408 17038 15464
rect 17094 15408 17099 15464
rect 9765 15406 17099 15408
rect 9765 15403 9831 15406
rect 17033 15403 17099 15406
rect 17772 15464 18939 15466
rect 17772 15408 18878 15464
rect 18934 15408 18939 15464
rect 17772 15406 18939 15408
rect 11237 15330 11303 15333
rect 17772 15330 17832 15406
rect 18873 15403 18939 15406
rect 19977 15466 20043 15469
rect 22134 15466 22140 15468
rect 19977 15464 22140 15466
rect 19977 15408 19982 15464
rect 20038 15408 22140 15464
rect 19977 15406 22140 15408
rect 19977 15403 20043 15406
rect 22134 15404 22140 15406
rect 22204 15404 22210 15468
rect 23841 15466 23907 15469
rect 26200 15466 27000 15496
rect 23841 15464 27000 15466
rect 23841 15408 23846 15464
rect 23902 15408 27000 15464
rect 23841 15406 27000 15408
rect 23841 15403 23907 15406
rect 26200 15376 27000 15406
rect 11237 15328 17832 15330
rect 11237 15272 11242 15328
rect 11298 15272 17832 15328
rect 11237 15270 17832 15272
rect 11237 15267 11303 15270
rect 19190 15268 19196 15332
rect 19260 15330 19266 15332
rect 20621 15330 20687 15333
rect 23381 15330 23447 15333
rect 19260 15328 20687 15330
rect 19260 15272 20626 15328
rect 20682 15272 20687 15328
rect 19260 15270 20687 15272
rect 19260 15268 19266 15270
rect 20621 15267 20687 15270
rect 20854 15328 23447 15330
rect 20854 15272 23386 15328
rect 23442 15272 23447 15328
rect 20854 15270 23447 15272
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 3785 15194 3851 15197
rect 4654 15194 4660 15196
rect 3785 15192 4660 15194
rect 3785 15136 3790 15192
rect 3846 15136 4660 15192
rect 3785 15134 4660 15136
rect 3785 15131 3851 15134
rect 4654 15132 4660 15134
rect 4724 15132 4730 15196
rect 8385 15194 8451 15197
rect 14038 15194 14044 15196
rect 8385 15192 14044 15194
rect 8385 15136 8390 15192
rect 8446 15136 14044 15192
rect 8385 15134 14044 15136
rect 8385 15131 8451 15134
rect 14038 15132 14044 15134
rect 14108 15132 14114 15196
rect 20529 15194 20595 15197
rect 20854 15194 20914 15270
rect 23381 15267 23447 15270
rect 22093 15194 22159 15197
rect 23473 15194 23539 15197
rect 20529 15192 20914 15194
rect 20529 15136 20534 15192
rect 20590 15136 20914 15192
rect 20529 15134 20914 15136
rect 22050 15192 23539 15194
rect 22050 15136 22098 15192
rect 22154 15136 23478 15192
rect 23534 15136 23539 15192
rect 22050 15134 23539 15136
rect 20529 15131 20595 15134
rect 22050 15131 22159 15134
rect 23473 15131 23539 15134
rect 2773 15058 2839 15061
rect 3366 15058 3372 15060
rect 2773 15056 3372 15058
rect 2773 15000 2778 15056
rect 2834 15000 3372 15056
rect 2773 14998 3372 15000
rect 2773 14995 2839 14998
rect 3366 14996 3372 14998
rect 3436 14996 3442 15060
rect 6729 15058 6795 15061
rect 22050 15058 22110 15131
rect 6729 15056 22110 15058
rect 6729 15000 6734 15056
rect 6790 15000 22110 15056
rect 6729 14998 22110 15000
rect 22553 15058 22619 15061
rect 26200 15058 27000 15088
rect 22553 15056 27000 15058
rect 22553 15000 22558 15056
rect 22614 15000 27000 15056
rect 22553 14998 27000 15000
rect 6729 14995 6795 14998
rect 22553 14995 22619 14998
rect 26200 14968 27000 14998
rect 8753 14922 8819 14925
rect 18454 14922 18460 14924
rect 8753 14920 18460 14922
rect 8753 14864 8758 14920
rect 8814 14864 18460 14920
rect 8753 14862 18460 14864
rect 8753 14859 8819 14862
rect 18454 14860 18460 14862
rect 18524 14860 18530 14924
rect 19006 14860 19012 14924
rect 19076 14922 19082 14924
rect 21950 14922 21956 14924
rect 19076 14862 21956 14922
rect 19076 14860 19082 14862
rect 21950 14860 21956 14862
rect 22020 14860 22026 14924
rect 4337 14786 4403 14789
rect 9990 14786 9996 14788
rect 4337 14784 9996 14786
rect 4337 14728 4342 14784
rect 4398 14728 9996 14784
rect 4337 14726 9996 14728
rect 4337 14723 4403 14726
rect 9990 14724 9996 14726
rect 10060 14724 10066 14788
rect 15142 14724 15148 14788
rect 15212 14786 15218 14788
rect 22185 14786 22251 14789
rect 15212 14784 22251 14786
rect 15212 14728 22190 14784
rect 22246 14728 22251 14784
rect 15212 14726 22251 14728
rect 15212 14724 15218 14726
rect 22185 14723 22251 14726
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 14641 14650 14707 14653
rect 22502 14650 22508 14652
rect 14641 14648 22508 14650
rect 14641 14592 14646 14648
rect 14702 14592 22508 14648
rect 14641 14590 22508 14592
rect 14641 14587 14707 14590
rect 22502 14588 22508 14590
rect 22572 14588 22578 14652
rect 23381 14650 23447 14653
rect 26200 14650 27000 14680
rect 23381 14648 27000 14650
rect 23381 14592 23386 14648
rect 23442 14592 27000 14648
rect 23381 14590 27000 14592
rect 23381 14587 23447 14590
rect 26200 14560 27000 14590
rect 2313 14514 2379 14517
rect 5533 14516 5599 14517
rect 2630 14514 2636 14516
rect 2313 14512 2636 14514
rect 2313 14456 2318 14512
rect 2374 14456 2636 14512
rect 2313 14454 2636 14456
rect 2313 14451 2379 14454
rect 2630 14452 2636 14454
rect 2700 14452 2706 14516
rect 5533 14514 5580 14516
rect 5488 14512 5580 14514
rect 5488 14456 5538 14512
rect 5488 14454 5580 14456
rect 5533 14452 5580 14454
rect 5644 14452 5650 14516
rect 9622 14452 9628 14516
rect 9692 14514 9698 14516
rect 9692 14454 15210 14514
rect 9692 14452 9698 14454
rect 5533 14451 5599 14452
rect 15150 14381 15210 14454
rect 7281 14378 7347 14381
rect 14549 14378 14615 14381
rect 15009 14378 15075 14381
rect 7281 14376 12450 14378
rect 7281 14320 7286 14376
rect 7342 14320 12450 14376
rect 7281 14318 12450 14320
rect 7281 14315 7347 14318
rect 10133 14242 10199 14245
rect 11094 14242 11100 14244
rect 10133 14240 11100 14242
rect 10133 14184 10138 14240
rect 10194 14184 11100 14240
rect 10133 14182 11100 14184
rect 10133 14179 10199 14182
rect 11094 14180 11100 14182
rect 11164 14180 11170 14244
rect 12390 14242 12450 14318
rect 14549 14376 15075 14378
rect 14549 14320 14554 14376
rect 14610 14320 15014 14376
rect 15070 14320 15075 14376
rect 14549 14318 15075 14320
rect 15150 14378 15259 14381
rect 23289 14378 23355 14381
rect 15150 14376 23355 14378
rect 15150 14320 15198 14376
rect 15254 14320 23294 14376
rect 23350 14320 23355 14376
rect 15150 14318 23355 14320
rect 14549 14315 14615 14318
rect 15009 14315 15075 14318
rect 15193 14315 15259 14318
rect 23289 14315 23355 14318
rect 16389 14242 16455 14245
rect 12390 14240 16455 14242
rect 12390 14184 16394 14240
rect 16450 14184 16455 14240
rect 12390 14182 16455 14184
rect 16389 14179 16455 14182
rect 23381 14242 23447 14245
rect 26200 14242 27000 14272
rect 23381 14240 27000 14242
rect 23381 14184 23386 14240
rect 23442 14184 27000 14240
rect 23381 14182 27000 14184
rect 23381 14179 23447 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 15653 14106 15719 14109
rect 22553 14106 22619 14109
rect 9216 14104 15719 14106
rect 9216 14048 15658 14104
rect 15714 14048 15719 14104
rect 9216 14046 15719 14048
rect 2313 13970 2379 13973
rect 7833 13970 7899 13973
rect 9216 13970 9276 14046
rect 15653 14043 15719 14046
rect 22142 14104 22619 14106
rect 22142 14048 22558 14104
rect 22614 14048 22619 14104
rect 22142 14046 22619 14048
rect 2313 13968 2790 13970
rect 2313 13912 2318 13968
rect 2374 13912 2790 13968
rect 2313 13910 2790 13912
rect 2313 13907 2379 13910
rect 2730 13834 2790 13910
rect 7833 13968 9276 13970
rect 7833 13912 7838 13968
rect 7894 13912 9276 13968
rect 7833 13910 9276 13912
rect 9673 13970 9739 13973
rect 19977 13970 20043 13973
rect 9673 13968 20043 13970
rect 9673 13912 9678 13968
rect 9734 13912 19982 13968
rect 20038 13912 20043 13968
rect 9673 13910 20043 13912
rect 7833 13907 7899 13910
rect 9673 13907 9739 13910
rect 19977 13907 20043 13910
rect 7925 13834 7991 13837
rect 2730 13832 7991 13834
rect 2730 13776 7930 13832
rect 7986 13776 7991 13832
rect 2730 13774 7991 13776
rect 7925 13771 7991 13774
rect 9673 13834 9739 13837
rect 9806 13834 9812 13836
rect 9673 13832 9812 13834
rect 9673 13776 9678 13832
rect 9734 13776 9812 13832
rect 9673 13774 9812 13776
rect 9673 13771 9739 13774
rect 9806 13772 9812 13774
rect 9876 13772 9882 13836
rect 13486 13772 13492 13836
rect 13556 13834 13562 13836
rect 13629 13834 13695 13837
rect 13556 13832 13695 13834
rect 13556 13776 13634 13832
rect 13690 13776 13695 13832
rect 13556 13774 13695 13776
rect 13556 13772 13562 13774
rect 13629 13771 13695 13774
rect 15285 13834 15351 13837
rect 16941 13834 17007 13837
rect 15285 13832 17007 13834
rect 15285 13776 15290 13832
rect 15346 13776 16946 13832
rect 17002 13776 17007 13832
rect 15285 13774 17007 13776
rect 15285 13771 15351 13774
rect 16941 13771 17007 13774
rect 19793 13834 19859 13837
rect 21081 13834 21147 13837
rect 19793 13832 21147 13834
rect 19793 13776 19798 13832
rect 19854 13776 21086 13832
rect 21142 13776 21147 13832
rect 19793 13774 21147 13776
rect 19793 13771 19859 13774
rect 21081 13771 21147 13774
rect 22142 13701 22202 14046
rect 22553 14043 22619 14046
rect 22318 13908 22324 13972
rect 22388 13970 22394 13972
rect 22921 13970 22987 13973
rect 22388 13968 22987 13970
rect 22388 13912 22926 13968
rect 22982 13912 22987 13968
rect 22388 13910 22987 13912
rect 22388 13908 22394 13910
rect 22921 13907 22987 13910
rect 24710 13908 24716 13972
rect 24780 13970 24786 13972
rect 24945 13970 25011 13973
rect 24780 13968 25011 13970
rect 24780 13912 24950 13968
rect 25006 13912 25011 13968
rect 24780 13910 25011 13912
rect 24780 13908 24786 13910
rect 24945 13907 25011 13910
rect 22553 13834 22619 13837
rect 26200 13834 27000 13864
rect 22553 13832 27000 13834
rect 22553 13776 22558 13832
rect 22614 13776 27000 13832
rect 22553 13774 27000 13776
rect 22553 13771 22619 13774
rect 26200 13744 27000 13774
rect 22093 13696 22202 13701
rect 22093 13640 22098 13696
rect 22154 13640 22202 13696
rect 22093 13638 22202 13640
rect 25405 13698 25471 13701
rect 25681 13698 25747 13701
rect 25405 13696 25747 13698
rect 25405 13640 25410 13696
rect 25466 13640 25686 13696
rect 25742 13640 25747 13696
rect 25405 13638 25747 13640
rect 22093 13635 22159 13638
rect 25405 13635 25471 13638
rect 25681 13635 25747 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 6361 13562 6427 13565
rect 9581 13562 9647 13565
rect 22277 13562 22343 13565
rect 6361 13560 9647 13562
rect 6361 13504 6366 13560
rect 6422 13504 9586 13560
rect 9642 13504 9647 13560
rect 6361 13502 9647 13504
rect 6361 13499 6427 13502
rect 9581 13499 9647 13502
rect 17174 13560 22343 13562
rect 17174 13504 22282 13560
rect 22338 13504 22343 13560
rect 17174 13502 22343 13504
rect 2129 13426 2195 13429
rect 17174 13426 17234 13502
rect 22277 13499 22343 13502
rect 2129 13424 17234 13426
rect 2129 13368 2134 13424
rect 2190 13368 17234 13424
rect 2129 13366 17234 13368
rect 17493 13426 17559 13429
rect 20437 13426 20503 13429
rect 17493 13424 20503 13426
rect 17493 13368 17498 13424
rect 17554 13368 20442 13424
rect 20498 13368 20503 13424
rect 17493 13366 20503 13368
rect 2129 13363 2195 13366
rect 17493 13363 17559 13366
rect 20437 13363 20503 13366
rect 22001 13426 22067 13429
rect 26200 13426 27000 13456
rect 22001 13424 27000 13426
rect 22001 13368 22006 13424
rect 22062 13368 27000 13424
rect 22001 13366 27000 13368
rect 22001 13363 22067 13366
rect 26200 13336 27000 13366
rect 5441 13290 5507 13293
rect 16982 13290 16988 13292
rect 5441 13288 16988 13290
rect 5441 13232 5446 13288
rect 5502 13232 16988 13288
rect 5441 13230 16988 13232
rect 5441 13227 5507 13230
rect 16982 13228 16988 13230
rect 17052 13228 17058 13292
rect 23422 13290 23428 13292
rect 17174 13230 23428 13290
rect 9673 13154 9739 13157
rect 13670 13154 13676 13156
rect 9673 13152 13676 13154
rect 9673 13096 9678 13152
rect 9734 13096 13676 13152
rect 9673 13094 13676 13096
rect 9673 13091 9739 13094
rect 13670 13092 13676 13094
rect 13740 13092 13746 13156
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 13854 13018 13860 13020
rect 9446 12958 13860 13018
rect 2129 12882 2195 12885
rect 2262 12882 2268 12884
rect 2129 12880 2268 12882
rect 2129 12824 2134 12880
rect 2190 12824 2268 12880
rect 2129 12822 2268 12824
rect 2129 12819 2195 12822
rect 2262 12820 2268 12822
rect 2332 12820 2338 12884
rect 6545 12882 6611 12885
rect 9446 12882 9506 12958
rect 13854 12956 13860 12958
rect 13924 12956 13930 13020
rect 6545 12880 9506 12882
rect 6545 12824 6550 12880
rect 6606 12824 9506 12880
rect 6545 12822 9506 12824
rect 9581 12882 9647 12885
rect 17174 12882 17234 13230
rect 23422 13228 23428 13230
rect 23492 13228 23498 13292
rect 18781 13154 18847 13157
rect 21817 13154 21883 13157
rect 18781 13152 21883 13154
rect 18781 13096 18786 13152
rect 18842 13096 21822 13152
rect 21878 13096 21883 13152
rect 18781 13094 21883 13096
rect 18781 13091 18847 13094
rect 21817 13091 21883 13094
rect 22277 13154 22343 13157
rect 25037 13154 25103 13157
rect 22277 13152 25103 13154
rect 22277 13096 22282 13152
rect 22338 13096 25042 13152
rect 25098 13096 25103 13152
rect 22277 13094 25103 13096
rect 22277 13091 22343 13094
rect 25037 13091 25103 13094
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 22553 13018 22619 13021
rect 26200 13018 27000 13048
rect 22553 13016 27000 13018
rect 22553 12960 22558 13016
rect 22614 12960 27000 13016
rect 22553 12958 27000 12960
rect 22553 12955 22619 12958
rect 26200 12928 27000 12958
rect 9581 12880 17234 12882
rect 9581 12824 9586 12880
rect 9642 12824 17234 12880
rect 9581 12822 17234 12824
rect 17769 12882 17835 12885
rect 18229 12882 18295 12885
rect 17769 12880 18295 12882
rect 17769 12824 17774 12880
rect 17830 12824 18234 12880
rect 18290 12824 18295 12880
rect 17769 12822 18295 12824
rect 6545 12819 6611 12822
rect 9581 12819 9647 12822
rect 17769 12819 17835 12822
rect 18229 12819 18295 12822
rect 5349 12746 5415 12749
rect 25681 12746 25747 12749
rect 5349 12744 25747 12746
rect 5349 12688 5354 12744
rect 5410 12688 25686 12744
rect 25742 12688 25747 12744
rect 5349 12686 25747 12688
rect 5349 12683 5415 12686
rect 25681 12683 25747 12686
rect 13537 12610 13603 12613
rect 18781 12610 18847 12613
rect 13537 12608 18847 12610
rect 13537 12552 13542 12608
rect 13598 12552 18786 12608
rect 18842 12552 18847 12608
rect 13537 12550 18847 12552
rect 13537 12547 13603 12550
rect 18781 12547 18847 12550
rect 25129 12610 25195 12613
rect 26200 12610 27000 12640
rect 25129 12608 27000 12610
rect 25129 12552 25134 12608
rect 25190 12552 27000 12608
rect 25129 12550 27000 12552
rect 25129 12547 25195 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 8293 12474 8359 12477
rect 16297 12474 16363 12477
rect 8293 12472 12818 12474
rect 8293 12416 8298 12472
rect 8354 12416 12818 12472
rect 8293 12414 12818 12416
rect 8293 12411 8359 12414
rect 3509 12338 3575 12341
rect 12758 12338 12818 12414
rect 13494 12472 16363 12474
rect 13494 12416 16302 12472
rect 16358 12416 16363 12472
rect 13494 12414 16363 12416
rect 13494 12338 13554 12414
rect 16297 12411 16363 12414
rect 16941 12474 17007 12477
rect 17861 12474 17927 12477
rect 16941 12472 17927 12474
rect 16941 12416 16946 12472
rect 17002 12416 17866 12472
rect 17922 12416 17927 12472
rect 16941 12414 17927 12416
rect 16941 12411 17007 12414
rect 17861 12411 17927 12414
rect 3509 12336 12634 12338
rect 3509 12280 3514 12336
rect 3570 12280 12634 12336
rect 3509 12278 12634 12280
rect 12758 12278 13554 12338
rect 15469 12340 15535 12341
rect 15469 12336 15516 12340
rect 15580 12338 15586 12340
rect 19793 12338 19859 12341
rect 20989 12338 21055 12341
rect 15469 12280 15474 12336
rect 3509 12275 3575 12278
rect 7005 12202 7071 12205
rect 9213 12202 9279 12205
rect 12382 12202 12388 12204
rect 7005 12200 8402 12202
rect 7005 12144 7010 12200
rect 7066 12144 8402 12200
rect 7005 12142 8402 12144
rect 7005 12139 7071 12142
rect 8342 12066 8402 12142
rect 9213 12200 12388 12202
rect 9213 12144 9218 12200
rect 9274 12144 12388 12200
rect 9213 12142 12388 12144
rect 9213 12139 9279 12142
rect 12382 12140 12388 12142
rect 12452 12140 12458 12204
rect 12574 12202 12634 12278
rect 15469 12276 15516 12280
rect 15580 12278 15626 12338
rect 19793 12336 21055 12338
rect 19793 12280 19798 12336
rect 19854 12280 20994 12336
rect 21050 12280 21055 12336
rect 19793 12278 21055 12280
rect 15580 12276 15586 12278
rect 15469 12275 15535 12276
rect 19793 12275 19859 12278
rect 20989 12275 21055 12278
rect 21817 12338 21883 12341
rect 24526 12338 24532 12340
rect 21817 12336 24532 12338
rect 21817 12280 21822 12336
rect 21878 12280 24532 12336
rect 21817 12278 24532 12280
rect 21817 12275 21883 12278
rect 24526 12276 24532 12278
rect 24596 12276 24602 12340
rect 12750 12202 12756 12204
rect 12574 12142 12756 12202
rect 12750 12140 12756 12142
rect 12820 12140 12826 12204
rect 15469 12202 15535 12205
rect 15878 12202 15884 12204
rect 15469 12200 15884 12202
rect 15469 12144 15474 12200
rect 15530 12144 15884 12200
rect 15469 12142 15884 12144
rect 15469 12139 15535 12142
rect 15878 12140 15884 12142
rect 15948 12140 15954 12204
rect 24761 12202 24827 12205
rect 26200 12202 27000 12232
rect 24761 12200 27000 12202
rect 24761 12144 24766 12200
rect 24822 12144 27000 12200
rect 24761 12142 27000 12144
rect 24761 12139 24827 12142
rect 26200 12112 27000 12142
rect 17534 12066 17540 12068
rect 8342 12006 17540 12066
rect 17534 12004 17540 12006
rect 17604 12004 17610 12068
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 12382 11868 12388 11932
rect 12452 11930 12458 11932
rect 12452 11870 15762 11930
rect 12452 11868 12458 11870
rect 7373 11794 7439 11797
rect 15469 11794 15535 11797
rect 7373 11792 15535 11794
rect 7373 11736 7378 11792
rect 7434 11736 15474 11792
rect 15530 11736 15535 11792
rect 7373 11734 15535 11736
rect 15702 11794 15762 11870
rect 21398 11794 21404 11796
rect 15702 11734 21404 11794
rect 7373 11731 7439 11734
rect 15469 11731 15535 11734
rect 21398 11732 21404 11734
rect 21468 11732 21474 11796
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 1945 11658 2011 11661
rect 15142 11658 15148 11660
rect 1945 11656 15148 11658
rect 1945 11600 1950 11656
rect 2006 11600 15148 11656
rect 1945 11598 15148 11600
rect 1945 11595 2011 11598
rect 15142 11596 15148 11598
rect 15212 11596 15218 11660
rect 16481 11658 16547 11661
rect 25957 11658 26023 11661
rect 16481 11656 26023 11658
rect 16481 11600 16486 11656
rect 16542 11600 25962 11656
rect 26018 11600 26023 11656
rect 16481 11598 26023 11600
rect 16481 11595 16547 11598
rect 25957 11595 26023 11598
rect 13721 11522 13787 11525
rect 19190 11522 19196 11524
rect 13721 11520 19196 11522
rect 13721 11464 13726 11520
rect 13782 11464 19196 11520
rect 13721 11462 19196 11464
rect 13721 11459 13787 11462
rect 19190 11460 19196 11462
rect 19260 11460 19266 11524
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 14549 11386 14615 11389
rect 21030 11386 21036 11388
rect 14549 11384 21036 11386
rect 14549 11328 14554 11384
rect 14610 11328 21036 11384
rect 14549 11326 21036 11328
rect 14549 11323 14615 11326
rect 21030 11324 21036 11326
rect 21100 11386 21106 11388
rect 21725 11386 21791 11389
rect 21100 11384 21791 11386
rect 21100 11328 21730 11384
rect 21786 11328 21791 11384
rect 21100 11326 21791 11328
rect 21100 11324 21106 11326
rect 21725 11323 21791 11326
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 5809 11250 5875 11253
rect 16757 11252 16823 11253
rect 16757 11250 16804 11252
rect 5809 11248 16804 11250
rect 16868 11250 16874 11252
rect 20437 11250 20503 11253
rect 20846 11250 20852 11252
rect 5809 11192 5814 11248
rect 5870 11192 16762 11248
rect 5809 11190 16804 11192
rect 5809 11187 5875 11190
rect 16757 11188 16804 11190
rect 16868 11190 16950 11250
rect 20437 11248 20852 11250
rect 20437 11192 20442 11248
rect 20498 11192 20852 11248
rect 20437 11190 20852 11192
rect 16868 11188 16874 11190
rect 16757 11187 16823 11188
rect 20437 11187 20503 11190
rect 20846 11188 20852 11190
rect 20916 11188 20922 11252
rect 5625 11114 5691 11117
rect 14549 11114 14615 11117
rect 5625 11112 14615 11114
rect 5625 11056 5630 11112
rect 5686 11056 14554 11112
rect 14610 11056 14615 11112
rect 5625 11054 14615 11056
rect 5625 11051 5691 11054
rect 14549 11051 14615 11054
rect 14774 11052 14780 11116
rect 14844 11114 14850 11116
rect 15009 11114 15075 11117
rect 14844 11112 15075 11114
rect 14844 11056 15014 11112
rect 15070 11056 15075 11112
rect 14844 11054 15075 11056
rect 14844 11052 14850 11054
rect 15009 11051 15075 11054
rect 18638 11052 18644 11116
rect 18708 11114 18714 11116
rect 18781 11114 18847 11117
rect 18708 11112 18847 11114
rect 18708 11056 18786 11112
rect 18842 11056 18847 11112
rect 18708 11054 18847 11056
rect 18708 11052 18714 11054
rect 18781 11051 18847 11054
rect 19885 11114 19951 11117
rect 20805 11114 20871 11117
rect 19885 11112 20871 11114
rect 19885 11056 19890 11112
rect 19946 11056 20810 11112
rect 20866 11056 20871 11112
rect 19885 11054 20871 11056
rect 19885 11051 19951 11054
rect 20805 11051 20871 11054
rect 25129 10978 25195 10981
rect 26200 10978 27000 11008
rect 25129 10976 27000 10978
rect 25129 10920 25134 10976
rect 25190 10920 27000 10976
rect 25129 10918 27000 10920
rect 25129 10915 25195 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 24669 10842 24735 10845
rect 18462 10840 24735 10842
rect 18462 10784 24674 10840
rect 24730 10784 24735 10840
rect 18462 10782 24735 10784
rect 3969 10706 4035 10709
rect 3969 10704 6930 10706
rect 3969 10648 3974 10704
rect 4030 10648 6930 10704
rect 3969 10646 6930 10648
rect 3969 10643 4035 10646
rect 6870 10570 6930 10646
rect 18462 10570 18522 10782
rect 24669 10779 24735 10782
rect 23974 10706 23980 10708
rect 6870 10510 18522 10570
rect 18784 10646 23980 10706
rect 17125 10434 17191 10437
rect 18784 10434 18844 10646
rect 23974 10644 23980 10646
rect 24044 10644 24050 10708
rect 19057 10570 19123 10573
rect 22686 10570 22692 10572
rect 19057 10568 22692 10570
rect 19057 10512 19062 10568
rect 19118 10512 22692 10568
rect 19057 10510 22692 10512
rect 19057 10507 19123 10510
rect 22686 10508 22692 10510
rect 22756 10508 22762 10572
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 17125 10432 18844 10434
rect 17125 10376 17130 10432
rect 17186 10376 18844 10432
rect 17125 10374 18844 10376
rect 17125 10371 17191 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 17217 10298 17283 10301
rect 20110 10298 20116 10300
rect 17217 10296 20116 10298
rect 17217 10240 17222 10296
rect 17278 10240 20116 10296
rect 17217 10238 20116 10240
rect 17217 10235 17283 10238
rect 20110 10236 20116 10238
rect 20180 10236 20186 10300
rect 14958 10100 14964 10164
rect 15028 10162 15034 10164
rect 15285 10162 15351 10165
rect 15028 10160 15351 10162
rect 15028 10104 15290 10160
rect 15346 10104 15351 10160
rect 15028 10102 15351 10104
rect 15028 10100 15034 10102
rect 15285 10099 15351 10102
rect 18321 10162 18387 10165
rect 23606 10162 23612 10164
rect 18321 10160 23612 10162
rect 18321 10104 18326 10160
rect 18382 10104 23612 10160
rect 18321 10102 23612 10104
rect 18321 10099 18387 10102
rect 23606 10100 23612 10102
rect 23676 10100 23682 10164
rect 24761 10162 24827 10165
rect 26200 10162 27000 10192
rect 24761 10160 27000 10162
rect 24761 10104 24766 10160
rect 24822 10104 27000 10160
rect 24761 10102 27000 10104
rect 24761 10099 24827 10102
rect 26200 10072 27000 10102
rect 20345 9890 20411 9893
rect 21214 9890 21220 9892
rect 20345 9888 21220 9890
rect 20345 9832 20350 9888
rect 20406 9832 21220 9888
rect 20345 9830 21220 9832
rect 20345 9827 20411 9830
rect 21214 9828 21220 9830
rect 21284 9828 21290 9892
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 19425 9754 19491 9757
rect 20294 9754 20300 9756
rect 19425 9752 20300 9754
rect 19425 9696 19430 9752
rect 19486 9696 20300 9752
rect 19425 9694 20300 9696
rect 19425 9691 19491 9694
rect 20294 9692 20300 9694
rect 20364 9692 20370 9756
rect 21222 9754 21282 9828
rect 21357 9754 21423 9757
rect 21222 9752 21423 9754
rect 21222 9696 21362 9752
rect 21418 9696 21423 9752
rect 21222 9694 21423 9696
rect 21357 9691 21423 9694
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 1761 9618 1827 9621
rect 15653 9620 15719 9621
rect 15653 9618 15700 9620
rect 1761 9616 6930 9618
rect 1761 9560 1766 9616
rect 1822 9560 6930 9616
rect 1761 9558 6930 9560
rect 15608 9616 15700 9618
rect 15608 9560 15658 9616
rect 15608 9558 15700 9560
rect 1761 9555 1827 9558
rect 6870 9482 6930 9558
rect 15653 9556 15700 9558
rect 15764 9556 15770 9620
rect 20529 9618 20595 9621
rect 20662 9618 20668 9620
rect 20529 9616 20668 9618
rect 20529 9560 20534 9616
rect 20590 9560 20668 9616
rect 20529 9558 20668 9560
rect 15653 9555 15719 9556
rect 20529 9555 20595 9558
rect 20662 9556 20668 9558
rect 20732 9556 20738 9620
rect 21173 9482 21239 9485
rect 22093 9482 22159 9485
rect 6870 9480 21239 9482
rect 6870 9424 21178 9480
rect 21234 9424 21239 9480
rect 6870 9422 21239 9424
rect 21173 9419 21239 9422
rect 22050 9480 22159 9482
rect 22050 9424 22098 9480
rect 22154 9424 22159 9480
rect 22050 9419 22159 9424
rect 22050 9349 22110 9419
rect 20989 9346 21055 9349
rect 21449 9346 21515 9349
rect 22001 9346 22110 9349
rect 20989 9344 21515 9346
rect 20989 9288 20994 9344
rect 21050 9288 21454 9344
rect 21510 9288 21515 9344
rect 20989 9286 21515 9288
rect 21966 9344 22110 9346
rect 21966 9288 22006 9344
rect 22062 9288 22110 9344
rect 21966 9286 22110 9288
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 20989 9283 21055 9286
rect 21449 9283 21515 9286
rect 22001 9283 22067 9286
rect 24853 9283 24919 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 18781 9210 18847 9213
rect 19006 9210 19012 9212
rect 18781 9208 19012 9210
rect 18781 9152 18786 9208
rect 18842 9152 19012 9208
rect 18781 9150 19012 9152
rect 18781 9147 18847 9150
rect 19006 9148 19012 9150
rect 19076 9148 19082 9212
rect 19149 9210 19215 9213
rect 21817 9210 21883 9213
rect 25957 9210 26023 9213
rect 19149 9208 21883 9210
rect 19149 9152 19154 9208
rect 19210 9152 21822 9208
rect 21878 9152 21883 9208
rect 19149 9150 21883 9152
rect 19149 9147 19215 9150
rect 21817 9147 21883 9150
rect 23798 9208 26023 9210
rect 23798 9152 25962 9208
rect 26018 9152 26023 9208
rect 23798 9150 26023 9152
rect 19333 9074 19399 9077
rect 23798 9074 23858 9150
rect 25957 9147 26023 9150
rect 26049 9074 26115 9077
rect 19333 9072 23858 9074
rect 19333 9016 19338 9072
rect 19394 9016 23858 9072
rect 19333 9014 23858 9016
rect 23982 9072 26115 9074
rect 23982 9016 26054 9072
rect 26110 9016 26115 9072
rect 23982 9014 26115 9016
rect 19333 9011 19399 9014
rect 16297 8938 16363 8941
rect 23982 8938 24042 9014
rect 26049 9011 26115 9014
rect 16297 8936 24042 8938
rect 16297 8880 16302 8936
rect 16358 8880 24042 8936
rect 16297 8878 24042 8880
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 16297 8875 16363 8878
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 20805 8802 20871 8805
rect 21030 8802 21036 8804
rect 20805 8800 21036 8802
rect 20805 8744 20810 8800
rect 20866 8744 21036 8800
rect 20805 8742 21036 8744
rect 20805 8739 20871 8742
rect 21030 8740 21036 8742
rect 21100 8740 21106 8804
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 19793 8666 19859 8669
rect 19926 8666 19932 8668
rect 19793 8664 19932 8666
rect 19793 8608 19798 8664
rect 19854 8608 19932 8664
rect 19793 8606 19932 8608
rect 19793 8603 19859 8606
rect 19926 8604 19932 8606
rect 19996 8604 20002 8668
rect 24945 8530 25011 8533
rect 26200 8530 27000 8560
rect 24945 8528 27000 8530
rect 24945 8472 24950 8528
rect 25006 8472 27000 8528
rect 24945 8470 27000 8472
rect 24945 8467 25011 8470
rect 26200 8440 27000 8470
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 19425 8122 19491 8125
rect 19558 8122 19564 8124
rect 19425 8120 19564 8122
rect 19425 8064 19430 8120
rect 19486 8064 19564 8120
rect 19425 8062 19564 8064
rect 19425 8059 19491 8062
rect 19558 8060 19564 8062
rect 19628 8060 19634 8124
rect 24853 8122 24919 8125
rect 26200 8122 27000 8152
rect 24853 8120 27000 8122
rect 24853 8064 24858 8120
rect 24914 8064 27000 8120
rect 24853 8062 27000 8064
rect 24853 8059 24919 8062
rect 26200 8032 27000 8062
rect 4981 7986 5047 7989
rect 25405 7986 25471 7989
rect 4981 7984 25471 7986
rect 4981 7928 4986 7984
rect 5042 7928 25410 7984
rect 25466 7928 25471 7984
rect 4981 7926 25471 7928
rect 4981 7923 5047 7926
rect 25405 7923 25471 7926
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 24485 6900 24551 6901
rect 24669 6900 24735 6901
rect 24485 6898 24532 6900
rect 24440 6896 24532 6898
rect 24440 6840 24490 6896
rect 24440 6838 24532 6840
rect 24485 6836 24532 6838
rect 24596 6836 24602 6900
rect 24669 6896 24716 6900
rect 24780 6898 24786 6900
rect 24945 6898 25011 6901
rect 26200 6898 27000 6928
rect 24669 6840 24674 6896
rect 24669 6836 24716 6840
rect 24780 6838 24826 6898
rect 24945 6896 27000 6898
rect 24945 6840 24950 6896
rect 25006 6840 27000 6896
rect 24945 6838 27000 6840
rect 24780 6836 24786 6838
rect 24485 6835 24551 6836
rect 24669 6835 24735 6836
rect 24945 6835 25011 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 22277 5268 22343 5269
rect 22277 5266 22324 5268
rect 22232 5264 22324 5266
rect 22232 5208 22282 5264
rect 22232 5206 22324 5208
rect 22277 5204 22324 5206
rect 22388 5204 22394 5268
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 22277 5203 22343 5204
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24853 4858 24919 4861
rect 26200 4858 27000 4888
rect 24853 4856 27000 4858
rect 24853 4800 24858 4856
rect 24914 4800 27000 4856
rect 24853 4798 27000 4800
rect 24853 4795 24919 4798
rect 26200 4768 27000 4798
rect 25497 4450 25563 4453
rect 26200 4450 27000 4480
rect 25497 4448 27000 4450
rect 25497 4392 25502 4448
rect 25558 4392 27000 4448
rect 25497 4390 27000 4392
rect 25497 4387 25563 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25129 4042 25195 4045
rect 26200 4042 27000 4072
rect 25129 4040 27000 4042
rect 25129 3984 25134 4040
rect 25190 3984 27000 4040
rect 25129 3982 27000 3984
rect 25129 3979 25195 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 24945 3226 25011 3229
rect 26200 3226 27000 3256
rect 24945 3224 27000 3226
rect 24945 3168 24950 3224
rect 25006 3168 27000 3224
rect 24945 3166 27000 3168
rect 24945 3163 25011 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22093 2002 22159 2005
rect 26200 2002 27000 2032
rect 22093 2000 27000 2002
rect 22093 1944 22098 2000
rect 22154 1944 27000 2000
rect 22093 1942 27000 1944
rect 22093 1939 22159 1942
rect 26200 1912 27000 1942
rect 22185 1594 22251 1597
rect 26200 1594 27000 1624
rect 22185 1592 27000 1594
rect 22185 1536 22190 1592
rect 22246 1536 27000 1592
rect 22185 1534 27000 1536
rect 22185 1531 22251 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 16620 26828 16684 26892
rect 10180 26692 10244 26756
rect 15332 26556 15396 26620
rect 21404 26420 21468 26484
rect 2636 26284 2700 26348
rect 5396 26148 5460 26212
rect 5580 26012 5644 26076
rect 2268 25740 2332 25804
rect 6500 25604 6564 25668
rect 7604 25332 7668 25396
rect 4660 25196 4724 25260
rect 16436 24924 16500 24988
rect 5948 24788 6012 24852
rect 7788 24652 7852 24716
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 18460 24380 18524 24444
rect 11652 24244 11716 24308
rect 8524 24108 8588 24172
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 23980 23972 24044 24036
rect 5764 23428 5828 23492
rect 9996 23488 10060 23492
rect 9996 23432 10046 23488
rect 10046 23432 10060 23488
rect 9996 23428 10060 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 14964 23564 15028 23628
rect 13860 23488 13924 23492
rect 13860 23432 13874 23488
rect 13874 23432 13924 23488
rect 13860 23428 13924 23432
rect 14044 23428 14108 23492
rect 15148 23428 15212 23492
rect 16068 23428 16132 23492
rect 19564 23428 19628 23492
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 12756 23156 12820 23220
rect 13676 23156 13740 23220
rect 9260 22884 9324 22948
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 16620 22340 16684 22404
rect 18644 22340 18708 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 16436 22204 16500 22268
rect 21956 22068 22020 22132
rect 9812 21796 9876 21860
rect 21404 21796 21468 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 11468 21660 11532 21724
rect 18460 21660 18524 21724
rect 13492 21524 13556 21588
rect 16068 21388 16132 21452
rect 17540 21448 17604 21452
rect 17540 21392 17554 21448
rect 17554 21392 17604 21448
rect 17540 21388 17604 21392
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 9628 20980 9692 21044
rect 5764 20708 5828 20772
rect 16620 20708 16684 20772
rect 17172 20708 17236 20772
rect 19932 20768 19996 20772
rect 19932 20712 19946 20768
rect 19946 20712 19996 20768
rect 19932 20708 19996 20712
rect 21220 20768 21284 20772
rect 21220 20712 21234 20768
rect 21234 20712 21284 20768
rect 21220 20708 21284 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 12572 20572 12636 20636
rect 15332 20572 15396 20636
rect 22508 20572 22572 20636
rect 15516 20164 15580 20228
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 12572 19892 12636 19956
rect 15700 20028 15764 20092
rect 16804 20164 16868 20228
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 20116 19620 20180 19684
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 15700 19484 15764 19548
rect 20668 19484 20732 19548
rect 14780 19348 14844 19412
rect 20852 19348 20916 19412
rect 22324 19348 22388 19412
rect 18460 19076 18524 19140
rect 20300 19212 20364 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 10916 18940 10980 19004
rect 18828 18940 18892 19004
rect 9260 18668 9324 18732
rect 23428 18668 23492 18732
rect 11100 18532 11164 18596
rect 15148 18532 15212 18596
rect 22140 18532 22204 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 7788 18396 7852 18460
rect 3372 17988 3436 18052
rect 5948 17988 6012 18052
rect 7604 17988 7668 18052
rect 11468 17988 11532 18052
rect 23612 17988 23676 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 8524 17852 8588 17916
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 16988 17172 17052 17236
rect 22324 17172 22388 17236
rect 11652 16900 11716 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 10180 16764 10244 16828
rect 11468 16824 11532 16828
rect 11468 16768 11518 16824
rect 11518 16768 11532 16824
rect 11468 16764 11532 16768
rect 15884 16764 15948 16828
rect 22692 16628 22756 16692
rect 24532 16628 24596 16692
rect 16436 16356 16500 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 6500 16220 6564 16284
rect 16988 16084 17052 16148
rect 10916 15812 10980 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 18828 15676 18892 15740
rect 5396 15540 5460 15604
rect 21404 15540 21468 15604
rect 22140 15404 22204 15468
rect 19196 15268 19260 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 4660 15132 4724 15196
rect 14044 15132 14108 15196
rect 3372 14996 3436 15060
rect 18460 14860 18524 14924
rect 19012 14860 19076 14924
rect 21956 14860 22020 14924
rect 9996 14724 10060 14788
rect 15148 14724 15212 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 22508 14588 22572 14652
rect 2636 14452 2700 14516
rect 5580 14512 5644 14516
rect 5580 14456 5594 14512
rect 5594 14456 5644 14512
rect 5580 14452 5644 14456
rect 9628 14452 9692 14516
rect 11100 14180 11164 14244
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 9812 13772 9876 13836
rect 13492 13772 13556 13836
rect 22324 13908 22388 13972
rect 24716 13908 24780 13972
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 16988 13228 17052 13292
rect 13676 13092 13740 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 2268 12820 2332 12884
rect 13860 12956 13924 13020
rect 23428 13228 23492 13292
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 15516 12336 15580 12340
rect 15516 12280 15530 12336
rect 15530 12280 15580 12336
rect 12388 12140 12452 12204
rect 15516 12276 15580 12280
rect 24532 12276 24596 12340
rect 12756 12140 12820 12204
rect 15884 12140 15948 12204
rect 17540 12004 17604 12068
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 12388 11868 12452 11932
rect 21404 11732 21468 11796
rect 15148 11596 15212 11660
rect 19196 11460 19260 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 21036 11324 21100 11388
rect 16804 11248 16868 11252
rect 16804 11192 16818 11248
rect 16818 11192 16868 11248
rect 16804 11188 16868 11192
rect 20852 11188 20916 11252
rect 14780 11052 14844 11116
rect 18644 11052 18708 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 23980 10644 24044 10708
rect 22692 10508 22756 10572
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 20116 10236 20180 10300
rect 14964 10100 15028 10164
rect 23612 10100 23676 10164
rect 21220 9828 21284 9892
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 20300 9692 20364 9756
rect 15700 9616 15764 9620
rect 15700 9560 15714 9616
rect 15714 9560 15764 9616
rect 15700 9556 15764 9560
rect 20668 9556 20732 9620
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 19012 9148 19076 9212
rect 21036 8740 21100 8804
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 19932 8604 19996 8668
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 19564 8060 19628 8124
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 24532 6896 24596 6900
rect 24532 6840 24546 6896
rect 24546 6840 24596 6896
rect 24532 6836 24596 6840
rect 24716 6896 24780 6900
rect 24716 6840 24730 6896
rect 24730 6840 24780 6896
rect 24716 6836 24780 6840
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 22324 5264 22388 5268
rect 22324 5208 22338 5264
rect 22338 5208 22388 5264
rect 22324 5204 22388 5208
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 16619 26892 16685 26893
rect 16619 26828 16620 26892
rect 16684 26828 16685 26892
rect 16619 26827 16685 26828
rect 10179 26756 10245 26757
rect 10179 26692 10180 26756
rect 10244 26692 10245 26756
rect 10179 26691 10245 26692
rect 2635 26348 2701 26349
rect 2635 26284 2636 26348
rect 2700 26284 2701 26348
rect 2635 26283 2701 26284
rect 2267 25804 2333 25805
rect 2267 25740 2268 25804
rect 2332 25740 2333 25804
rect 2267 25739 2333 25740
rect 2270 12885 2330 25739
rect 2638 14517 2698 26283
rect 5395 26212 5461 26213
rect 5395 26148 5396 26212
rect 5460 26148 5461 26212
rect 5395 26147 5461 26148
rect 4659 25260 4725 25261
rect 4659 25196 4660 25260
rect 4724 25196 4725 25260
rect 4659 25195 4725 25196
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 3371 18052 3437 18053
rect 3371 17988 3372 18052
rect 3436 17988 3437 18052
rect 3371 17987 3437 17988
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 3374 15061 3434 17987
rect 4662 15197 4722 25195
rect 5398 15605 5458 26147
rect 5579 26076 5645 26077
rect 5579 26012 5580 26076
rect 5644 26012 5645 26076
rect 5579 26011 5645 26012
rect 5395 15604 5461 15605
rect 5395 15540 5396 15604
rect 5460 15540 5461 15604
rect 5395 15539 5461 15540
rect 4659 15196 4725 15197
rect 4659 15132 4660 15196
rect 4724 15132 4725 15196
rect 4659 15131 4725 15132
rect 3371 15060 3437 15061
rect 3371 14996 3372 15060
rect 3436 14996 3437 15060
rect 3371 14995 3437 14996
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2635 14516 2701 14517
rect 2635 14452 2636 14516
rect 2700 14452 2701 14516
rect 2635 14451 2701 14452
rect 2944 13632 3264 14656
rect 5582 14517 5642 26011
rect 6499 25668 6565 25669
rect 6499 25604 6500 25668
rect 6564 25604 6565 25668
rect 6499 25603 6565 25604
rect 5947 24852 6013 24853
rect 5947 24788 5948 24852
rect 6012 24788 6013 24852
rect 5947 24787 6013 24788
rect 5763 23492 5829 23493
rect 5763 23428 5764 23492
rect 5828 23428 5829 23492
rect 5763 23427 5829 23428
rect 5766 20773 5826 23427
rect 5763 20772 5829 20773
rect 5763 20708 5764 20772
rect 5828 20708 5829 20772
rect 5763 20707 5829 20708
rect 5950 18053 6010 24787
rect 5947 18052 6013 18053
rect 5947 17988 5948 18052
rect 6012 17988 6013 18052
rect 5947 17987 6013 17988
rect 6502 16285 6562 25603
rect 7603 25396 7669 25397
rect 7603 25332 7604 25396
rect 7668 25332 7669 25396
rect 7603 25331 7669 25332
rect 7606 18053 7666 25331
rect 7787 24716 7853 24717
rect 7787 24652 7788 24716
rect 7852 24652 7853 24716
rect 7787 24651 7853 24652
rect 7790 18461 7850 24651
rect 7944 23968 8264 24528
rect 8523 24172 8589 24173
rect 8523 24108 8524 24172
rect 8588 24108 8589 24172
rect 8523 24107 8589 24108
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7787 18460 7853 18461
rect 7787 18396 7788 18460
rect 7852 18396 7853 18460
rect 7787 18395 7853 18396
rect 7603 18052 7669 18053
rect 7603 17988 7604 18052
rect 7668 17988 7669 18052
rect 7603 17987 7669 17988
rect 7944 17440 8264 18464
rect 8526 17917 8586 24107
rect 9995 23492 10061 23493
rect 9995 23428 9996 23492
rect 10060 23428 10061 23492
rect 9995 23427 10061 23428
rect 9259 22948 9325 22949
rect 9259 22884 9260 22948
rect 9324 22884 9325 22948
rect 9259 22883 9325 22884
rect 9262 18733 9322 22883
rect 9811 21860 9877 21861
rect 9811 21796 9812 21860
rect 9876 21796 9877 21860
rect 9811 21795 9877 21796
rect 9627 21044 9693 21045
rect 9627 20980 9628 21044
rect 9692 20980 9693 21044
rect 9627 20979 9693 20980
rect 9259 18732 9325 18733
rect 9259 18668 9260 18732
rect 9324 18668 9325 18732
rect 9259 18667 9325 18668
rect 8523 17916 8589 17917
rect 8523 17852 8524 17916
rect 8588 17852 8589 17916
rect 8523 17851 8589 17852
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 6499 16284 6565 16285
rect 6499 16220 6500 16284
rect 6564 16220 6565 16284
rect 6499 16219 6565 16220
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 5579 14516 5645 14517
rect 5579 14452 5580 14516
rect 5644 14452 5645 14516
rect 5579 14451 5645 14452
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2267 12884 2333 12885
rect 2267 12820 2268 12884
rect 2332 12820 2333 12884
rect 2267 12819 2333 12820
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 14176 8264 15200
rect 9630 14517 9690 20979
rect 9627 14516 9693 14517
rect 9627 14452 9628 14516
rect 9692 14452 9693 14516
rect 9627 14451 9693 14452
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 9814 13837 9874 21795
rect 9998 14789 10058 23427
rect 10182 16829 10242 26691
rect 15331 26620 15397 26621
rect 15331 26556 15332 26620
rect 15396 26556 15397 26620
rect 15331 26555 15397 26556
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 11651 24308 11717 24309
rect 11651 24244 11652 24308
rect 11716 24244 11717 24308
rect 11651 24243 11717 24244
rect 11467 21724 11533 21725
rect 11467 21660 11468 21724
rect 11532 21660 11533 21724
rect 11467 21659 11533 21660
rect 10915 19004 10981 19005
rect 10915 18940 10916 19004
rect 10980 18940 10981 19004
rect 10915 18939 10981 18940
rect 10179 16828 10245 16829
rect 10179 16764 10180 16828
rect 10244 16764 10245 16828
rect 10179 16763 10245 16764
rect 10918 15877 10978 18939
rect 11099 18596 11165 18597
rect 11099 18532 11100 18596
rect 11164 18532 11165 18596
rect 11099 18531 11165 18532
rect 10915 15876 10981 15877
rect 10915 15812 10916 15876
rect 10980 15812 10981 15876
rect 10915 15811 10981 15812
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 11102 14245 11162 18531
rect 11470 18053 11530 21659
rect 11467 18052 11533 18053
rect 11467 17988 11468 18052
rect 11532 17988 11533 18052
rect 11467 17987 11533 17988
rect 11470 16829 11530 17987
rect 11654 16965 11714 24243
rect 12944 23424 13264 24448
rect 14963 23628 15029 23629
rect 14963 23564 14964 23628
rect 15028 23564 15029 23628
rect 14963 23563 15029 23564
rect 13859 23492 13925 23493
rect 13859 23428 13860 23492
rect 13924 23428 13925 23492
rect 13859 23427 13925 23428
rect 14043 23492 14109 23493
rect 14043 23428 14044 23492
rect 14108 23428 14109 23492
rect 14043 23427 14109 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12755 23220 12821 23221
rect 12755 23156 12756 23220
rect 12820 23156 12821 23220
rect 12755 23155 12821 23156
rect 12571 20636 12637 20637
rect 12571 20572 12572 20636
rect 12636 20572 12637 20636
rect 12571 20571 12637 20572
rect 12574 19957 12634 20571
rect 12571 19956 12637 19957
rect 12571 19892 12572 19956
rect 12636 19892 12637 19956
rect 12571 19891 12637 19892
rect 11651 16964 11717 16965
rect 11651 16900 11652 16964
rect 11716 16900 11717 16964
rect 11651 16899 11717 16900
rect 11467 16828 11533 16829
rect 11467 16764 11468 16828
rect 11532 16764 11533 16828
rect 11467 16763 11533 16764
rect 11099 14244 11165 14245
rect 11099 14180 11100 14244
rect 11164 14180 11165 14244
rect 11099 14179 11165 14180
rect 9811 13836 9877 13837
rect 9811 13772 9812 13836
rect 9876 13772 9877 13836
rect 9811 13771 9877 13772
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 12758 12205 12818 23155
rect 12944 22336 13264 23360
rect 13675 23220 13741 23221
rect 13675 23156 13676 23220
rect 13740 23156 13741 23220
rect 13675 23155 13741 23156
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 13491 21588 13557 21589
rect 13491 21524 13492 21588
rect 13556 21524 13557 21588
rect 13491 21523 13557 21524
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13494 13837 13554 21523
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 13678 13157 13738 23155
rect 13675 13156 13741 13157
rect 13675 13092 13676 13156
rect 13740 13092 13741 13156
rect 13675 13091 13741 13092
rect 13862 13021 13922 23427
rect 14046 15197 14106 23427
rect 14779 19412 14845 19413
rect 14779 19348 14780 19412
rect 14844 19348 14845 19412
rect 14779 19347 14845 19348
rect 14043 15196 14109 15197
rect 14043 15132 14044 15196
rect 14108 15132 14109 15196
rect 14043 15131 14109 15132
rect 13859 13020 13925 13021
rect 13859 12956 13860 13020
rect 13924 12956 13925 13020
rect 13859 12955 13925 12956
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12387 12204 12453 12205
rect 12387 12140 12388 12204
rect 12452 12140 12453 12204
rect 12387 12139 12453 12140
rect 12755 12204 12821 12205
rect 12755 12140 12756 12204
rect 12820 12140 12821 12204
rect 12755 12139 12821 12140
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 12390 11933 12450 12139
rect 12387 11932 12453 11933
rect 12387 11868 12388 11932
rect 12452 11868 12453 11932
rect 12387 11867 12453 11868
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 14782 11117 14842 19347
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 14966 10165 15026 23563
rect 15147 23492 15213 23493
rect 15147 23428 15148 23492
rect 15212 23428 15213 23492
rect 15147 23427 15213 23428
rect 15150 18597 15210 23427
rect 15334 20637 15394 26555
rect 16435 24988 16501 24989
rect 16435 24924 16436 24988
rect 16500 24924 16501 24988
rect 16435 24923 16501 24924
rect 16067 23492 16133 23493
rect 16067 23428 16068 23492
rect 16132 23428 16133 23492
rect 16067 23427 16133 23428
rect 16070 21453 16130 23427
rect 16438 22269 16498 24923
rect 16622 22405 16682 26827
rect 21403 26484 21469 26485
rect 21403 26420 21404 26484
rect 21468 26420 21469 26484
rect 21403 26419 21469 26420
rect 17944 23968 18264 24528
rect 18459 24444 18525 24445
rect 18459 24380 18460 24444
rect 18524 24380 18525 24444
rect 18459 24379 18525 24380
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 16619 22404 16685 22405
rect 16619 22340 16620 22404
rect 16684 22340 16685 22404
rect 16619 22339 16685 22340
rect 16435 22268 16501 22269
rect 16435 22204 16436 22268
rect 16500 22204 16501 22268
rect 16435 22203 16501 22204
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 16067 21452 16133 21453
rect 16067 21388 16068 21452
rect 16132 21388 16133 21452
rect 16067 21387 16133 21388
rect 17539 21452 17605 21453
rect 17539 21388 17540 21452
rect 17604 21388 17605 21452
rect 17539 21387 17605 21388
rect 16619 20772 16685 20773
rect 16619 20770 16620 20772
rect 16438 20710 16620 20770
rect 15331 20636 15397 20637
rect 15331 20572 15332 20636
rect 15396 20572 15397 20636
rect 15331 20571 15397 20572
rect 15515 20228 15581 20229
rect 15515 20164 15516 20228
rect 15580 20164 15581 20228
rect 15515 20163 15581 20164
rect 15147 18596 15213 18597
rect 15147 18532 15148 18596
rect 15212 18532 15213 18596
rect 15147 18531 15213 18532
rect 15147 14788 15213 14789
rect 15147 14724 15148 14788
rect 15212 14724 15213 14788
rect 15147 14723 15213 14724
rect 15150 11661 15210 14723
rect 15518 12341 15578 20163
rect 15699 20092 15765 20093
rect 15699 20028 15700 20092
rect 15764 20028 15765 20092
rect 15699 20027 15765 20028
rect 15702 19549 15762 20027
rect 15699 19548 15765 19549
rect 15699 19484 15700 19548
rect 15764 19484 15765 19548
rect 15699 19483 15765 19484
rect 15515 12340 15581 12341
rect 15515 12276 15516 12340
rect 15580 12276 15581 12340
rect 15515 12275 15581 12276
rect 15147 11660 15213 11661
rect 15147 11596 15148 11660
rect 15212 11596 15213 11660
rect 15147 11595 15213 11596
rect 14963 10164 15029 10165
rect 14963 10100 14964 10164
rect 15028 10100 15029 10164
rect 14963 10099 15029 10100
rect 15702 9621 15762 19483
rect 15883 16828 15949 16829
rect 15883 16764 15884 16828
rect 15948 16764 15949 16828
rect 15883 16763 15949 16764
rect 15886 12205 15946 16763
rect 16438 16421 16498 20710
rect 16619 20708 16620 20710
rect 16684 20708 16685 20772
rect 16619 20707 16685 20708
rect 17171 20772 17237 20773
rect 17171 20708 17172 20772
rect 17236 20708 17237 20772
rect 17171 20707 17237 20708
rect 16803 20228 16869 20229
rect 16803 20164 16804 20228
rect 16868 20164 16869 20228
rect 16803 20163 16869 20164
rect 16435 16420 16501 16421
rect 16435 16356 16436 16420
rect 16500 16356 16501 16420
rect 16435 16355 16501 16356
rect 15883 12204 15949 12205
rect 15883 12140 15884 12204
rect 15948 12140 15949 12204
rect 15883 12139 15949 12140
rect 16806 11253 16866 20163
rect 16987 17236 17053 17237
rect 16987 17172 16988 17236
rect 17052 17172 17053 17236
rect 16987 17171 17053 17172
rect 16990 16149 17050 17171
rect 16987 16148 17053 16149
rect 16987 16084 16988 16148
rect 17052 16084 17053 16148
rect 16987 16083 17053 16084
rect 16987 13292 17053 13293
rect 16987 13228 16988 13292
rect 17052 13290 17053 13292
rect 17174 13290 17234 20707
rect 17052 13230 17234 13290
rect 17052 13228 17053 13230
rect 16987 13227 17053 13228
rect 17542 12069 17602 21387
rect 17944 20704 18264 21728
rect 18462 21725 18522 24379
rect 19563 23492 19629 23493
rect 19563 23428 19564 23492
rect 19628 23428 19629 23492
rect 19563 23427 19629 23428
rect 18643 22404 18709 22405
rect 18643 22340 18644 22404
rect 18708 22340 18709 22404
rect 18643 22339 18709 22340
rect 18459 21724 18525 21725
rect 18459 21660 18460 21724
rect 18524 21660 18525 21724
rect 18459 21659 18525 21660
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18459 19140 18525 19141
rect 18459 19076 18460 19140
rect 18524 19076 18525 19140
rect 18459 19075 18525 19076
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 18462 14925 18522 19075
rect 18459 14924 18525 14925
rect 18459 14860 18460 14924
rect 18524 14860 18525 14924
rect 18459 14859 18525 14860
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17539 12068 17605 12069
rect 17539 12004 17540 12068
rect 17604 12004 17605 12068
rect 17539 12003 17605 12004
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 16803 11252 16869 11253
rect 16803 11188 16804 11252
rect 16868 11188 16869 11252
rect 16803 11187 16869 11188
rect 17944 10912 18264 11936
rect 18646 11117 18706 22339
rect 18827 19004 18893 19005
rect 18827 18940 18828 19004
rect 18892 18940 18893 19004
rect 18827 18939 18893 18940
rect 18830 15741 18890 18939
rect 18827 15740 18893 15741
rect 18827 15676 18828 15740
rect 18892 15676 18893 15740
rect 18827 15675 18893 15676
rect 19195 15332 19261 15333
rect 19195 15268 19196 15332
rect 19260 15268 19261 15332
rect 19195 15267 19261 15268
rect 19011 14924 19077 14925
rect 19011 14860 19012 14924
rect 19076 14860 19077 14924
rect 19011 14859 19077 14860
rect 18643 11116 18709 11117
rect 18643 11052 18644 11116
rect 18708 11052 18709 11116
rect 18643 11051 18709 11052
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 15699 9620 15765 9621
rect 15699 9556 15700 9620
rect 15764 9556 15765 9620
rect 15699 9555 15765 9556
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 19014 9213 19074 14859
rect 19198 11525 19258 15267
rect 19195 11524 19261 11525
rect 19195 11460 19196 11524
rect 19260 11460 19261 11524
rect 19195 11459 19261 11460
rect 19011 9212 19077 9213
rect 19011 9148 19012 9212
rect 19076 9148 19077 9212
rect 19011 9147 19077 9148
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 19566 8125 19626 23427
rect 21406 21861 21466 26419
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 23979 24036 24045 24037
rect 23979 23972 23980 24036
rect 24044 23972 24045 24036
rect 23979 23971 24045 23972
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 21955 22132 22021 22133
rect 21955 22068 21956 22132
rect 22020 22068 22021 22132
rect 21955 22067 22021 22068
rect 21403 21860 21469 21861
rect 21403 21796 21404 21860
rect 21468 21796 21469 21860
rect 21403 21795 21469 21796
rect 19931 20772 19997 20773
rect 19931 20708 19932 20772
rect 19996 20708 19997 20772
rect 19931 20707 19997 20708
rect 21219 20772 21285 20773
rect 21219 20708 21220 20772
rect 21284 20708 21285 20772
rect 21219 20707 21285 20708
rect 19934 8669 19994 20707
rect 20115 19684 20181 19685
rect 20115 19620 20116 19684
rect 20180 19620 20181 19684
rect 20115 19619 20181 19620
rect 20118 10301 20178 19619
rect 20667 19548 20733 19549
rect 20667 19484 20668 19548
rect 20732 19484 20733 19548
rect 20667 19483 20733 19484
rect 20299 19276 20365 19277
rect 20299 19212 20300 19276
rect 20364 19212 20365 19276
rect 20299 19211 20365 19212
rect 20115 10300 20181 10301
rect 20115 10236 20116 10300
rect 20180 10236 20181 10300
rect 20115 10235 20181 10236
rect 20302 9757 20362 19211
rect 20299 9756 20365 9757
rect 20299 9692 20300 9756
rect 20364 9692 20365 9756
rect 20299 9691 20365 9692
rect 20670 9621 20730 19483
rect 20851 19412 20917 19413
rect 20851 19348 20852 19412
rect 20916 19348 20917 19412
rect 20851 19347 20917 19348
rect 20854 11253 20914 19347
rect 21035 11388 21101 11389
rect 21035 11324 21036 11388
rect 21100 11324 21101 11388
rect 21035 11323 21101 11324
rect 20851 11252 20917 11253
rect 20851 11188 20852 11252
rect 20916 11188 20917 11252
rect 20851 11187 20917 11188
rect 20667 9620 20733 9621
rect 20667 9556 20668 9620
rect 20732 9556 20733 9620
rect 20667 9555 20733 9556
rect 21038 8805 21098 11323
rect 21222 9893 21282 20707
rect 21403 15604 21469 15605
rect 21403 15540 21404 15604
rect 21468 15540 21469 15604
rect 21403 15539 21469 15540
rect 21406 11797 21466 15539
rect 21958 14925 22018 22067
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22507 20636 22573 20637
rect 22507 20572 22508 20636
rect 22572 20572 22573 20636
rect 22507 20571 22573 20572
rect 22323 19412 22389 19413
rect 22323 19348 22324 19412
rect 22388 19348 22389 19412
rect 22323 19347 22389 19348
rect 22139 18596 22205 18597
rect 22139 18532 22140 18596
rect 22204 18532 22205 18596
rect 22139 18531 22205 18532
rect 22142 15469 22202 18531
rect 22326 17237 22386 19347
rect 22323 17236 22389 17237
rect 22323 17172 22324 17236
rect 22388 17172 22389 17236
rect 22323 17171 22389 17172
rect 22139 15468 22205 15469
rect 22139 15404 22140 15468
rect 22204 15404 22205 15468
rect 22139 15403 22205 15404
rect 21955 14924 22021 14925
rect 21955 14860 21956 14924
rect 22020 14860 22021 14924
rect 21955 14859 22021 14860
rect 22510 14653 22570 20571
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 23427 18732 23493 18733
rect 23427 18668 23428 18732
rect 23492 18668 23493 18732
rect 23427 18667 23493 18668
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22691 16692 22757 16693
rect 22691 16628 22692 16692
rect 22756 16628 22757 16692
rect 22691 16627 22757 16628
rect 22507 14652 22573 14653
rect 22507 14588 22508 14652
rect 22572 14588 22573 14652
rect 22507 14587 22573 14588
rect 22323 13972 22389 13973
rect 22323 13908 22324 13972
rect 22388 13908 22389 13972
rect 22323 13907 22389 13908
rect 21403 11796 21469 11797
rect 21403 11732 21404 11796
rect 21468 11732 21469 11796
rect 21403 11731 21469 11732
rect 21219 9892 21285 9893
rect 21219 9828 21220 9892
rect 21284 9828 21285 9892
rect 21219 9827 21285 9828
rect 21035 8804 21101 8805
rect 21035 8740 21036 8804
rect 21100 8740 21101 8804
rect 21035 8739 21101 8740
rect 19931 8668 19997 8669
rect 19931 8604 19932 8668
rect 19996 8604 19997 8668
rect 19931 8603 19997 8604
rect 19563 8124 19629 8125
rect 19563 8060 19564 8124
rect 19628 8060 19629 8124
rect 19563 8059 19629 8060
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 22326 5269 22386 13907
rect 22694 10573 22754 16627
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 23430 13293 23490 18667
rect 23611 18052 23677 18053
rect 23611 17988 23612 18052
rect 23676 17988 23677 18052
rect 23611 17987 23677 17988
rect 23427 13292 23493 13293
rect 23427 13228 23428 13292
rect 23492 13228 23493 13292
rect 23427 13227 23493 13228
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22691 10572 22757 10573
rect 22691 10508 22692 10572
rect 22756 10508 22757 10572
rect 22691 10507 22757 10508
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 23614 10165 23674 17987
rect 23982 10709 24042 23971
rect 24531 16692 24597 16693
rect 24531 16628 24532 16692
rect 24596 16628 24597 16692
rect 24531 16627 24597 16628
rect 24534 12341 24594 16627
rect 24715 13972 24781 13973
rect 24715 13908 24716 13972
rect 24780 13908 24781 13972
rect 24715 13907 24781 13908
rect 24531 12340 24597 12341
rect 24531 12276 24532 12340
rect 24596 12276 24597 12340
rect 24531 12275 24597 12276
rect 23979 10708 24045 10709
rect 23979 10644 23980 10708
rect 24044 10644 24045 10708
rect 23979 10643 24045 10644
rect 23611 10164 23677 10165
rect 23611 10100 23612 10164
rect 23676 10100 23677 10164
rect 23611 10099 23677 10100
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 24534 6901 24594 12275
rect 24718 6901 24778 13907
rect 24531 6900 24597 6901
rect 24531 6836 24532 6900
rect 24596 6836 24597 6900
rect 24531 6835 24597 6836
rect 24715 6900 24781 6901
rect 24715 6836 24716 6900
rect 24780 6836 24781 6900
rect 24715 6835 24781 6836
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22323 5268 22389 5269
rect 22323 5204 22324 5268
rect 22388 5204 22389 5268
rect 22323 5203 22389 5204
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 18584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1679235063
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1679235063
transform 1 0 25024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1679235063
transform 1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1679235063
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1679235063
transform 1 0 21896 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1679235063
transform 1 0 23736 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1679235063
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1679235063
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1679235063
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1679235063
transform 1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19136 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1679235063
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1679235063
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1679235063
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1679235063
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1679235063
transform 1 0 20424 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1679235063
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1679235063
transform 1 0 19136 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1679235063
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _098_
timestamp 1679235063
transform 1 0 17848 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _099_
timestamp 1679235063
transform 1 0 17388 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1679235063
transform 1 0 14812 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _101_
timestamp 1679235063
transform 1 0 16100 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1679235063
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1679235063
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _108_
timestamp 1679235063
transform 1 0 6440 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1679235063
transform 1 0 5152 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1679235063
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _115_
timestamp 1679235063
transform 1 0 6992 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _116_
timestamp 1679235063
transform 1 0 3220 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _117_
timestamp 1679235063
transform 1 0 3220 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 23736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1679235063
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _123_
timestamp 1679235063
transform 1 0 4508 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _124_
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1679235063
transform 1 0 1932 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1679235063
transform 1 0 4508 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _129_
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1679235063
transform 1 0 4048 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 7728 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 24380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 24840 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 24840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 22080 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 8372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1679235063
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1679235063
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1679235063
transform 1 0 24656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1679235063
transform 1 0 25116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1679235063
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1679235063
transform 1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1679235063
transform 1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_prog_clk_A
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_prog_clk_A
timestamp 1679235063
transform 1 0 14996 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_prog_clk_A
timestamp 1679235063
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_prog_clk_A
timestamp 1679235063
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_prog_clk_A
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_prog_clk_A
timestamp 1679235063
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_prog_clk_A
timestamp 1679235063
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold21_A
timestamp 1679235063
transform 1 0 4968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold24_A
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold27_A
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold38_A
timestamp 1679235063
transform 1 0 6440 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold39_A
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold42_A
timestamp 1679235063
transform 1 0 6440 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold46_A
timestamp 1679235063
transform 1 0 3864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold54_A
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold68_A
timestamp 1679235063
transform 1 0 3496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold69_A
timestamp 1679235063
transform 1 0 2852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold70_A
timestamp 1679235063
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1679235063
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1679235063
transform 1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 5060 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 2024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 21620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 20516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 21528 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 5428 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 2576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 21344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 5796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 20240 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 2668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 1656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 1472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 2852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 2852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 1656 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 25300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 18860 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 22172 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 20884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 3864 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 17756 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 12696 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 15272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21252 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 1472 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 1472 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 6440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 6440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_4.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 4140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 25208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_8.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_10.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 1472 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20608 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23828 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 25300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 1656 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 16192 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 13708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 2852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16008 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 15088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18860 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17112 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1679235063
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1679235063
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1679235063
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1679235063
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1679235063
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1679235063
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1679235063
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1679235063
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1679235063
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1679235063
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1679235063
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1679235063
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1679235063
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1679235063
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1679235063
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1679235063
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1679235063
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1679235063
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1679235063
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1679235063
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1679235063
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1679235063
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1679235063
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1679235063
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1679235063
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1679235063
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1679235063
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1679235063
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1679235063
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1679235063
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1679235063
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1679235063
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1679235063
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1679235063
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1679235063
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1679235063
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1679235063
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1679235063
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1679235063
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1679235063
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1679235063
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1679235063
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1679235063
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1679235063
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1679235063
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1679235063
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1679235063
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1679235063
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1679235063
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1679235063
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1679235063
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1679235063
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1679235063
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1679235063
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1679235063
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1679235063
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1679235063
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1679235063
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1679235063
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_259
timestamp 1679235063
transform 1 0 24932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1679235063
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1679235063
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1679235063
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1679235063
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1679235063
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1679235063
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1679235063
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1679235063
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1679235063
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1679235063
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1679235063
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1679235063
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1679235063
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1679235063
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1679235063
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1679235063
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1679235063
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1679235063
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1679235063
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1679235063
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1679235063
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1679235063
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1679235063
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1679235063
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1679235063
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1679235063
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1679235063
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1679235063
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1679235063
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1679235063
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1679235063
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_225
timestamp 1679235063
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1679235063
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1679235063
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1679235063
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_263
timestamp 1679235063
transform 1 0 25300 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1679235063
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1679235063
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1679235063
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1679235063
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1679235063
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1679235063
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1679235063
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1679235063
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1679235063
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1679235063
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1679235063
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1679235063
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1679235063
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1679235063
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1679235063
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1679235063
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1679235063
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1679235063
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1679235063
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1679235063
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1679235063
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1679235063
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1679235063
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1679235063
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1679235063
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1679235063
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1679235063
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1679235063
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1679235063
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1679235063
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1679235063
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1679235063
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1679235063
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1679235063
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1679235063
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1679235063
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1679235063
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_213
timestamp 1679235063
transform 1 0 20700 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_220
timestamp 1679235063
transform 1 0 21344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_226
timestamp 1679235063
transform 1 0 21896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1679235063
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_259
timestamp 1679235063
transform 1 0 24932 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1679235063
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1679235063
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1679235063
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1679235063
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1679235063
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1679235063
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1679235063
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1679235063
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1679235063
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1679235063
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1679235063
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1679235063
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1679235063
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1679235063
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1679235063
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1679235063
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1679235063
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1679235063
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1679235063
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_213
timestamp 1679235063
transform 1 0 20700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_217
timestamp 1679235063
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1679235063
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1679235063
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1679235063
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1679235063
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1679235063
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1679235063
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1679235063
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1679235063
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1679235063
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1679235063
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1679235063
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1679235063
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1679235063
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1679235063
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1679235063
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1679235063
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1679235063
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1679235063
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1679235063
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_216
timestamp 1679235063
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 1679235063
transform 1 0 21712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1679235063
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1679235063
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_255
timestamp 1679235063
transform 1 0 24564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1679235063
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1679235063
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1679235063
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1679235063
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1679235063
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1679235063
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1679235063
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1679235063
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1679235063
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1679235063
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1679235063
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1679235063
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1679235063
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_180
timestamp 1679235063
transform 1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1679235063
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_188
timestamp 1679235063
transform 1 0 18400 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1679235063
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_206
timestamp 1679235063
transform 1 0 20056 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1679235063
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1679235063
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1679235063
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1679235063
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1679235063
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1679235063
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1679235063
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1679235063
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1679235063
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1679235063
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1679235063
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1679235063
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1679235063
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1679235063
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1679235063
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1679235063
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1679235063
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1679235063
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1679235063
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1679235063
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1679235063
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp 1679235063
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1679235063
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1679235063
transform 1 0 21528 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1679235063
transform 1 0 22172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1679235063
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1679235063
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1679235063
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1679235063
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1679235063
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1679235063
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1679235063
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1679235063
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1679235063
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1679235063
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1679235063
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1679235063
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1679235063
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1679235063
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1679235063
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1679235063
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1679235063
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp 1679235063
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_199
timestamp 1679235063
transform 1 0 19412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_206
timestamp 1679235063
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1679235063
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1679235063
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1679235063
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1679235063
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1679235063
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1679235063
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1679235063
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1679235063
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1679235063
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1679235063
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1679235063
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1679235063
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_122
timestamp 1679235063
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1679235063
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1679235063
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_161
timestamp 1679235063
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1679235063
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_180
timestamp 1679235063
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_187
timestamp 1679235063
transform 1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1679235063
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1679235063
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1679235063
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1679235063
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_229
timestamp 1679235063
transform 1 0 22172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 1679235063
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1679235063
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1679235063
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1679235063
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1679235063
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1679235063
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1679235063
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1679235063
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1679235063
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1679235063
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1679235063
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1679235063
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1679235063
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_145
timestamp 1679235063
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1679235063
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_154
timestamp 1679235063
transform 1 0 15272 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1679235063
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1679235063
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_174
timestamp 1679235063
transform 1 0 17112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_181
timestamp 1679235063
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1679235063
transform 1 0 18400 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1679235063
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_202
timestamp 1679235063
transform 1 0 19688 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_206
timestamp 1679235063
transform 1 0 20056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1679235063
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1679235063
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1679235063
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1679235063
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1679235063
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1679235063
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1679235063
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1679235063
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1679235063
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1679235063
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1679235063
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1679235063
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1679235063
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1679235063
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1679235063
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_155
timestamp 1679235063
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1679235063
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_169
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_176
timestamp 1679235063
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_180
timestamp 1679235063
transform 1 0 17664 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1679235063
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1679235063
transform 1 0 18584 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1679235063
transform 1 0 19412 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1679235063
transform 1 0 19872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1679235063
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_241
timestamp 1679235063
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_245
timestamp 1679235063
transform 1 0 23644 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1679235063
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1679235063
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1679235063
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1679235063
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1679235063
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1679235063
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1679235063
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1679235063
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1679235063
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1679235063
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1679235063
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1679235063
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_125
timestamp 1679235063
transform 1 0 12604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_133
timestamp 1679235063
transform 1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1679235063
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_145
timestamp 1679235063
transform 1 0 14444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1679235063
transform 1 0 15732 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1679235063
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_171
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_174
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1679235063
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1679235063
transform 1 0 19136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1679235063
transform 1 0 19504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1679235063
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1679235063
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1679235063
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1679235063
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1679235063
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1679235063
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1679235063
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1679235063
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1679235063
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1679235063
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1679235063
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1679235063
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1679235063
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1679235063
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_148
timestamp 1679235063
transform 1 0 14720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_156
timestamp 1679235063
transform 1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1679235063
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1679235063
transform 1 0 18032 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_188
timestamp 1679235063
transform 1 0 18400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_207
timestamp 1679235063
transform 1 0 20148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1679235063
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_227
timestamp 1679235063
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_231
timestamp 1679235063
transform 1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1679235063
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1679235063
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1679235063
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1679235063
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1679235063
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1679235063
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1679235063
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1679235063
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1679235063
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1679235063
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1679235063
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_118
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1679235063
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1679235063
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1679235063
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1679235063
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1679235063
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1679235063
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_219
timestamp 1679235063
transform 1 0 21252 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1679235063
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_12
timestamp 1679235063
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1679235063
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1679235063
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1679235063
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1679235063
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1679235063
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1679235063
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1679235063
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_109
timestamp 1679235063
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1679235063
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1679235063
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1679235063
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1679235063
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1679235063
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1679235063
transform 1 0 18676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1679235063
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1679235063
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_263
timestamp 1679235063
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1679235063
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1679235063
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1679235063
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1679235063
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1679235063
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1679235063
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1679235063
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1679235063
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1679235063
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1679235063
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1679235063
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1679235063
transform 1 0 14812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1679235063
transform 1 0 15456 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1679235063
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1679235063
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1679235063
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_221
timestamp 1679235063
transform 1 0 21436 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1679235063
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1679235063
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1679235063
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_8
timestamp 1679235063
transform 1 0 1840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1679235063
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_19
timestamp 1679235063
transform 1 0 2852 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1679235063
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1679235063
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1679235063
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_66
timestamp 1679235063
transform 1 0 7176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1679235063
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1679235063
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1679235063
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1679235063
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1679235063
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_199
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1679235063
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1679235063
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1679235063
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1679235063
transform 1 0 1932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1679235063
transform 1 0 2392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_18
timestamp 1679235063
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_26
timestamp 1679235063
transform 1 0 3496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1679235063
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1679235063
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_47
timestamp 1679235063
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1679235063
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1679235063
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1679235063
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1679235063
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1679235063
transform 1 0 7912 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1679235063
transform 1 0 8648 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1679235063
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_96
timestamp 1679235063
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1679235063
transform 1 0 10580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_121
timestamp 1679235063
transform 1 0 12236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1679235063
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_161
timestamp 1679235063
transform 1 0 15916 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1679235063
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1679235063
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_210
timestamp 1679235063
transform 1 0 20424 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1679235063
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1679235063
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1679235063
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_14
timestamp 1679235063
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_35
timestamp 1679235063
transform 1 0 4324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1679235063
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1679235063
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1679235063
transform 1 0 6900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1679235063
transform 1 0 7544 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_76
timestamp 1679235063
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_92
timestamp 1679235063
transform 1 0 9568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_96
timestamp 1679235063
transform 1 0 9936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1679235063
transform 1 0 10304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1679235063
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1679235063
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1679235063
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1679235063
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1679235063
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1679235063
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_238
timestamp 1679235063
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_263
timestamp 1679235063
transform 1 0 25300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1679235063
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1679235063
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1679235063
transform 1 0 3496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1679235063
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_42
timestamp 1679235063
transform 1 0 4968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1679235063
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_49
timestamp 1679235063
transform 1 0 5612 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_69
timestamp 1679235063
transform 1 0 7452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1679235063
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1679235063
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1679235063
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_98
timestamp 1679235063
transform 1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1679235063
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_139
timestamp 1679235063
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1679235063
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1679235063
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_191
timestamp 1679235063
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1679235063
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1679235063
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1679235063
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1679235063
transform 1 0 22724 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1679235063
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1679235063
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1679235063
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_31
timestamp 1679235063
transform 1 0 3956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1679235063
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1679235063
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1679235063
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1679235063
transform 1 0 7360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1679235063
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_90
timestamp 1679235063
transform 1 0 9384 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1679235063
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1679235063
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1679235063
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1679235063
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1679235063
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1679235063
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1679235063
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1679235063
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1679235063
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1679235063
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1679235063
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1679235063
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1679235063
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1679235063
transform 1 0 2484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_33
timestamp 1679235063
transform 1 0 4140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_47
timestamp 1679235063
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_61
timestamp 1679235063
transform 1 0 6716 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1679235063
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1679235063
transform 1 0 8464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1679235063
transform 1 0 8924 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1679235063
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1679235063
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1679235063
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1679235063
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1679235063
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1679235063
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1679235063
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_263
timestamp 1679235063
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1679235063
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1679235063
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_35
timestamp 1679235063
transform 1 0 4324 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1679235063
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1679235063
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1679235063
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_72
timestamp 1679235063
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1679235063
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 1679235063
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1679235063
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1679235063
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1679235063
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1679235063
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1679235063
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_263
timestamp 1679235063
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1679235063
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_19
timestamp 1679235063
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1679235063
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_47
timestamp 1679235063
transform 1 0 5428 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1679235063
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_73
timestamp 1679235063
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1679235063
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_135
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1679235063
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1679235063
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1679235063
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1679235063
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1679235063
transform 1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1679235063
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_219
timestamp 1679235063
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1679235063
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1679235063
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1679235063
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1679235063
transform 1 0 25116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1679235063
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1679235063
transform 1 0 2484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1679235063
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_47
timestamp 1679235063
transform 1 0 5428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1679235063
transform 1 0 5796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1679235063
transform 1 0 6256 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1679235063
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_70
timestamp 1679235063
transform 1 0 7544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1679235063
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1679235063
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1679235063
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1679235063
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1679235063
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1679235063
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1679235063
transform 1 0 18676 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1679235063
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1679235063
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1679235063
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_263
timestamp 1679235063
transform 1 0 25300 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1679235063
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1679235063
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1679235063
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1679235063
transform 1 0 4324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1679235063
transform 1 0 5612 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_53
timestamp 1679235063
transform 1 0 5980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1679235063
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1679235063
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1679235063
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1679235063
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1679235063
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1679235063
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1679235063
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1679235063
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1679235063
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_265
timestamp 1679235063
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1679235063
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_12
timestamp 1679235063
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_19
timestamp 1679235063
transform 1 0 2852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1679235063
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_45
timestamp 1679235063
transform 1 0 5244 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1679235063
transform 1 0 5520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1679235063
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_70
timestamp 1679235063
transform 1 0 7544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1679235063
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1679235063
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1679235063
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1679235063
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1679235063
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1679235063
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1679235063
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1679235063
transform 1 0 19780 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_207
timestamp 1679235063
transform 1 0 20148 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1679235063
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1679235063
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1679235063
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_5
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_23
timestamp 1679235063
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_28
timestamp 1679235063
transform 1 0 3680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1679235063
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1679235063
transform 1 0 4784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 1679235063
transform 1 0 5152 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_60
timestamp 1679235063
transform 1 0 6624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_70
timestamp 1679235063
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1679235063
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1679235063
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1679235063
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1679235063
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1679235063
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1679235063
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1679235063
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1679235063
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1679235063
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1679235063
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_219
timestamp 1679235063
transform 1 0 21252 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1679235063
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1679235063
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1679235063
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_8
timestamp 1679235063
transform 1 0 1840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_34
timestamp 1679235063
transform 1 0 4232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_48
timestamp 1679235063
transform 1 0 5520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_55
timestamp 1679235063
transform 1 0 6164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1679235063
transform 1 0 6624 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1679235063
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1679235063
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1679235063
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1679235063
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1679235063
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1679235063
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_175
timestamp 1679235063
transform 1 0 17204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1679235063
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_193
timestamp 1679235063
transform 1 0 18860 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_208
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_214
timestamp 1679235063
transform 1 0 20792 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1679235063
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1679235063
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1679235063
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1679235063
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_42
timestamp 1679235063
transform 1 0 4968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1679235063
transform 1 0 6624 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_70
timestamp 1679235063
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1679235063
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1679235063
transform 1 0 11868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_128
timestamp 1679235063
transform 1 0 12880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1679235063
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_155
timestamp 1679235063
transform 1 0 15364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_159
timestamp 1679235063
transform 1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1679235063
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1679235063
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1679235063
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1679235063
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1679235063
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1679235063
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_241
timestamp 1679235063
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1679235063
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_8
timestamp 1679235063
transform 1 0 1840 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_59
timestamp 1679235063
transform 1 0 6532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_79
timestamp 1679235063
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1679235063
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_104
timestamp 1679235063
transform 1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_108
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1679235063
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1679235063
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1679235063
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_155
timestamp 1679235063
transform 1 0 15364 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1679235063
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1679235063
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1679235063
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1679235063
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1679235063
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1679235063
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1679235063
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1679235063
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1679235063
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1679235063
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1679235063
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1679235063
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1679235063
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_130
timestamp 1679235063
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1679235063
transform 1 0 13616 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1679235063
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1679235063
transform 1 0 15824 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_171
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1679235063
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1679235063
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1679235063
transform 1 0 21252 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1679235063
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1679235063
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_8
timestamp 1679235063
transform 1 0 1840 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1679235063
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_42
timestamp 1679235063
transform 1 0 4968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_89
timestamp 1679235063
transform 1 0 9292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1679235063
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1679235063
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_128
timestamp 1679235063
transform 1 0 12880 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1679235063
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1679235063
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1679235063
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1679235063
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1679235063
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_207
timestamp 1679235063
transform 1 0 20148 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1679235063
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1679235063
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_63
timestamp 1679235063
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_68
timestamp 1679235063
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1679235063
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1679235063
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1679235063
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1679235063
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1679235063
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1679235063
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_217
timestamp 1679235063
transform 1 0 21068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1679235063
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1679235063
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_240
timestamp 1679235063
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1679235063
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1679235063
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_8
timestamp 1679235063
transform 1 0 1840 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1679235063
transform 1 0 4048 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1679235063
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1679235063
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1679235063
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1679235063
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1679235063
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1679235063
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_184
timestamp 1679235063
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1679235063
transform 1 0 18768 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1679235063
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1679235063
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_60
timestamp 1679235063
transform 1 0 6624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1679235063
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_117
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_135
timestamp 1679235063
transform 1 0 13524 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_139
timestamp 1679235063
transform 1 0 13892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_150
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1679235063
transform 1 0 15364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1679235063
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1679235063
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_205
timestamp 1679235063
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_218
timestamp 1679235063
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_227
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_250
timestamp 1679235063
transform 1 0 24104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1679235063
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_151
timestamp 1679235063
transform 1 0 14996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_163
timestamp 1679235063
transform 1 0 16100 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_167
timestamp 1679235063
transform 1 0 16468 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_179
timestamp 1679235063
transform 1 0 17572 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_183
timestamp 1679235063
transform 1 0 17940 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6808 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20516 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold3
timestamp 1679235063
transform 1 0 1656 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 15640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5
timestamp 1679235063
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1679235063
transform 1 0 20516 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold8
timestamp 1679235063
transform 1 0 24564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold10
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 18400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold13
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold14
timestamp 1679235063
transform 1 0 6808 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 21896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold16
timestamp 1679235063
transform 1 0 7912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold18
timestamp 1679235063
transform 1 0 14260 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold19
timestamp 1679235063
transform 1 0 23000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1679235063
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1679235063
transform 1 0 1656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold27
timestamp 1679235063
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 4232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 10488 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1679235063
transform 1 0 6808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1679235063
transform 1 0 7820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1679235063
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 17940 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1679235063
transform 1 0 5704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold39
timestamp 1679235063
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 11868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold42
timestamp 1679235063
transform 1 0 6808 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1679235063
transform 1 0 12880 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1679235063
transform 1 0 15364 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 24196 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold52
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold53
timestamp 1679235063
transform 1 0 20240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1679235063
transform 1 0 6716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 9292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 17296 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 21436 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1679235063
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 9292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 16928 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold68
timestamp 1679235063
transform 1 0 4600 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold69
timestamp 1679235063
transform 1 0 1656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold70
timestamp 1679235063
transform 1 0 11960 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold71
timestamp 1679235063
transform 1 0 24196 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1679235063
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1679235063
transform 1 0 4048 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1679235063
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1679235063
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1679235063
transform 1 0 2576 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1679235063
transform 1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 8648 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1679235063
transform 1 0 16376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1679235063
transform 1 0 6624 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1679235063
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1679235063
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1679235063
transform 1 0 18768 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1679235063
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1679235063
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1679235063
transform 1 0 15088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1679235063
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1679235063
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1679235063
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 18032 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 9200 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 9660 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1679235063
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1679235063
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1679235063
transform 1 0 7268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1679235063
transform 1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1679235063
transform 1 0 2576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 20516 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1679235063
transform 1 0 4508 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 5796 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1679235063
transform 1 0 5336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1679235063
transform 1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1679235063
transform 1 0 4508 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1679235063
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 19412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1679235063
transform 1 0 4692 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 2576 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 3220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1679235063
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 5980 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1679235063
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1679235063
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1679235063
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1679235063
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1679235063
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1679235063
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1679235063
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1679235063
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1679235063
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1679235063
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1679235063
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1679235063
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1679235063
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1679235063
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22172 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23276 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22816 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21344 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18032 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9016 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10488 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__151 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19596 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__157
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__126
timestamp 1679235063
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 22540 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__131
timestamp 1679235063
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__132
timestamp 1679235063
transform 1 0 5888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__152
timestamp 1679235063
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20424 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__124
timestamp 1679235063
transform 1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__125
timestamp 1679235063
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__127
timestamp 1679235063
transform 1 0 17940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__128
timestamp 1679235063
transform 1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__129
timestamp 1679235063
transform 1 0 21252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20424 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__130
timestamp 1679235063
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__133
timestamp 1679235063
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__139
timestamp 1679235063
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20240 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__144
timestamp 1679235063
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 20332 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__149
timestamp 1679235063
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__150
timestamp 1679235063
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__134
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13800 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9292 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__135
timestamp 1679235063
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16468 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__136
timestamp 1679235063
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4508 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9476 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__137
timestamp 1679235063
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__138
timestamp 1679235063
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__140
timestamp 1679235063
transform 1 0 3956 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__141
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__142
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__143
timestamp 1679235063
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__145
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6440 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__146
timestamp 1679235063
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__147
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10396 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__148
timestamp 1679235063
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal2 6762 1571 6762 1571 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal1 19412 12750 19412 12750 0 chanx_right_in[0]
rlabel metal1 16744 15606 16744 15606 0 chanx_right_in[10]
rlabel metal3 18446 17544 18446 17544 0 chanx_right_in[11]
rlabel metal2 16514 18037 16514 18037 0 chanx_right_in[12]
rlabel metal2 2162 18785 2162 18785 0 chanx_right_in[13]
rlabel metal1 14950 14280 14950 14280 0 chanx_right_in[14]
rlabel metal2 23414 19023 23414 19023 0 chanx_right_in[15]
rlabel metal3 5451 10676 5451 10676 0 chanx_right_in[16]
rlabel metal1 4186 15334 4186 15334 0 chanx_right_in[17]
rlabel metal2 12558 11628 12558 11628 0 chanx_right_in[18]
rlabel metal2 21758 22984 21758 22984 0 chanx_right_in[19]
rlabel metal1 19826 10540 19826 10540 0 chanx_right_in[1]
rlabel metal2 22494 23885 22494 23885 0 chanx_right_in[20]
rlabel metal1 6578 17646 6578 17646 0 chanx_right_in[21]
rlabel metal1 2392 22202 2392 22202 0 chanx_right_in[22]
rlabel metal3 26228 22372 26228 22372 0 chanx_right_in[23]
rlabel metal3 21367 19380 21367 19380 0 chanx_right_in[24]
rlabel metal2 26220 23188 26220 23188 0 chanx_right_in[25]
rlabel metal2 26266 23596 26266 23596 0 chanx_right_in[26]
rlabel metal3 25193 24004 25193 24004 0 chanx_right_in[27]
rlabel metal2 26128 22508 26128 22508 0 chanx_right_in[28]
rlabel metal2 22126 24565 22126 24565 0 chanx_right_in[29]
rlabel metal2 22632 12716 22632 12716 0 chanx_right_in[2]
rlabel metal1 21206 13872 21206 13872 0 chanx_right_in[3]
rlabel metal1 19872 9962 19872 9962 0 chanx_right_in[4]
rlabel metal1 16468 11050 16468 11050 0 chanx_right_in[5]
rlabel metal1 20378 8058 20378 8058 0 chanx_right_in[6]
rlabel metal3 10833 12172 10833 12172 0 chanx_right_in[7]
rlabel metal3 17204 16184 17204 16184 0 chanx_right_in[8]
rlabel metal1 20148 14790 20148 14790 0 chanx_right_in[9]
rlabel metal3 25722 748 25722 748 0 chanx_right_out[0]
rlabel metal1 24104 5270 24104 5270 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24426 6766 24426 6766 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal2 24794 6953 24794 6953 0 chanx_right_out[17]
rlabel metal1 24380 7922 24380 7922 0 chanx_right_out[18]
rlabel metal1 24012 8398 24012 8398 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 25162 8177 25162 8177 0 chanx_right_out[20]
rlabel metal1 24380 9010 24380 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal2 24794 9265 24794 9265 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 25162 10285 25162 10285 0 chanx_right_out[25]
rlabel metal1 24380 11186 24380 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24794 11373 24794 11373 0 chanx_right_out[28]
rlabel metal3 25768 12580 25768 12580 0 chanx_right_out[29]
rlabel metal3 24296 1564 24296 1564 0 chanx_right_out[2]
rlabel metal1 20792 2618 20792 2618 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25676 3196 25676 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal2 25162 3553 25162 3553 0 chanx_right_out[8]
rlabel metal3 25952 4420 25952 4420 0 chanx_right_out[9]
rlabel metal1 6026 14042 6026 14042 0 chany_top_in[0]
rlabel metal1 8970 20910 8970 20910 0 chany_top_in[10]
rlabel metal2 16790 25833 16790 25833 0 chany_top_in[11]
rlabel metal2 17158 25969 17158 25969 0 chany_top_in[12]
rlabel metal3 15111 23188 15111 23188 0 chany_top_in[13]
rlabel metal2 21758 8092 21758 8092 0 chany_top_in[14]
rlabel metal2 17986 26265 17986 26265 0 chany_top_in[15]
rlabel metal2 18630 25901 18630 25901 0 chany_top_in[16]
rlabel metal2 18998 26037 18998 26037 0 chany_top_in[17]
rlabel metal2 19366 26173 19366 26173 0 chany_top_in[18]
rlabel metal2 3082 18428 3082 18428 0 chany_top_in[19]
rlabel metal2 12834 24616 12834 24616 0 chany_top_in[1]
rlabel metal2 19826 26231 19826 26231 0 chany_top_in[20]
rlabel metal2 2346 14433 2346 14433 0 chany_top_in[21]
rlabel metal2 20746 26248 20746 26248 0 chany_top_in[22]
rlabel via3 21229 20740 21229 20740 0 chany_top_in[23]
rlabel metal2 21429 26724 21429 26724 0 chany_top_in[24]
rlabel metal1 20332 9486 20332 9486 0 chany_top_in[25]
rlabel metal2 22310 25612 22310 25612 0 chany_top_in[26]
rlabel via1 22402 26333 22402 26333 0 chany_top_in[27]
rlabel metal1 2622 16694 2622 16694 0 chany_top_in[28]
rlabel metal1 19182 8942 19182 8942 0 chany_top_in[29]
rlabel metal3 12604 12240 12604 12240 0 chany_top_in[2]
rlabel metal1 13754 23120 13754 23120 0 chany_top_in[3]
rlabel metal2 12466 15946 12466 15946 0 chany_top_in[4]
rlabel metal3 14329 23460 14329 23460 0 chany_top_in[5]
rlabel via2 2162 12835 2162 12835 0 chany_top_in[6]
rlabel metal2 19642 24276 19642 24276 0 chany_top_in[7]
rlabel via2 2346 13923 2346 13923 0 chany_top_in[8]
rlabel metal2 15778 15079 15778 15079 0 chany_top_in[9]
rlabel metal1 1978 19278 1978 19278 0 chany_top_out[0]
rlabel metal1 4692 23766 4692 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4876 24242 4876 24242 0 chany_top_out[13]
rlabel metal1 7130 20978 7130 20978 0 chany_top_out[14]
rlabel metal1 7590 21454 7590 21454 0 chany_top_out[15]
rlabel metal1 6716 23630 6716 23630 0 chany_top_out[16]
rlabel metal1 7130 23154 7130 23154 0 chany_top_out[17]
rlabel metal2 8326 24184 8326 24184 0 chany_top_out[18]
rlabel metal1 7268 24106 7268 24106 0 chany_top_out[19]
rlabel metal1 2438 19890 2438 19890 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8832 23154 8832 23154 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9660 23766 9660 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal2 10994 24242 10994 24242 0 chany_top_out[26]
rlabel metal2 12650 23120 12650 23120 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel metal1 12627 24242 12627 24242 0 chany_top_out[29]
rlabel metal2 2438 23606 2438 23606 0 chany_top_out[2]
rlabel metal1 3082 20366 3082 20366 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4416 23290 4416 23290 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3956 23154 3956 23154 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal2 21574 20944 21574 20944 0 clknet_0_prog_clk
rlabel metal1 10488 13158 10488 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15640 15538 15640 15538 0 clknet_3_1__leaf_prog_clk
rlabel via1 9062 20978 9062 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 13570 20468 13570 20468 0 clknet_3_3__leaf_prog_clk
rlabel metal1 19504 14042 19504 14042 0 clknet_3_4__leaf_prog_clk
rlabel metal1 20838 13362 20838 13362 0 clknet_3_5__leaf_prog_clk
rlabel metal1 19826 18734 19826 18734 0 clknet_3_6__leaf_prog_clk
rlabel metal2 23322 22848 23322 22848 0 clknet_3_7__leaf_prog_clk
rlabel metal2 6854 5746 6854 5746 0 net1
rlabel metal2 2714 17272 2714 17272 0 net10
rlabel metal1 3542 15946 3542 15946 0 net100
rlabel metal1 12006 19278 12006 19278 0 net101
rlabel metal2 17250 18020 17250 18020 0 net102
rlabel metal1 23920 22066 23920 22066 0 net103
rlabel metal1 4830 24106 4830 24106 0 net104
rlabel metal2 2162 23001 2162 23001 0 net105
rlabel metal1 5152 16422 5152 16422 0 net106
rlabel metal1 4922 17170 4922 17170 0 net107
rlabel metal1 1886 17782 1886 17782 0 net108
rlabel metal1 4738 18802 4738 18802 0 net109
rlabel metal1 9568 23018 9568 23018 0 net11
rlabel metal2 10074 18938 10074 18938 0 net110
rlabel metal2 2070 20519 2070 20519 0 net111
rlabel metal1 4646 17714 4646 17714 0 net112
rlabel metal2 1886 21284 1886 21284 0 net113
rlabel metal3 7199 14756 7199 14756 0 net114
rlabel metal1 4232 14586 4232 14586 0 net115
rlabel metal1 2300 20910 2300 20910 0 net116
rlabel metal4 12604 20264 12604 20264 0 net117
rlabel metal1 2392 21998 2392 21998 0 net118
rlabel metal1 2990 21556 2990 21556 0 net119
rlabel metal1 15226 19686 15226 19686 0 net12
rlabel metal1 4094 20842 4094 20842 0 net120
rlabel metal1 5428 16626 5428 16626 0 net121
rlabel metal2 2254 22916 2254 22916 0 net122
rlabel metal2 18630 24276 18630 24276 0 net123
rlabel metal2 20838 10013 20838 10013 0 net124
rlabel metal3 20470 13804 20470 13804 0 net125
rlabel metal1 25898 23018 25898 23018 0 net126
rlabel metal1 17710 10098 17710 10098 0 net127
rlabel metal1 19044 12818 19044 12818 0 net128
rlabel metal1 20976 7854 20976 7854 0 net129
rlabel metal2 12880 20298 12880 20298 0 net13
rlabel metal2 23414 8874 23414 8874 0 net130
rlabel metal3 15801 16796 15801 16796 0 net131
rlabel metal3 17204 18360 17204 18360 0 net132
rlabel metal1 19918 19686 19918 19686 0 net133
rlabel metal2 14214 21869 14214 21869 0 net134
rlabel metal1 12650 21488 12650 21488 0 net135
rlabel metal1 1564 15130 1564 15130 0 net136
rlabel metal1 8648 14382 8648 14382 0 net137
rlabel metal1 8418 15572 8418 15572 0 net138
rlabel metal1 23736 22950 23736 22950 0 net139
rlabel metal2 15594 18649 15594 18649 0 net14
rlabel metal1 6716 13226 6716 13226 0 net140
rlabel metal1 12558 20502 12558 20502 0 net141
rlabel metal2 12190 19856 12190 19856 0 net142
rlabel metal1 4692 14042 4692 14042 0 net143
rlabel metal1 18768 13362 18768 13362 0 net144
rlabel metal1 10212 16082 10212 16082 0 net145
rlabel metal1 13524 15470 13524 15470 0 net146
rlabel metal1 14306 16048 14306 16048 0 net147
rlabel metal1 15272 19346 15272 19346 0 net148
rlabel metal1 20792 23834 20792 23834 0 net149
rlabel metal2 16882 19669 16882 19669 0 net15
rlabel via2 13846 23477 13846 23477 0 net150
rlabel metal1 20884 19414 20884 19414 0 net151
rlabel via2 14306 17731 14306 17731 0 net152
rlabel metal2 1978 11849 1978 11849 0 net153
rlabel metal1 13478 13464 13478 13464 0 net154
rlabel metal1 23644 14246 23644 14246 0 net155
rlabel metal1 25438 13226 25438 13226 0 net156
rlabel metal1 5198 19890 5198 19890 0 net157
rlabel metal1 19320 13906 19320 13906 0 net158
rlabel metal1 21206 15402 21206 15402 0 net159
rlabel metal1 2024 16422 2024 16422 0 net16
rlabel metal1 13846 23800 13846 23800 0 net160
rlabel metal2 21206 11458 21206 11458 0 net161
rlabel via2 1610 23035 1610 23035 0 net162
rlabel metal2 16330 11696 16330 11696 0 net163
rlabel metal2 21482 11628 21482 11628 0 net164
rlabel metal1 15134 17306 15134 17306 0 net165
rlabel metal2 17250 16422 17250 16422 0 net166
rlabel metal2 19734 16830 19734 16830 0 net167
rlabel metal2 8602 20672 8602 20672 0 net168
rlabel metal1 25254 12954 25254 12954 0 net169
rlabel metal2 17940 21862 17940 21862 0 net17
rlabel metal2 19090 11220 19090 11220 0 net170
rlabel metal2 20286 18989 20286 18989 0 net171
rlabel metal1 21666 16150 21666 16150 0 net172
rlabel via2 19734 20859 19734 20859 0 net173
rlabel metal1 19642 15096 19642 15096 0 net174
rlabel metal2 16514 20944 16514 20944 0 net175
rlabel metal1 21022 14892 21022 14892 0 net176
rlabel metal2 14030 17068 14030 17068 0 net177
rlabel metal2 19182 16150 19182 16150 0 net178
rlabel metal2 13110 11934 13110 11934 0 net179
rlabel via3 19941 20740 19941 20740 0 net18
rlabel metal2 16790 11169 16790 11169 0 net180
rlabel metal1 11178 16150 11178 16150 0 net181
rlabel metal1 6486 20570 6486 20570 0 net182
rlabel metal1 18170 23596 18170 23596 0 net183
rlabel metal1 24794 13294 24794 13294 0 net184
rlabel metal1 8924 18326 8924 18326 0 net185
rlabel metal2 22126 23817 22126 23817 0 net186
rlabel metal1 7406 20366 7406 20366 0 net187
rlabel metal2 10994 14620 10994 14620 0 net188
rlabel metal3 12788 23460 12788 23460 0 net189
rlabel via2 19458 8075 19458 8075 0 net19
rlabel metal2 14582 14620 14582 14620 0 net190
rlabel metal1 10028 17578 10028 17578 0 net191
rlabel metal1 14759 22202 14759 22202 0 net192
rlabel metal1 23736 14926 23736 14926 0 net193
rlabel metal1 13386 19278 13386 19278 0 net194
rlabel metal1 18446 12342 18446 12342 0 net195
rlabel metal2 25254 10132 25254 10132 0 net196
rlabel metal3 17204 13056 17204 13056 0 net197
rlabel metal2 20010 23494 20010 23494 0 net198
rlabel metal1 16284 18802 16284 18802 0 net199
rlabel metal1 17802 6630 17802 6630 0 net2
rlabel metal2 18814 10251 18814 10251 0 net20
rlabel metal2 12098 13090 12098 13090 0 net200
rlabel metal1 20746 20026 20746 20026 0 net201
rlabel metal1 11822 17578 11822 17578 0 net202
rlabel metal2 12282 14552 12282 14552 0 net203
rlabel metal1 15456 15130 15456 15130 0 net204
rlabel metal1 6716 21046 6716 21046 0 net205
rlabel metal1 14490 20366 14490 20366 0 net206
rlabel metal2 12098 15062 12098 15062 0 net207
rlabel metal1 14444 22542 14444 22542 0 net208
rlabel metal1 14168 13226 14168 13226 0 net209
rlabel metal3 20585 19652 20585 19652 0 net21
rlabel metal2 20010 13090 20010 13090 0 net210
rlabel metal2 11040 23324 11040 23324 0 net211
rlabel metal1 22678 17102 22678 17102 0 net212
rlabel metal1 22264 23834 22264 23834 0 net213
rlabel metal1 10948 19754 10948 19754 0 net214
rlabel metal1 17572 13362 17572 13362 0 net215
rlabel metal1 20056 11254 20056 11254 0 net216
rlabel metal2 21666 9554 21666 9554 0 net217
rlabel metal1 15870 12886 15870 12886 0 net218
rlabel metal1 8970 19414 8970 19414 0 net219
rlabel metal3 16629 19380 16629 19380 0 net22
rlabel metal1 21344 10778 21344 10778 0 net220
rlabel metal1 25162 11322 25162 11322 0 net221
rlabel metal1 17572 10778 17572 10778 0 net222
rlabel metal1 9752 16218 9752 16218 0 net223
rlabel metal1 17434 23494 17434 23494 0 net224
rlabel metal1 8602 21590 8602 21590 0 net225
rlabel metal1 12006 17272 12006 17272 0 net226
rlabel metal2 23506 23834 23506 23834 0 net227
rlabel via2 17158 22661 17158 22661 0 net228
rlabel metal1 14536 16490 14536 16490 0 net229
rlabel metal1 14996 10234 14996 10234 0 net23
rlabel metal2 17342 18836 17342 18836 0 net230
rlabel metal1 18998 4794 18998 4794 0 net24
rlabel metal1 17112 17646 17112 17646 0 net25
rlabel metal1 19688 16082 19688 16082 0 net26
rlabel metal3 16146 13804 16146 13804 0 net27
rlabel metal1 16974 9146 16974 9146 0 net28
rlabel metal2 12558 18717 12558 18717 0 net29
rlabel metal1 17618 16422 17618 16422 0 net3
rlabel metal2 13662 21954 13662 21954 0 net30
rlabel metal1 19136 14586 19136 14586 0 net31
rlabel metal3 7705 12172 7705 12172 0 net32
rlabel metal2 15226 14569 15226 14569 0 net33
rlabel metal1 21528 12750 21528 12750 0 net34
rlabel metal2 6762 14943 6762 14943 0 net35
rlabel metal1 19320 18190 19320 18190 0 net36
rlabel metal3 20815 19516 20815 19516 0 net37
rlabel via2 1886 16099 1886 16099 0 net38
rlabel metal1 20930 18156 20930 18156 0 net39
rlabel via2 15870 17323 15870 17323 0 net4
rlabel metal2 15134 15011 15134 15011 0 net40
rlabel metal2 19366 18751 19366 18751 0 net41
rlabel metal2 1886 17375 1886 17375 0 net42
rlabel metal2 11730 10846 11730 10846 0 net43
rlabel metal2 5382 14399 5382 14399 0 net44
rlabel metal2 20010 14688 20010 14688 0 net45
rlabel metal2 23644 23052 23644 23052 0 net46
rlabel metal1 19642 9418 19642 9418 0 net47
rlabel metal2 17066 15572 17066 15572 0 net48
rlabel metal2 19366 9197 19366 9197 0 net49
rlabel metal2 17250 18207 17250 18207 0 net5
rlabel metal1 23644 23834 23644 23834 0 net50
rlabel metal1 25070 24310 25070 24310 0 net51
rlabel metal1 9384 12342 9384 12342 0 net52
rlabel metal2 22494 22321 22494 22321 0 net53
rlabel metal2 21758 11237 21758 11237 0 net54
rlabel metal3 17756 22712 17756 22712 0 net55
rlabel metal2 17250 6528 17250 6528 0 net56
rlabel metal2 16422 15181 16422 15181 0 net57
rlabel metal1 1978 12920 1978 12920 0 net58
rlabel metal1 18860 18666 18860 18666 0 net59
rlabel metal1 1978 18632 1978 18632 0 net6
rlabel metal1 2162 14008 2162 14008 0 net60
rlabel metal1 11707 10098 11707 10098 0 net61
rlabel metal2 1518 18088 1518 18088 0 net62
rlabel metal1 20286 2482 20286 2482 0 net63
rlabel metal2 20102 7038 20102 7038 0 net64
rlabel via2 22310 5219 22310 5219 0 net65
rlabel metal2 23736 13668 23736 13668 0 net66
rlabel metal1 22862 5610 22862 5610 0 net67
rlabel metal2 22218 7004 22218 7004 0 net68
rlabel metal1 19458 7412 19458 7412 0 net69
rlabel metal1 11592 14042 11592 14042 0 net7
rlabel metal1 21390 6732 21390 6732 0 net70
rlabel metal1 16284 13838 16284 13838 0 net71
rlabel metal2 23598 14348 23598 14348 0 net72
rlabel metal2 22402 8602 22402 8602 0 net73
rlabel metal1 25898 17034 25898 17034 0 net74
rlabel metal1 21482 3502 21482 3502 0 net75
rlabel metal2 23506 6766 23506 6766 0 net76
rlabel metal2 22678 8228 22678 8228 0 net77
rlabel metal1 20516 9146 20516 9146 0 net78
rlabel metal1 19182 8568 19182 8568 0 net79
rlabel metal1 10258 14518 10258 14518 0 net8
rlabel metal2 21574 10268 21574 10268 0 net80
rlabel metal1 20746 6868 20746 6868 0 net81
rlabel metal2 18906 9962 18906 9962 0 net82
rlabel metal1 17710 7956 17710 7956 0 net83
rlabel metal1 15134 10676 15134 10676 0 net84
rlabel metal2 21850 11322 21850 11322 0 net85
rlabel metal1 20700 4114 20700 4114 0 net86
rlabel metal1 18446 3060 18446 3060 0 net87
rlabel metal1 22862 2346 22862 2346 0 net88
rlabel metal2 22310 3196 22310 3196 0 net89
rlabel metal2 16514 17323 16514 17323 0 net9
rlabel metal1 23782 3502 23782 3502 0 net90
rlabel metal2 22126 5372 22126 5372 0 net91
rlabel metal2 23966 6460 23966 6460 0 net92
rlabel metal1 22862 4624 22862 4624 0 net93
rlabel metal1 1978 19380 1978 19380 0 net94
rlabel metal3 19067 21692 19067 21692 0 net95
rlabel metal1 19044 21454 19044 21454 0 net96
rlabel metal2 2622 20468 2622 20468 0 net97
rlabel metal3 4416 21964 4416 21964 0 net98
rlabel metal1 5267 17306 5267 17306 0 net99
rlabel metal2 18998 15606 18998 15606 0 prog_clk
rlabel metal2 24518 24677 24518 24677 0 prog_reset
rlabel metal2 1518 19754 1518 19754 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 24886 23766 24886 23766 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 25998 26044 25998 26044 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 26090 26452 26090 26452 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 14536 17170 14536 17170 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal1 20056 19278 20056 19278 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal1 17618 21420 17618 21420 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel via2 16514 11611 16514 11611 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal1 14858 16082 14858 16082 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal2 20286 10234 20286 10234 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 20838 10608 20838 10608 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal2 21482 19975 21482 19975 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 24058 16218 24058 16218 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22494 17714 22494 17714 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 24564 13838 24564 13838 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24564 14926 24564 14926 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal2 23782 13056 23782 13056 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal2 19734 10812 19734 10812 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal1 1748 21522 1748 21522 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 22586 22508 22586 22508 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 21528 13838 21528 13838 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 23828 13498 23828 13498 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 21482 16456 21482 16456 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 23874 16082 23874 16082 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal1 20240 15538 20240 15538 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal1 20792 17102 20792 17102 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal1 20010 14484 20010 14484 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal1 18722 15504 18722 15504 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal2 24058 23341 24058 23341 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal1 23092 22950 23092 22950 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17158 13498 17158 13498 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18446 14586 18446 14586 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 19136 12682 19136 12682 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 18124 18802 18124 18802 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20700 12682 20700 12682 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal1 19182 11866 19182 11866 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal1 21160 11526 21160 11526 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 25254 22474 25254 22474 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 23368 22134 23368 22134 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 25162 23596 25162 23596 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15824 19278 15824 19278 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal1 11868 9146 11868 9146 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 15088 23630 15088 23630 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 14904 21454 14904 21454 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal2 16054 22916 16054 22916 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 7866 20502 7866 20502 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal1 14536 19482 14536 19482 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal2 12006 21080 12006 21080 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal1 16790 22066 16790 22066 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 9246 22066 9246 22066 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal1 13570 22712 13570 22712 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 10626 19142 10626 19142 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 7958 20026 7958 20026 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 18722 20519 18722 20519 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal2 17342 20366 17342 20366 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 9982 18802 9982 18802 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal2 9338 17238 9338 17238 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12650 19108 12650 19108 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel metal2 14214 19737 14214 19737 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 11546 16490 11546 16490 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 14398 20910 14398 20910 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 11408 15334 11408 15334 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal1 13524 15878 13524 15878 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 20976 23222 20976 23222 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal3 20263 19108 20263 19108 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 11086 15572 11086 15572 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal1 13110 14518 13110 14518 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 13432 12206 13432 12206 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 13800 13498 13800 13498 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14214 14518 14214 14518 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 17250 13158 17250 13158 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16146 14994 16146 14994 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 17066 23154 17066 23154 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal1 1702 22644 1702 22644 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal2 16790 22746 16790 22746 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 10166 9044 10166 9044 0 sb_0__0_.mux_right_track_0.out
rlabel metal1 19136 19346 19136 19346 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 19482 20056 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal4 18492 17000 18492 17000 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15502 10234 15502 10234 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 24196 21862 24196 21862 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 23023 16660 23023 16660 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19228 8466 19228 8466 0 sb_0__0_.mux_right_track_12.out
rlabel metal1 22494 15980 22494 15980 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 19941 15300 19941 15300 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19642 9316 19642 9316 0 sb_0__0_.mux_right_track_14.out
rlabel metal2 23874 18224 23874 18224 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16882 12614 16882 12614 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 18722 8228 18722 8228 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 23690 14450 23690 14450 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23092 14246 23092 14246 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20562 6290 20562 6290 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 25208 13158 25208 13158 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20654 8432 20654 8432 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14490 10404 14490 10404 0 sb_0__0_.mux_right_track_2.out
rlabel metal1 22448 22406 22448 22406 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14720 9690 14720 9690 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 6766 20470 6766 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 21160 14042 21160 14042 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 7378 20792 7378 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19182 7412 19182 7412 0 sb_0__0_.mux_right_track_30.out
rlabel metal1 21252 15538 21252 15538 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 15334 21160 15334 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18446 8330 18446 8330 0 sb_0__0_.mux_right_track_32.out
rlabel metal2 20010 18428 20010 18428 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19366 15334 19366 15334 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25070 6426 25070 6426 0 sb_0__0_.mux_right_track_34.out
rlabel metal1 19872 14450 19872 14450 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19412 14246 19412 14246 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 18998 13396 18998 13396 0 sb_0__0_.mux_right_track_4.out
rlabel metal1 24840 20026 24840 20026 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24288 22950 24288 22950 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21942 6698 21942 6698 0 sb_0__0_.mux_right_track_44.out
rlabel metal2 17526 16048 17526 16048 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17066 11662 17066 11662 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 5202 23414 5202 0 sb_0__0_.mux_right_track_46.out
rlabel metal2 18630 13515 18630 13515 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18814 12070 18814 12070 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 5576 20470 5576 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20332 12886 20332 12886 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19918 12614 19918 12614 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 2414 24702 2414 0 sb_0__0_.mux_right_track_50.out
rlabel metal2 20562 15742 20562 15742 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21781 5202 21781 5202 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17664 7514 17664 7514 0 sb_0__0_.mux_right_track_6.out
rlabel metal1 24748 24038 24748 24038 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22540 21862 22540 21862 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18170 7514 18170 7514 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21298 6596 21298 6596 0 sb_0__0_.mux_right_track_8.out
rlabel metal1 24886 23494 24886 23494 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25070 18870 25070 18870 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4048 24038 4048 24038 0 sb_0__0_.mux_top_track_0.out
rlabel metal2 14306 19176 14306 19176 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17388 19482 17388 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 19482 14858 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7958 14586 7958 14586 0 sb_0__0_.mux_top_track_10.out
rlabel metal2 17710 21760 17710 21760 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14122 15215 14122 15215 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 4002 19516 4002 19516 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 15456 21114 15456 21114 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12282 20842 12282 20842 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2185 17646 2185 17646 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 15456 21862 15456 21862 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7222 19482 7222 19482 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5198 15130 5198 15130 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 15502 21012 15502 21012 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9476 21862 9476 21862 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 4738 16116 4738 16116 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 10902 19958 10902 19958 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 2162 15436 2162 15436 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3910 14926 3910 14926 0 sb_0__0_.mux_top_track_2.out
rlabel via2 20838 21131 20838 21131 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17756 21114 17756 21114 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3358 16082 3358 16082 0 sb_0__0_.mux_top_track_28.out
rlabel metal1 15180 18394 15180 18394 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3634 18326 3634 18326 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4692 14586 4692 14586 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 16606 20026 16606 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4922 15045 4922 15045 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3910 13804 3910 13804 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 16836 18054 16836 18054 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 4554 13906 4554 13906 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5980 15674 5980 15674 0 sb_0__0_.mux_top_track_34.out
rlabel metal2 14122 16864 14122 16864 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 6026 15980 6026 15980 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4094 13702 4094 13702 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 19918 22746 19918 22746 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 23885 12466 23885 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 6486 16184 6486 16184 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 13386 15912 13386 15912 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 6670 15708 6670 15708 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4600 13498 4600 13498 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13202 15606 13202 15606 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12742 14042 12742 14042 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8556 20774 8556 20774 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 16882 16218 16882 16218 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12604 16218 12604 16218 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5014 12818 5014 12818 0 sb_0__0_.mux_top_track_50.out
rlabel metal1 15318 17850 15318 17850 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8786 18836 8786 18836 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7084 14042 7084 14042 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 15456 21318 15456 21318 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17618 23460 17618 23460 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15686 15385 15686 15385 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 2346 15130 2346 15130 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 18768 22474 18768 22474 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14122 24327 14122 24327 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18032 20774 18032 20774 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 17526 17170 17526 17170 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 1610 22066 1610 22066 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 15410 21454 15410 21454 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
