magic
tech sky130A
magscale 1 2
timestamp 1681041005
<< viali >>
rect 3985 54281 4019 54315
rect 14565 54281 14599 54315
rect 16405 54281 16439 54315
rect 24501 54281 24535 54315
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 14105 54213 14139 54247
rect 18429 54213 18463 54247
rect 21465 54213 21499 54247
rect 23305 54213 23339 54247
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 11897 54145 11931 54179
rect 12357 54145 12391 54179
rect 14841 54145 14875 54179
rect 15577 54145 15611 54179
rect 16129 54145 16163 54179
rect 16865 54145 16899 54179
rect 17601 54145 17635 54179
rect 18981 54145 19015 54179
rect 19441 54145 19475 54179
rect 20177 54145 20211 54179
rect 20913 54145 20947 54179
rect 22017 54145 22051 54179
rect 22753 54145 22787 54179
rect 23765 54145 23799 54179
rect 24961 54145 24995 54179
rect 3249 54077 3283 54111
rect 12817 54077 12851 54111
rect 17785 54009 17819 54043
rect 3801 53941 3835 53975
rect 11713 53941 11747 53975
rect 15025 53941 15059 53975
rect 15761 53941 15795 53975
rect 17049 53941 17083 53975
rect 18521 53941 18555 53975
rect 19625 53941 19659 53975
rect 20361 53941 20395 53975
rect 21097 53941 21131 53975
rect 22201 53941 22235 53975
rect 22937 53941 22971 53975
rect 23949 53941 23983 53975
rect 25237 53941 25271 53975
rect 16405 53737 16439 53771
rect 18889 53737 18923 53771
rect 21281 53669 21315 53703
rect 23121 53669 23155 53703
rect 3249 53601 3283 53635
rect 6561 53601 6595 53635
rect 8401 53601 8435 53635
rect 11069 53601 11103 53635
rect 12725 53601 12759 53635
rect 24409 53601 24443 53635
rect 2237 53533 2271 53567
rect 3985 53533 4019 53567
rect 5549 53533 5583 53567
rect 7297 53533 7331 53567
rect 10609 53533 10643 53567
rect 12449 53533 12483 53567
rect 14289 53533 14323 53567
rect 14841 53533 14875 53567
rect 15669 53533 15703 53567
rect 16129 53533 16163 53567
rect 16681 53533 16715 53567
rect 17601 53533 17635 53567
rect 18245 53533 18279 53567
rect 18705 53533 18739 53567
rect 19441 53533 19475 53567
rect 20269 53533 20303 53567
rect 20729 53533 20763 53567
rect 21097 53533 21131 53567
rect 22017 53533 22051 53567
rect 22661 53533 22695 53567
rect 23305 53533 23339 53567
rect 23857 53533 23891 53567
rect 24593 53533 24627 53567
rect 25053 53533 25087 53567
rect 15853 53465 15887 53499
rect 18429 53465 18463 53499
rect 20453 53465 20487 53499
rect 24041 53465 24075 53499
rect 4629 53397 4663 53431
rect 14473 53397 14507 53431
rect 16865 53397 16899 53431
rect 17417 53397 17451 53431
rect 19625 53397 19659 53431
rect 21833 53397 21867 53431
rect 22477 53397 22511 53431
rect 25237 53397 25271 53431
rect 17325 53193 17359 53227
rect 19533 53193 19567 53227
rect 19717 53193 19751 53227
rect 21005 53193 21039 53227
rect 21833 53193 21867 53227
rect 22293 53193 22327 53227
rect 22569 53193 22603 53227
rect 23029 53193 23063 53227
rect 3985 53125 4019 53159
rect 5825 53125 5859 53159
rect 9137 53125 9171 53159
rect 13829 53125 13863 53159
rect 21189 53125 21223 53159
rect 1685 53057 1719 53091
rect 2973 53057 3007 53091
rect 4721 53057 4755 53091
rect 7941 53057 7975 53091
rect 9781 53057 9815 53091
rect 11897 53057 11931 53091
rect 14657 53057 14691 53091
rect 14933 53057 14967 53091
rect 16129 53057 16163 53091
rect 16405 53057 16439 53091
rect 19073 53057 19107 53091
rect 19349 53057 19383 53091
rect 20545 53057 20579 53091
rect 20821 53057 20855 53091
rect 23489 53057 23523 53091
rect 24133 53057 24167 53091
rect 24409 53057 24443 53091
rect 24777 53057 24811 53091
rect 25053 53057 25087 53091
rect 10333 52989 10367 53023
rect 12357 52989 12391 53023
rect 14013 52921 14047 52955
rect 2329 52853 2363 52887
rect 14473 52853 14507 52887
rect 15945 52853 15979 52887
rect 18889 52853 18923 52887
rect 20361 52853 20395 52887
rect 23305 52853 23339 52887
rect 23949 52853 23983 52887
rect 25237 52853 25271 52887
rect 12633 52649 12667 52683
rect 14105 52649 14139 52683
rect 24593 52649 24627 52683
rect 25237 52581 25271 52615
rect 3249 52513 3283 52547
rect 3985 52513 4019 52547
rect 4261 52513 4295 52547
rect 7757 52513 7791 52547
rect 11253 52513 11287 52547
rect 2237 52445 2271 52479
rect 5457 52445 5491 52479
rect 6561 52445 6595 52479
rect 7389 52445 7423 52479
rect 10793 52445 10827 52479
rect 12817 52445 12851 52479
rect 13645 52445 13679 52479
rect 24777 52445 24811 52479
rect 25053 52445 25087 52479
rect 13461 52377 13495 52411
rect 2237 52105 2271 52139
rect 7021 52105 7055 52139
rect 11713 52105 11747 52139
rect 12357 52105 12391 52139
rect 13277 52105 13311 52139
rect 25329 52105 25363 52139
rect 6929 52037 6963 52071
rect 1593 51969 1627 52003
rect 2973 51969 3007 52003
rect 4813 51969 4847 52003
rect 8033 51969 8067 52003
rect 9689 51969 9723 52003
rect 11897 51969 11931 52003
rect 12541 51969 12575 52003
rect 3341 51901 3375 51935
rect 5089 51901 5123 51935
rect 8493 51901 8527 51935
rect 10149 51901 10183 51935
rect 25513 51765 25547 51799
rect 10241 51561 10275 51595
rect 2881 51425 2915 51459
rect 7573 51425 7607 51459
rect 2237 51357 2271 51391
rect 3985 51357 4019 51391
rect 5457 51357 5491 51391
rect 7113 51357 7147 51391
rect 10425 51357 10459 51391
rect 25053 51357 25087 51391
rect 6193 51289 6227 51323
rect 4629 51221 4663 51255
rect 25237 51221 25271 51255
rect 1593 51017 1627 51051
rect 6929 51017 6963 51051
rect 9597 50949 9631 50983
rect 1777 50881 1811 50915
rect 2513 50881 2547 50915
rect 4261 50881 4295 50915
rect 6837 50881 6871 50915
rect 7757 50881 7791 50915
rect 9413 50881 9447 50915
rect 24777 50881 24811 50915
rect 25053 50881 25087 50915
rect 2789 50813 2823 50847
rect 4629 50813 4663 50847
rect 7481 50813 7515 50847
rect 25237 50677 25271 50711
rect 6837 50473 6871 50507
rect 9229 50473 9263 50507
rect 3249 50337 3283 50371
rect 3985 50337 4019 50371
rect 5089 50337 5123 50371
rect 2237 50269 2271 50303
rect 4261 50269 4295 50303
rect 7021 50269 7055 50303
rect 9413 50269 9447 50303
rect 25421 50133 25455 50167
rect 6561 49929 6595 49963
rect 25145 49929 25179 49963
rect 3157 49861 3191 49895
rect 4261 49861 4295 49895
rect 6377 49861 6411 49895
rect 9321 49861 9355 49895
rect 1961 49793 1995 49827
rect 3985 49793 4019 49827
rect 9137 49793 9171 49827
rect 25329 49793 25363 49827
rect 6009 49725 6043 49759
rect 11621 49385 11655 49419
rect 2053 49249 2087 49283
rect 1777 49181 1811 49215
rect 11805 49181 11839 49215
rect 24869 49181 24903 49215
rect 25329 49181 25363 49215
rect 3341 49045 3375 49079
rect 25145 49045 25179 49079
rect 12725 48841 12759 48875
rect 12909 48705 12943 48739
rect 25513 48501 25547 48535
rect 24869 48093 24903 48127
rect 25329 48093 25363 48127
rect 1685 48025 1719 48059
rect 2145 48025 2179 48059
rect 1777 47957 1811 47991
rect 17693 47957 17727 47991
rect 25145 47957 25179 47991
rect 9137 47753 9171 47787
rect 17233 47753 17267 47787
rect 18429 47753 18463 47787
rect 9321 47617 9355 47651
rect 17325 47617 17359 47651
rect 18521 47617 18555 47651
rect 19073 47617 19107 47651
rect 24501 47617 24535 47651
rect 17417 47549 17451 47583
rect 18613 47549 18647 47583
rect 24777 47549 24811 47583
rect 16865 47413 16899 47447
rect 18061 47413 18095 47447
rect 9873 47209 9907 47243
rect 15932 47209 15966 47243
rect 18153 47141 18187 47175
rect 25145 47141 25179 47175
rect 10241 47073 10275 47107
rect 15669 47073 15703 47107
rect 17417 47073 17451 47107
rect 18613 47073 18647 47107
rect 18797 47073 18831 47107
rect 22477 47073 22511 47107
rect 22661 47073 22695 47107
rect 22385 47005 22419 47039
rect 25329 47005 25363 47039
rect 10517 46937 10551 46971
rect 12265 46937 12299 46971
rect 14197 46937 14231 46971
rect 18521 46937 18555 46971
rect 19257 46937 19291 46971
rect 21649 46937 21683 46971
rect 24869 46937 24903 46971
rect 11989 46869 12023 46903
rect 17693 46869 17727 46903
rect 22017 46869 22051 46903
rect 7205 46665 7239 46699
rect 10885 46665 10919 46699
rect 18613 46665 18647 46699
rect 20821 46665 20855 46699
rect 22661 46665 22695 46699
rect 22753 46665 22787 46699
rect 12633 46597 12667 46631
rect 7389 46529 7423 46563
rect 11069 46529 11103 46563
rect 12357 46461 12391 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 16865 46461 16899 46495
rect 17141 46461 17175 46495
rect 19073 46461 19107 46495
rect 19349 46461 19383 46495
rect 22845 46461 22879 46495
rect 23305 46461 23339 46495
rect 24501 46461 24535 46495
rect 24777 46461 24811 46495
rect 14105 46325 14139 46359
rect 16313 46325 16347 46359
rect 21097 46325 21131 46359
rect 21925 46325 21959 46359
rect 22293 46325 22327 46359
rect 8125 46121 8159 46155
rect 9137 46121 9171 46155
rect 10701 46121 10735 46155
rect 18705 46121 18739 46155
rect 25421 46121 25455 46155
rect 10057 46053 10091 46087
rect 1869 45985 1903 46019
rect 11345 45985 11379 46019
rect 11897 45985 11931 46019
rect 12173 45985 12207 46019
rect 14105 45985 14139 46019
rect 20177 45985 20211 46019
rect 20361 45985 20395 46019
rect 21373 45985 21407 46019
rect 21465 45985 21499 46019
rect 1593 45917 1627 45951
rect 9321 45917 9355 45951
rect 10241 45917 10275 45951
rect 23213 45917 23247 45951
rect 23489 45917 23523 45951
rect 8033 45849 8067 45883
rect 8493 45849 8527 45883
rect 11069 45849 11103 45883
rect 19441 45849 19475 45883
rect 11161 45781 11195 45815
rect 13645 45781 13679 45815
rect 16405 45781 16439 45815
rect 19717 45781 19751 45815
rect 20085 45781 20119 45815
rect 20913 45781 20947 45815
rect 21281 45781 21315 45815
rect 24501 45781 24535 45815
rect 1409 45577 1443 45611
rect 16405 45577 16439 45611
rect 20177 45577 20211 45611
rect 23765 45577 23799 45611
rect 8861 45509 8895 45543
rect 9229 45441 9263 45475
rect 11253 45441 11287 45475
rect 24041 45441 24075 45475
rect 24777 45441 24811 45475
rect 9505 45373 9539 45407
rect 11529 45373 11563 45407
rect 14381 45373 14415 45407
rect 14657 45373 14691 45407
rect 18429 45373 18463 45407
rect 18705 45373 18739 45407
rect 20453 45373 20487 45407
rect 22017 45373 22051 45407
rect 22293 45373 22327 45407
rect 24501 45373 24535 45407
rect 10977 45305 11011 45339
rect 20729 45305 20763 45339
rect 12173 45237 12207 45271
rect 16129 45237 16163 45271
rect 9321 45033 9355 45067
rect 11621 45033 11655 45067
rect 12449 45033 12483 45067
rect 13001 45033 13035 45067
rect 15380 45033 15414 45067
rect 16865 45033 16899 45067
rect 7941 44965 7975 44999
rect 13553 44897 13587 44931
rect 15117 44897 15151 44931
rect 24409 44897 24443 44931
rect 12357 44829 12391 44863
rect 19533 44829 19567 44863
rect 21557 44829 21591 44863
rect 22293 44829 22327 44863
rect 7757 44761 7791 44795
rect 9229 44761 9263 44795
rect 11161 44761 11195 44795
rect 11529 44761 11563 44795
rect 19809 44761 19843 44795
rect 22569 44761 22603 44795
rect 6469 44693 6503 44727
rect 7113 44693 7147 44727
rect 8309 44693 8343 44727
rect 9781 44693 9815 44727
rect 13369 44693 13403 44727
rect 13461 44693 13495 44727
rect 17141 44693 17175 44727
rect 21281 44693 21315 44727
rect 24041 44693 24075 44727
rect 25513 44693 25547 44727
rect 5825 44489 5859 44523
rect 6745 44489 6779 44523
rect 8033 44489 8067 44523
rect 11069 44489 11103 44523
rect 11897 44489 11931 44523
rect 14933 44489 14967 44523
rect 15393 44489 15427 44523
rect 18613 44489 18647 44523
rect 21281 44489 21315 44523
rect 24041 44489 24075 44523
rect 7573 44421 7607 44455
rect 13461 44421 13495 44455
rect 18889 44421 18923 44455
rect 21557 44421 21591 44455
rect 6009 44353 6043 44387
rect 6653 44353 6687 44387
rect 7389 44353 7423 44387
rect 8217 44353 8251 44387
rect 8953 44353 8987 44387
rect 10977 44353 11011 44387
rect 12265 44353 12299 44387
rect 13185 44353 13219 44387
rect 24501 44353 24535 44387
rect 9137 44285 9171 44319
rect 12357 44285 12391 44319
rect 12449 44285 12483 44319
rect 15209 44285 15243 44319
rect 16865 44285 16899 44319
rect 17141 44285 17175 44319
rect 19533 44285 19567 44319
rect 19809 44285 19843 44319
rect 22293 44285 22327 44319
rect 22569 44285 22603 44319
rect 24777 44285 24811 44319
rect 9505 44217 9539 44251
rect 11621 44149 11655 44183
rect 8401 43945 8435 43979
rect 11621 43945 11655 43979
rect 21649 43945 21683 43979
rect 24133 43945 24167 43979
rect 25421 43945 25455 43979
rect 6929 43877 6963 43911
rect 9137 43809 9171 43843
rect 22477 43809 22511 43843
rect 22661 43809 22695 43843
rect 8585 43741 8619 43775
rect 6745 43673 6779 43707
rect 9413 43673 9447 43707
rect 11529 43673 11563 43707
rect 11989 43673 12023 43707
rect 22385 43673 22419 43707
rect 7205 43605 7239 43639
rect 10885 43605 10919 43639
rect 17969 43605 18003 43639
rect 22017 43605 22051 43639
rect 25329 43605 25363 43639
rect 7757 43401 7791 43435
rect 8585 43401 8619 43435
rect 9505 43401 9539 43435
rect 10609 43401 10643 43435
rect 15025 43401 15059 43435
rect 15117 43401 15151 43435
rect 15669 43401 15703 43435
rect 17417 43401 17451 43435
rect 17509 43401 17543 43435
rect 20085 43401 20119 43435
rect 20453 43401 20487 43435
rect 21373 43401 21407 43435
rect 21649 43401 21683 43435
rect 22477 43401 22511 43435
rect 9597 43333 9631 43367
rect 11069 43333 11103 43367
rect 12633 43333 12667 43367
rect 16681 43333 16715 43367
rect 23857 43333 23891 43367
rect 1685 43265 1719 43299
rect 2145 43265 2179 43299
rect 7941 43265 7975 43299
rect 8493 43265 8527 43299
rect 10517 43265 10551 43299
rect 22385 43265 22419 43299
rect 9689 43197 9723 43231
rect 12357 43197 12391 43231
rect 15209 43197 15243 43231
rect 17693 43197 17727 43231
rect 18337 43197 18371 43231
rect 18613 43197 18647 43231
rect 22661 43197 22695 43231
rect 23581 43197 23615 43231
rect 1869 43129 1903 43163
rect 9137 43129 9171 43163
rect 14657 43129 14691 43163
rect 14105 43061 14139 43095
rect 17049 43061 17083 43095
rect 22017 43061 22051 43095
rect 25329 43061 25363 43095
rect 8677 42857 8711 42891
rect 8953 42857 8987 42891
rect 9137 42857 9171 42891
rect 9597 42857 9631 42891
rect 12909 42857 12943 42891
rect 14289 42857 14323 42891
rect 19796 42857 19830 42891
rect 25329 42857 25363 42891
rect 23443 42789 23477 42823
rect 4997 42721 5031 42755
rect 9321 42721 9355 42755
rect 10793 42721 10827 42755
rect 14841 42721 14875 42755
rect 17785 42721 17819 42755
rect 18153 42721 18187 42755
rect 19533 42721 19567 42755
rect 22293 42721 22327 42755
rect 22477 42721 22511 42755
rect 17601 42653 17635 42687
rect 18337 42653 18371 42687
rect 23213 42653 23247 42687
rect 4813 42585 4847 42619
rect 5273 42585 5307 42619
rect 11069 42585 11103 42619
rect 15117 42585 15151 42619
rect 17509 42585 17543 42619
rect 22201 42585 22235 42619
rect 8309 42517 8343 42551
rect 10333 42517 10367 42551
rect 12541 42517 12575 42551
rect 16589 42517 16623 42551
rect 17141 42517 17175 42551
rect 21281 42517 21315 42551
rect 21833 42517 21867 42551
rect 24501 42517 24535 42551
rect 4353 42313 4387 42347
rect 5089 42313 5123 42347
rect 6745 42313 6779 42347
rect 9689 42313 9723 42347
rect 11805 42313 11839 42347
rect 13001 42313 13035 42347
rect 15393 42313 15427 42347
rect 15853 42313 15887 42347
rect 16865 42313 16899 42347
rect 17233 42313 17267 42347
rect 18153 42313 18187 42347
rect 21281 42313 21315 42347
rect 25237 42313 25271 42347
rect 10149 42245 10183 42279
rect 12265 42245 12299 42279
rect 15761 42245 15795 42279
rect 21557 42245 21591 42279
rect 22017 42245 22051 42279
rect 3893 42177 3927 42211
rect 4261 42177 4295 42211
rect 4997 42177 5031 42211
rect 6653 42177 6687 42211
rect 7481 42177 7515 42211
rect 10057 42177 10091 42211
rect 12173 42177 12207 42211
rect 13369 42177 13403 42211
rect 14197 42177 14231 42211
rect 17877 42177 17911 42211
rect 18613 42177 18647 42211
rect 18889 42177 18923 42211
rect 20637 42177 20671 42211
rect 7757 42109 7791 42143
rect 10241 42109 10275 42143
rect 12449 42109 12483 42143
rect 13461 42109 13495 42143
rect 13645 42109 13679 42143
rect 15945 42109 15979 42143
rect 17325 42109 17359 42143
rect 17417 42109 17451 42143
rect 19625 42109 19659 42143
rect 20729 42109 20763 42143
rect 20821 42109 20855 42143
rect 22845 42109 22879 42143
rect 23489 42109 23523 42143
rect 23765 42109 23799 42143
rect 5549 41973 5583 42007
rect 7205 41973 7239 42007
rect 9229 41973 9263 42007
rect 10701 41973 10735 42007
rect 16405 41973 16439 42007
rect 20269 41973 20303 42007
rect 5181 41769 5215 41803
rect 7665 41769 7699 41803
rect 8125 41769 8159 41803
rect 10701 41769 10735 41803
rect 17325 41769 17359 41803
rect 24593 41769 24627 41803
rect 8033 41701 8067 41735
rect 21189 41701 21223 41735
rect 21649 41701 21683 41735
rect 22845 41701 22879 41735
rect 25145 41701 25179 41735
rect 5917 41633 5951 41667
rect 10057 41633 10091 41667
rect 11253 41633 11287 41667
rect 12817 41633 12851 41667
rect 16681 41633 16715 41667
rect 16773 41633 16807 41667
rect 18613 41633 18647 41667
rect 18797 41633 18831 41667
rect 19717 41633 19751 41667
rect 22293 41633 22327 41667
rect 23305 41633 23339 41667
rect 23397 41633 23431 41667
rect 9321 41565 9355 41599
rect 11989 41565 12023 41599
rect 13185 41565 13219 41599
rect 19441 41565 19475 41599
rect 24501 41565 24535 41599
rect 25329 41565 25363 41599
rect 5089 41497 5123 41531
rect 6193 41497 6227 41531
rect 11161 41497 11195 41531
rect 16589 41497 16623 41531
rect 18521 41497 18555 41531
rect 22109 41497 22143 41531
rect 23213 41497 23247 41531
rect 24225 41497 24259 41531
rect 5641 41429 5675 41463
rect 11069 41429 11103 41463
rect 16221 41429 16255 41463
rect 18153 41429 18187 41463
rect 22017 41429 22051 41463
rect 24869 41429 24903 41463
rect 3341 41225 3375 41259
rect 8033 41225 8067 41259
rect 10977 41225 11011 41259
rect 11713 41225 11747 41259
rect 15761 41225 15795 41259
rect 18981 41225 19015 41259
rect 19901 41225 19935 41259
rect 21097 41225 21131 41259
rect 22017 41225 22051 41259
rect 24685 41225 24719 41259
rect 23213 41157 23247 41191
rect 1777 41089 1811 41123
rect 2053 41089 2087 41123
rect 3249 41089 3283 41123
rect 3709 41089 3743 41123
rect 8953 41089 8987 41123
rect 12081 41089 12115 41123
rect 12173 41089 12207 41123
rect 13645 41089 13679 41123
rect 16865 41089 16899 41123
rect 19809 41089 19843 41123
rect 25329 41089 25363 41123
rect 9229 41021 9263 41055
rect 12265 41021 12299 41055
rect 13921 41021 13955 41055
rect 17141 41021 17175 41055
rect 20085 41021 20119 41055
rect 21189 41021 21223 41055
rect 21281 41021 21315 41055
rect 22937 41021 22971 41055
rect 15393 40953 15427 40987
rect 1593 40885 1627 40919
rect 10701 40885 10735 40919
rect 18613 40885 18647 40919
rect 19165 40885 19199 40919
rect 19441 40885 19475 40919
rect 20729 40885 20763 40919
rect 25145 40885 25179 40919
rect 8585 40681 8619 40715
rect 10609 40681 10643 40715
rect 14749 40681 14783 40715
rect 16313 40681 16347 40715
rect 20913 40681 20947 40715
rect 24041 40681 24075 40715
rect 24409 40681 24443 40715
rect 9229 40613 9263 40647
rect 11069 40613 11103 40647
rect 14841 40613 14875 40647
rect 25145 40613 25179 40647
rect 6469 40545 6503 40579
rect 9873 40545 9907 40579
rect 11529 40545 11563 40579
rect 11713 40545 11747 40579
rect 13277 40545 13311 40579
rect 15669 40545 15703 40579
rect 15853 40545 15887 40579
rect 17141 40545 17175 40579
rect 17233 40545 17267 40579
rect 21465 40545 21499 40579
rect 22937 40545 22971 40579
rect 23121 40545 23155 40579
rect 6193 40477 6227 40511
rect 13001 40477 13035 40511
rect 15577 40477 15611 40511
rect 21373 40477 21407 40511
rect 22845 40477 22879 40511
rect 24685 40477 24719 40511
rect 25329 40477 25363 40511
rect 9597 40409 9631 40443
rect 11345 40409 11379 40443
rect 11805 40409 11839 40443
rect 13093 40409 13127 40443
rect 13737 40409 13771 40443
rect 21925 40409 21959 40443
rect 22201 40409 22235 40443
rect 24225 40409 24259 40443
rect 24869 40409 24903 40443
rect 7941 40341 7975 40375
rect 8309 40341 8343 40375
rect 8769 40341 8803 40375
rect 9689 40341 9723 40375
rect 10333 40341 10367 40375
rect 12173 40341 12207 40375
rect 12633 40341 12667 40375
rect 15209 40341 15243 40375
rect 16681 40341 16715 40375
rect 17049 40341 17083 40375
rect 20361 40341 20395 40375
rect 21281 40341 21315 40375
rect 22477 40341 22511 40375
rect 7297 40137 7331 40171
rect 11529 40137 11563 40171
rect 12265 40137 12299 40171
rect 15577 40137 15611 40171
rect 18245 40137 18279 40171
rect 18705 40137 18739 40171
rect 19809 40137 19843 40171
rect 25237 40137 25271 40171
rect 7665 40069 7699 40103
rect 10517 40069 10551 40103
rect 15025 40069 15059 40103
rect 15945 40069 15979 40103
rect 18613 40069 18647 40103
rect 20177 40069 20211 40103
rect 8493 40001 8527 40035
rect 12909 40001 12943 40035
rect 20821 40001 20855 40035
rect 22293 40001 22327 40035
rect 22569 40001 22603 40035
rect 23489 40001 23523 40035
rect 7757 39933 7791 39967
rect 7849 39933 7883 39967
rect 8769 39933 8803 39967
rect 10977 39933 11011 39967
rect 13185 39933 13219 39967
rect 16037 39933 16071 39967
rect 16129 39933 16163 39967
rect 18797 39933 18831 39967
rect 20269 39933 20303 39967
rect 20361 39933 20395 39967
rect 23765 39933 23799 39967
rect 14657 39797 14691 39831
rect 16681 39797 16715 39831
rect 21005 39797 21039 39831
rect 6653 39593 6687 39627
rect 9781 39593 9815 39627
rect 18797 39593 18831 39627
rect 19073 39593 19107 39627
rect 21281 39593 21315 39627
rect 15577 39525 15611 39559
rect 22661 39525 22695 39559
rect 4905 39457 4939 39491
rect 7113 39457 7147 39491
rect 10241 39457 10275 39491
rect 10333 39457 10367 39491
rect 10977 39457 11011 39491
rect 13921 39457 13955 39491
rect 14841 39457 14875 39491
rect 15025 39457 15059 39491
rect 16221 39457 16255 39491
rect 19901 39457 19935 39491
rect 20085 39457 20119 39491
rect 21741 39457 21775 39491
rect 21925 39457 21959 39491
rect 23305 39457 23339 39491
rect 25053 39457 25087 39491
rect 25145 39457 25179 39491
rect 13093 39389 13127 39423
rect 21649 39389 21683 39423
rect 23121 39389 23155 39423
rect 24961 39389 24995 39423
rect 5181 39321 5215 39355
rect 11253 39321 11287 39355
rect 14749 39321 14783 39355
rect 19809 39321 19843 39355
rect 23029 39321 23063 39355
rect 23857 39321 23891 39355
rect 7021 39253 7055 39287
rect 9137 39253 9171 39287
rect 10149 39253 10183 39287
rect 12725 39253 12759 39287
rect 13277 39253 13311 39287
rect 14381 39253 14415 39287
rect 15945 39253 15979 39287
rect 16037 39253 16071 39287
rect 18613 39253 18647 39287
rect 19441 39253 19475 39287
rect 20453 39253 20487 39287
rect 22293 39253 22327 39287
rect 24593 39253 24627 39287
rect 8217 39049 8251 39083
rect 9505 39049 9539 39083
rect 10793 39049 10827 39083
rect 14289 39049 14323 39083
rect 15301 39049 15335 39083
rect 19165 39049 19199 39083
rect 19533 39049 19567 39083
rect 20729 39049 20763 39083
rect 24501 39049 24535 39083
rect 8309 38981 8343 39015
rect 9597 38981 9631 39015
rect 18337 38981 18371 39015
rect 19625 38981 19659 39015
rect 22385 38981 22419 39015
rect 12081 38913 12115 38947
rect 15393 38913 15427 38947
rect 15945 38913 15979 38947
rect 24685 38913 24719 38947
rect 25329 38913 25363 38947
rect 9689 38845 9723 38879
rect 10885 38845 10919 38879
rect 10977 38845 11011 38879
rect 12357 38845 12391 38879
rect 15577 38845 15611 38879
rect 16865 38845 16899 38879
rect 18429 38845 18463 38879
rect 18613 38845 18647 38879
rect 19717 38845 19751 38879
rect 20821 38845 20855 38879
rect 20913 38845 20947 38879
rect 22109 38845 22143 38879
rect 24225 38845 24259 38879
rect 8677 38777 8711 38811
rect 10425 38777 10459 38811
rect 13829 38777 13863 38811
rect 7389 38709 7423 38743
rect 8493 38709 8527 38743
rect 9137 38709 9171 38743
rect 11529 38709 11563 38743
rect 14933 38709 14967 38743
rect 17969 38709 18003 38743
rect 20361 38709 20395 38743
rect 23857 38709 23891 38743
rect 25145 38709 25179 38743
rect 7849 38505 7883 38539
rect 10425 38505 10459 38539
rect 11897 38505 11931 38539
rect 14289 38505 14323 38539
rect 19441 38505 19475 38539
rect 20637 38505 20671 38539
rect 18153 38437 18187 38471
rect 22017 38437 22051 38471
rect 5733 38369 5767 38403
rect 7205 38369 7239 38403
rect 8493 38369 8527 38403
rect 9689 38369 9723 38403
rect 9781 38369 9815 38403
rect 10977 38369 11011 38403
rect 12357 38369 12391 38403
rect 12449 38369 12483 38403
rect 13921 38369 13955 38403
rect 14841 38369 14875 38403
rect 16221 38369 16255 38403
rect 18705 38369 18739 38403
rect 19993 38369 20027 38403
rect 21097 38369 21131 38403
rect 21189 38369 21223 38403
rect 22477 38369 22511 38403
rect 22569 38369 22603 38403
rect 23765 38369 23799 38403
rect 25145 38369 25179 38403
rect 1777 38301 1811 38335
rect 2053 38301 2087 38335
rect 5457 38301 5491 38335
rect 8217 38301 8251 38335
rect 14749 38301 14783 38335
rect 15945 38301 15979 38335
rect 18521 38301 18555 38335
rect 21005 38301 21039 38335
rect 25053 38301 25087 38335
rect 9597 38233 9631 38267
rect 19901 38233 19935 38267
rect 22385 38233 22419 38267
rect 23581 38233 23615 38267
rect 23673 38233 23707 38267
rect 1593 38165 1627 38199
rect 7573 38165 7607 38199
rect 8309 38165 8343 38199
rect 9229 38165 9263 38199
rect 10793 38165 10827 38199
rect 10885 38165 10919 38199
rect 12265 38165 12299 38199
rect 12909 38165 12943 38199
rect 13277 38165 13311 38199
rect 14657 38165 14691 38199
rect 17693 38165 17727 38199
rect 18613 38165 18647 38199
rect 19809 38165 19843 38199
rect 21649 38165 21683 38199
rect 23213 38165 23247 38199
rect 24593 38165 24627 38199
rect 24961 38165 24995 38199
rect 5273 37961 5307 37995
rect 5733 37961 5767 37995
rect 9137 37961 9171 37995
rect 10057 37961 10091 37995
rect 11713 37961 11747 37995
rect 12357 37961 12391 37995
rect 12725 37961 12759 37995
rect 15485 37961 15519 37995
rect 17233 37961 17267 37995
rect 18061 37961 18095 37995
rect 18337 37961 18371 37995
rect 18981 37961 19015 37995
rect 21557 37961 21591 37995
rect 22017 37961 22051 37995
rect 6837 37893 6871 37927
rect 11345 37893 11379 37927
rect 17877 37893 17911 37927
rect 18521 37893 18555 37927
rect 19441 37893 19475 37927
rect 20637 37893 20671 37927
rect 21281 37893 21315 37927
rect 22477 37893 22511 37927
rect 23121 37893 23155 37927
rect 23857 37893 23891 37927
rect 5641 37825 5675 37859
rect 9413 37825 9447 37859
rect 10425 37825 10459 37859
rect 14381 37825 14415 37859
rect 15393 37825 15427 37859
rect 17325 37825 17359 37859
rect 19349 37825 19383 37859
rect 20729 37825 20763 37859
rect 22385 37825 22419 37859
rect 23213 37825 23247 37859
rect 5825 37757 5859 37791
rect 6561 37757 6595 37791
rect 8585 37757 8619 37791
rect 8953 37757 8987 37791
rect 10517 37757 10551 37791
rect 10609 37757 10643 37791
rect 12817 37757 12851 37791
rect 13001 37757 13035 37791
rect 13553 37757 13587 37791
rect 15669 37757 15703 37791
rect 17509 37757 17543 37791
rect 19625 37757 19659 37791
rect 20913 37757 20947 37791
rect 22661 37757 22695 37791
rect 23581 37757 23615 37791
rect 25329 37757 25363 37791
rect 15025 37689 15059 37723
rect 16405 37689 16439 37723
rect 20269 37689 20303 37723
rect 14105 37621 14139 37655
rect 16129 37621 16163 37655
rect 16865 37621 16899 37655
rect 18613 37621 18647 37655
rect 8585 37417 8619 37451
rect 10425 37417 10459 37451
rect 10609 37417 10643 37451
rect 14933 37417 14967 37451
rect 12449 37349 12483 37383
rect 12909 37349 12943 37383
rect 14565 37349 14599 37383
rect 17325 37349 17359 37383
rect 7113 37281 7147 37315
rect 10977 37281 11011 37315
rect 11805 37281 11839 37315
rect 13369 37281 13403 37315
rect 13461 37281 13495 37315
rect 15485 37281 15519 37315
rect 16589 37281 16623 37315
rect 16681 37281 16715 37315
rect 17877 37281 17911 37315
rect 19073 37281 19107 37315
rect 24041 37281 24075 37315
rect 24225 37281 24259 37315
rect 24593 37281 24627 37315
rect 6837 37213 6871 37247
rect 9873 37213 9907 37247
rect 11621 37213 11655 37247
rect 13277 37213 13311 37247
rect 17785 37213 17819 37247
rect 21097 37213 21131 37247
rect 21465 37213 21499 37247
rect 22201 37213 22235 37247
rect 25329 37213 25363 37247
rect 9137 37145 9171 37179
rect 11713 37145 11747 37179
rect 16497 37145 16531 37179
rect 17693 37145 17727 37179
rect 19441 37145 19475 37179
rect 20177 37145 20211 37179
rect 11253 37077 11287 37111
rect 12633 37077 12667 37111
rect 14197 37077 14231 37111
rect 14473 37077 14507 37111
rect 15301 37077 15335 37111
rect 15393 37077 15427 37111
rect 16129 37077 16163 37111
rect 18521 37077 18555 37111
rect 20729 37077 20763 37111
rect 23765 37077 23799 37111
rect 24777 37077 24811 37111
rect 25145 37077 25179 37111
rect 7481 36873 7515 36907
rect 7941 36873 7975 36907
rect 9045 36873 9079 36907
rect 12173 36873 12207 36907
rect 12633 36873 12667 36907
rect 13829 36873 13863 36907
rect 15025 36873 15059 36907
rect 15577 36873 15611 36907
rect 17049 36873 17083 36907
rect 17417 36873 17451 36907
rect 20361 36873 20395 36907
rect 20453 36873 20487 36907
rect 21005 36873 21039 36907
rect 24593 36873 24627 36907
rect 10241 36805 10275 36839
rect 11529 36805 11563 36839
rect 12081 36805 12115 36839
rect 12541 36805 12575 36839
rect 23121 36805 23155 36839
rect 3985 36737 4019 36771
rect 7849 36737 7883 36771
rect 9413 36737 9447 36771
rect 9505 36737 9539 36771
rect 13737 36737 13771 36771
rect 14933 36737 14967 36771
rect 16681 36737 16715 36771
rect 17509 36737 17543 36771
rect 22845 36737 22879 36771
rect 25329 36737 25363 36771
rect 4261 36669 4295 36703
rect 5733 36669 5767 36703
rect 8033 36669 8067 36703
rect 9597 36669 9631 36703
rect 10977 36669 11011 36703
rect 12725 36669 12759 36703
rect 14013 36669 14047 36703
rect 15117 36669 15151 36703
rect 15853 36669 15887 36703
rect 17601 36669 17635 36703
rect 20545 36669 20579 36703
rect 11805 36601 11839 36635
rect 19349 36601 19383 36635
rect 6101 36533 6135 36567
rect 8769 36533 8803 36567
rect 13369 36533 13403 36567
rect 14565 36533 14599 36567
rect 19993 36533 20027 36567
rect 25145 36533 25179 36567
rect 7665 36329 7699 36363
rect 9137 36329 9171 36363
rect 12173 36329 12207 36363
rect 12725 36329 12759 36363
rect 14289 36329 14323 36363
rect 19441 36329 19475 36363
rect 25145 36329 25179 36363
rect 16129 36261 16163 36295
rect 23305 36261 23339 36295
rect 8217 36193 8251 36227
rect 9689 36193 9723 36227
rect 12449 36193 12483 36227
rect 13185 36193 13219 36227
rect 13369 36193 13403 36227
rect 14933 36193 14967 36227
rect 15761 36193 15795 36227
rect 16681 36193 16715 36227
rect 19073 36193 19107 36227
rect 19993 36193 20027 36227
rect 21281 36193 21315 36227
rect 21465 36193 21499 36227
rect 23765 36193 23799 36227
rect 23949 36193 23983 36227
rect 1777 36125 1811 36159
rect 2053 36125 2087 36159
rect 9597 36125 9631 36159
rect 16589 36125 16623 36159
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 8125 36057 8159 36091
rect 13829 36057 13863 36091
rect 14749 36057 14783 36091
rect 16497 36057 16531 36091
rect 17325 36057 17359 36091
rect 19901 36057 19935 36091
rect 1593 35989 1627 36023
rect 8033 35989 8067 36023
rect 9505 35989 9539 36023
rect 13093 35989 13127 36023
rect 14657 35989 14691 36023
rect 19809 35989 19843 36023
rect 20821 35989 20855 36023
rect 21189 35989 21223 36023
rect 23673 35989 23707 36023
rect 6009 35785 6043 35819
rect 14473 35785 14507 35819
rect 19349 35785 19383 35819
rect 24869 35785 24903 35819
rect 10149 35717 10183 35751
rect 14013 35717 14047 35751
rect 17877 35717 17911 35751
rect 4261 35649 4295 35683
rect 20177 35649 20211 35683
rect 23121 35649 23155 35683
rect 4537 35581 4571 35615
rect 8125 35581 8159 35615
rect 8401 35581 8435 35615
rect 11713 35581 11747 35615
rect 11989 35581 12023 35615
rect 17601 35581 17635 35615
rect 20269 35581 20303 35615
rect 20361 35581 20395 35615
rect 22477 35581 22511 35615
rect 23397 35581 23431 35615
rect 13461 35513 13495 35547
rect 6469 35445 6503 35479
rect 9873 35445 9907 35479
rect 13737 35445 13771 35479
rect 19809 35445 19843 35479
rect 20913 35445 20947 35479
rect 25237 35445 25271 35479
rect 25421 35445 25455 35479
rect 9321 35241 9355 35275
rect 13001 35241 13035 35275
rect 17141 35241 17175 35275
rect 21557 35241 21591 35275
rect 7849 35173 7883 35207
rect 6101 35105 6135 35139
rect 6377 35105 6411 35139
rect 9873 35105 9907 35139
rect 13553 35105 13587 35139
rect 15393 35105 15427 35139
rect 17417 35105 17451 35139
rect 19441 35105 19475 35139
rect 21189 35105 21223 35139
rect 21833 35105 21867 35139
rect 13461 35037 13495 35071
rect 22293 35037 22327 35071
rect 25329 35037 25363 35071
rect 9689 34969 9723 35003
rect 9781 34969 9815 35003
rect 15669 34969 15703 35003
rect 19717 34969 19751 35003
rect 22569 34969 22603 35003
rect 8125 34901 8159 34935
rect 13369 34901 13403 34935
rect 24041 34901 24075 34935
rect 24501 34901 24535 34935
rect 25145 34901 25179 34935
rect 8309 34697 8343 34731
rect 10609 34697 10643 34731
rect 13737 34697 13771 34731
rect 15577 34697 15611 34731
rect 15945 34697 15979 34731
rect 21097 34697 21131 34731
rect 21189 34697 21223 34731
rect 22385 34697 22419 34731
rect 23581 34697 23615 34731
rect 24409 34697 24443 34731
rect 25145 34697 25179 34731
rect 6837 34629 6871 34663
rect 16037 34629 16071 34663
rect 20269 34629 20303 34663
rect 6561 34561 6595 34595
rect 8861 34561 8895 34595
rect 22477 34561 22511 34595
rect 24593 34561 24627 34595
rect 25329 34561 25363 34595
rect 11713 34493 11747 34527
rect 13461 34493 13495 34527
rect 16129 34493 16163 34527
rect 21281 34493 21315 34527
rect 22569 34493 22603 34527
rect 23673 34493 23707 34527
rect 23765 34493 23799 34527
rect 23213 34425 23247 34459
rect 9124 34357 9158 34391
rect 10977 34357 11011 34391
rect 11976 34357 12010 34391
rect 20729 34357 20763 34391
rect 22017 34357 22051 34391
rect 5812 34153 5846 34187
rect 9137 34153 9171 34187
rect 12173 34153 12207 34187
rect 17693 34153 17727 34187
rect 20545 34153 20579 34187
rect 23305 34153 23339 34187
rect 25329 34153 25363 34187
rect 21097 34085 21131 34119
rect 5549 34017 5583 34051
rect 7297 34017 7331 34051
rect 9689 34017 9723 34051
rect 10701 34017 10735 34051
rect 13461 34017 13495 34051
rect 13553 34017 13587 34051
rect 15945 34017 15979 34051
rect 19073 34017 19107 34051
rect 19993 34017 20027 34051
rect 21649 34017 21683 34051
rect 22753 34017 22787 34051
rect 22937 34017 22971 34051
rect 7757 33949 7791 33983
rect 10425 33949 10459 33983
rect 12449 33949 12483 33983
rect 19809 33949 19843 33983
rect 21557 33949 21591 33983
rect 24777 33949 24811 33983
rect 9505 33881 9539 33915
rect 16221 33881 16255 33915
rect 19901 33881 19935 33915
rect 25421 33881 25455 33915
rect 7573 33813 7607 33847
rect 8493 33813 8527 33847
rect 9597 33813 9631 33847
rect 13001 33813 13035 33847
rect 13369 33813 13403 33847
rect 14105 33813 14139 33847
rect 17969 33813 18003 33847
rect 19441 33813 19475 33847
rect 20637 33813 20671 33847
rect 21465 33813 21499 33847
rect 22293 33813 22327 33847
rect 22661 33813 22695 33847
rect 24593 33813 24627 33847
rect 10425 33609 10459 33643
rect 10885 33609 10919 33643
rect 12909 33609 12943 33643
rect 13369 33609 13403 33643
rect 19809 33609 19843 33643
rect 20269 33609 20303 33643
rect 20729 33609 20763 33643
rect 21281 33609 21315 33643
rect 22661 33609 22695 33643
rect 25237 33609 25271 33643
rect 1777 33473 1811 33507
rect 2053 33473 2087 33507
rect 10793 33473 10827 33507
rect 13277 33473 13311 33507
rect 14105 33473 14139 33507
rect 18061 33473 18095 33507
rect 20637 33473 20671 33507
rect 23489 33473 23523 33507
rect 5365 33405 5399 33439
rect 9781 33405 9815 33439
rect 10977 33405 11011 33439
rect 12817 33405 12851 33439
rect 13461 33405 13495 33439
rect 14381 33405 14415 33439
rect 18337 33405 18371 33439
rect 20913 33405 20947 33439
rect 22017 33405 22051 33439
rect 23765 33405 23799 33439
rect 1593 33269 1627 33303
rect 7205 33269 7239 33303
rect 12541 33269 12575 33303
rect 15853 33269 15887 33303
rect 16129 33269 16163 33303
rect 7481 33065 7515 33099
rect 9413 33065 9447 33099
rect 10609 33065 10643 33099
rect 11161 33065 11195 33099
rect 12173 33065 12207 33099
rect 25145 33065 25179 33099
rect 7021 32997 7055 33031
rect 14289 32997 14323 33031
rect 17141 32997 17175 33031
rect 22937 32997 22971 33031
rect 5273 32929 5307 32963
rect 8125 32929 8159 32963
rect 10057 32929 10091 32963
rect 10885 32929 10919 32963
rect 11621 32929 11655 32963
rect 11805 32929 11839 32963
rect 14749 32929 14783 32963
rect 14841 32929 14875 32963
rect 16681 32929 16715 32963
rect 20269 32929 20303 32963
rect 20361 32929 20395 32963
rect 21649 32929 21683 32963
rect 9781 32861 9815 32895
rect 15761 32861 15795 32895
rect 16589 32861 16623 32895
rect 17325 32861 17359 32895
rect 20177 32861 20211 32895
rect 21373 32861 21407 32895
rect 22385 32861 22419 32895
rect 24869 32861 24903 32895
rect 25329 32861 25363 32895
rect 5549 32793 5583 32827
rect 7941 32793 7975 32827
rect 11529 32793 11563 32827
rect 19441 32793 19475 32827
rect 7849 32725 7883 32759
rect 9873 32725 9907 32759
rect 14657 32725 14691 32759
rect 16129 32725 16163 32759
rect 16497 32725 16531 32759
rect 17969 32725 18003 32759
rect 19809 32725 19843 32759
rect 21005 32725 21039 32759
rect 21465 32725 21499 32759
rect 22201 32725 22235 32759
rect 22661 32725 22695 32759
rect 4629 32521 4663 32555
rect 4997 32521 5031 32555
rect 5365 32521 5399 32555
rect 6929 32521 6963 32555
rect 11989 32521 12023 32555
rect 17325 32521 17359 32555
rect 19257 32521 19291 32555
rect 21189 32521 21223 32555
rect 21833 32521 21867 32555
rect 25145 32521 25179 32555
rect 5457 32453 5491 32487
rect 14841 32453 14875 32487
rect 17233 32453 17267 32487
rect 7573 32385 7607 32419
rect 12357 32385 12391 32419
rect 13185 32385 13219 32419
rect 14565 32385 14599 32419
rect 18429 32385 18463 32419
rect 18521 32385 18555 32419
rect 19073 32385 19107 32419
rect 20269 32385 20303 32419
rect 21097 32385 21131 32419
rect 22385 32385 22419 32419
rect 23029 32385 23063 32419
rect 24869 32385 24903 32419
rect 25329 32385 25363 32419
rect 5549 32317 5583 32351
rect 7849 32317 7883 32351
rect 9873 32317 9907 32351
rect 11713 32317 11747 32351
rect 12449 32317 12483 32351
rect 12541 32317 12575 32351
rect 16313 32317 16347 32351
rect 17509 32317 17543 32351
rect 18613 32317 18647 32351
rect 21373 32317 21407 32351
rect 9321 32181 9355 32215
rect 10333 32181 10367 32215
rect 16865 32181 16899 32215
rect 18061 32181 18095 32215
rect 20085 32181 20119 32215
rect 20729 32181 20763 32215
rect 22201 32181 22235 32215
rect 22845 32181 22879 32215
rect 23305 32181 23339 32215
rect 7941 31977 7975 32011
rect 8585 31977 8619 32011
rect 11161 31977 11195 32011
rect 16405 31977 16439 32011
rect 18061 31977 18095 32011
rect 25145 31977 25179 32011
rect 13921 31909 13955 31943
rect 14289 31909 14323 31943
rect 19441 31909 19475 31943
rect 20637 31909 20671 31943
rect 21925 31909 21959 31943
rect 6193 31841 6227 31875
rect 6469 31841 6503 31875
rect 9689 31841 9723 31875
rect 13645 31841 13679 31875
rect 14841 31841 14875 31875
rect 16957 31841 16991 31875
rect 18245 31841 18279 31875
rect 19993 31841 20027 31875
rect 21189 31841 21223 31875
rect 22385 31841 22419 31875
rect 22569 31841 22603 31875
rect 8309 31773 8343 31807
rect 9402 31773 9436 31807
rect 14749 31773 14783 31807
rect 16865 31773 16899 31807
rect 18429 31773 18463 31807
rect 19901 31773 19935 31807
rect 21097 31773 21131 31807
rect 24133 31773 24167 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 19809 31705 19843 31739
rect 21005 31705 21039 31739
rect 22293 31705 22327 31739
rect 9137 31637 9171 31671
rect 11437 31637 11471 31671
rect 14657 31637 14691 31671
rect 16773 31637 16807 31671
rect 7481 31433 7515 31467
rect 8677 31433 8711 31467
rect 9045 31433 9079 31467
rect 18337 31433 18371 31467
rect 20729 31433 20763 31467
rect 21557 31433 21591 31467
rect 25145 31433 25179 31467
rect 9781 31365 9815 31399
rect 14933 31365 14967 31399
rect 22477 31365 22511 31399
rect 1777 31297 1811 31331
rect 7849 31297 7883 31331
rect 7941 31297 7975 31331
rect 17509 31297 17543 31331
rect 17601 31297 17635 31331
rect 18705 31297 18739 31331
rect 19901 31297 19935 31331
rect 24593 31297 24627 31331
rect 25329 31297 25363 31331
rect 2053 31229 2087 31263
rect 7205 31229 7239 31263
rect 8125 31229 8159 31263
rect 9137 31229 9171 31263
rect 9321 31229 9355 31263
rect 12909 31229 12943 31263
rect 13185 31229 13219 31263
rect 16773 31229 16807 31263
rect 17785 31229 17819 31263
rect 18797 31229 18831 31263
rect 18889 31229 18923 31263
rect 19993 31229 20027 31263
rect 20177 31229 20211 31263
rect 22201 31229 22235 31263
rect 19533 31161 19567 31195
rect 14657 31093 14691 31127
rect 17141 31093 17175 31127
rect 20545 31093 20579 31127
rect 23949 31093 23983 31127
rect 24409 31093 24443 31127
rect 12817 30889 12851 30923
rect 20453 30889 20487 30923
rect 23029 30889 23063 30923
rect 24869 30889 24903 30923
rect 12449 30821 12483 30855
rect 25145 30821 25179 30855
rect 3985 30753 4019 30787
rect 7941 30753 7975 30787
rect 9597 30753 9631 30787
rect 9873 30753 9907 30787
rect 13369 30753 13403 30787
rect 16221 30753 16255 30787
rect 16497 30753 16531 30787
rect 19901 30753 19935 30787
rect 19993 30753 20027 30787
rect 22569 30753 22603 30787
rect 12265 30685 12299 30719
rect 13185 30685 13219 30719
rect 18245 30685 18279 30719
rect 19809 30685 19843 30719
rect 23857 30685 23891 30719
rect 25329 30685 25363 30719
rect 4169 30617 4203 30651
rect 5825 30617 5859 30651
rect 11621 30617 11655 30651
rect 13277 30617 13311 30651
rect 13921 30617 13955 30651
rect 22385 30617 22419 30651
rect 8493 30549 8527 30583
rect 11345 30549 11379 30583
rect 15853 30549 15887 30583
rect 17969 30549 18003 30583
rect 19441 30549 19475 30583
rect 22017 30549 22051 30583
rect 22477 30549 22511 30583
rect 23673 30549 23707 30583
rect 8953 30277 8987 30311
rect 12541 30277 12575 30311
rect 23673 30277 23707 30311
rect 25421 30277 25455 30311
rect 10793 30209 10827 30243
rect 11713 30209 11747 30243
rect 14473 30209 14507 30243
rect 17969 30209 18003 30243
rect 18613 30209 18647 30243
rect 19625 30209 19659 30243
rect 23397 30209 23431 30243
rect 10149 30141 10183 30175
rect 10885 30141 10919 30175
rect 10977 30141 11011 30175
rect 16221 30141 16255 30175
rect 16957 30141 16991 30175
rect 18061 30141 18095 30175
rect 18245 30141 18279 30175
rect 25145 30141 25179 30175
rect 10425 30005 10459 30039
rect 12265 30005 12299 30039
rect 14736 30005 14770 30039
rect 17601 30005 17635 30039
rect 18797 30005 18831 30039
rect 19441 30005 19475 30039
rect 7297 29801 7331 29835
rect 7849 29801 7883 29835
rect 9505 29801 9539 29835
rect 13737 29801 13771 29835
rect 16037 29801 16071 29835
rect 12633 29733 12667 29767
rect 21557 29733 21591 29767
rect 4261 29665 4295 29699
rect 8401 29665 8435 29699
rect 9229 29665 9263 29699
rect 10057 29665 10091 29699
rect 11989 29665 12023 29699
rect 13185 29665 13219 29699
rect 17509 29665 17543 29699
rect 18797 29665 18831 29699
rect 20085 29665 20119 29699
rect 20269 29665 20303 29699
rect 22201 29665 22235 29699
rect 23397 29665 23431 29699
rect 23581 29665 23615 29699
rect 13001 29597 13035 29631
rect 17417 29597 17451 29631
rect 19993 29597 20027 29631
rect 21925 29597 21959 29631
rect 25329 29597 25363 29631
rect 4445 29529 4479 29563
rect 6101 29529 6135 29563
rect 7481 29529 7515 29563
rect 8309 29529 8343 29563
rect 9873 29529 9907 29563
rect 11805 29529 11839 29563
rect 13093 29529 13127 29563
rect 14749 29529 14783 29563
rect 17325 29529 17359 29563
rect 18613 29529 18647 29563
rect 8217 29461 8251 29495
rect 9045 29461 9079 29495
rect 9965 29461 9999 29495
rect 11437 29461 11471 29495
rect 11897 29461 11931 29495
rect 16957 29461 16991 29495
rect 18153 29461 18187 29495
rect 18521 29461 18555 29495
rect 19625 29461 19659 29495
rect 20913 29461 20947 29495
rect 22017 29461 22051 29495
rect 22937 29461 22971 29495
rect 23305 29461 23339 29495
rect 25145 29461 25179 29495
rect 12909 29257 12943 29291
rect 14197 29257 14231 29291
rect 15301 29257 15335 29291
rect 16037 29257 16071 29291
rect 17233 29257 17267 29291
rect 17325 29257 17359 29291
rect 17969 29257 18003 29291
rect 22385 29257 22419 29291
rect 23949 29257 23983 29291
rect 25329 29257 25363 29291
rect 25513 29257 25547 29291
rect 9781 29189 9815 29223
rect 16221 29189 16255 29223
rect 21557 29189 21591 29223
rect 24685 29189 24719 29223
rect 13001 29121 13035 29155
rect 14105 29121 14139 29155
rect 19717 29121 19751 29155
rect 20453 29121 20487 29155
rect 20545 29121 20579 29155
rect 22477 29121 22511 29155
rect 23673 29121 23707 29155
rect 24133 29121 24167 29155
rect 7757 29053 7791 29087
rect 9505 29053 9539 29087
rect 13093 29053 13127 29087
rect 14381 29053 14415 29087
rect 15393 29053 15427 29087
rect 15485 29053 15519 29087
rect 16405 29053 16439 29087
rect 17417 29053 17451 29087
rect 20637 29053 20671 29087
rect 21097 29053 21131 29087
rect 22661 29053 22695 29087
rect 12541 28985 12575 29019
rect 13737 28985 13771 29019
rect 14933 28985 14967 29019
rect 16865 28985 16899 29019
rect 18061 28985 18095 29019
rect 20085 28985 20119 29019
rect 22017 28985 22051 29019
rect 24869 28985 24903 29019
rect 8020 28917 8054 28951
rect 12817 28713 12851 28747
rect 16773 28713 16807 28747
rect 21189 28645 21223 28679
rect 2053 28577 2087 28611
rect 4261 28577 4295 28611
rect 5641 28577 5675 28611
rect 6561 28577 6595 28611
rect 6837 28577 6871 28611
rect 8309 28577 8343 28611
rect 10885 28577 10919 28611
rect 13369 28577 13403 28611
rect 14841 28577 14875 28611
rect 16221 28577 16255 28611
rect 17693 28577 17727 28611
rect 17785 28577 17819 28611
rect 19441 28577 19475 28611
rect 1777 28509 1811 28543
rect 10609 28509 10643 28543
rect 14657 28509 14691 28543
rect 16037 28509 16071 28543
rect 16129 28509 16163 28543
rect 17601 28509 17635 28543
rect 24041 28509 24075 28543
rect 24777 28509 24811 28543
rect 4445 28441 4479 28475
rect 19717 28441 19751 28475
rect 21465 28441 21499 28475
rect 8677 28373 8711 28407
rect 12357 28373 12391 28407
rect 13185 28373 13219 28407
rect 13277 28373 13311 28407
rect 13921 28373 13955 28407
rect 14289 28373 14323 28407
rect 14749 28373 14783 28407
rect 15301 28373 15335 28407
rect 15669 28373 15703 28407
rect 17233 28373 17267 28407
rect 23857 28373 23891 28407
rect 24593 28373 24627 28407
rect 2053 28169 2087 28203
rect 3755 28169 3789 28203
rect 10333 28169 10367 28203
rect 12633 28169 12667 28203
rect 15945 28169 15979 28203
rect 16865 28169 16899 28203
rect 18337 28169 18371 28203
rect 19533 28169 19567 28203
rect 20177 28169 20211 28203
rect 24133 28169 24167 28203
rect 16773 28101 16807 28135
rect 24685 28101 24719 28135
rect 2237 28033 2271 28067
rect 3652 28033 3686 28067
rect 13185 28033 13219 28067
rect 18245 28033 18279 28067
rect 19441 28033 19475 28067
rect 22017 28033 22051 28067
rect 8309 27965 8343 27999
rect 8585 27965 8619 27999
rect 16037 27965 16071 27999
rect 16221 27965 16255 27999
rect 18521 27965 18555 27999
rect 19717 27965 19751 27999
rect 22293 27965 22327 27999
rect 10057 27897 10091 27931
rect 17049 27897 17083 27931
rect 24869 27897 24903 27931
rect 13277 27829 13311 27863
rect 15117 27829 15151 27863
rect 15577 27829 15611 27863
rect 17509 27829 17543 27863
rect 17877 27829 17911 27863
rect 19073 27829 19107 27863
rect 23765 27829 23799 27863
rect 6456 27625 6490 27659
rect 18705 27625 18739 27659
rect 24225 27625 24259 27659
rect 7941 27557 7975 27591
rect 8309 27557 8343 27591
rect 8401 27557 8435 27591
rect 20085 27557 20119 27591
rect 6193 27489 6227 27523
rect 15669 27489 15703 27523
rect 20545 27489 20579 27523
rect 20637 27489 20671 27523
rect 21925 27489 21959 27523
rect 11161 27421 11195 27455
rect 15577 27421 15611 27455
rect 16129 27421 16163 27455
rect 18337 27421 18371 27455
rect 24685 27421 24719 27455
rect 11437 27353 11471 27387
rect 22201 27353 22235 27387
rect 24869 27353 24903 27387
rect 12909 27285 12943 27319
rect 13277 27285 13311 27319
rect 15117 27285 15151 27319
rect 15485 27285 15519 27319
rect 16405 27285 16439 27319
rect 18153 27285 18187 27319
rect 18981 27285 19015 27319
rect 19809 27285 19843 27319
rect 20453 27285 20487 27319
rect 23673 27285 23707 27319
rect 25237 27285 25271 27319
rect 3203 27081 3237 27115
rect 15117 27081 15151 27115
rect 15209 27081 15243 27115
rect 17601 27081 17635 27115
rect 19993 27081 20027 27115
rect 10517 27013 10551 27047
rect 25145 27013 25179 27047
rect 3132 26945 3166 26979
rect 3709 26945 3743 26979
rect 6561 26945 6595 26979
rect 9137 26945 9171 26979
rect 12541 26945 12575 26979
rect 17969 26945 18003 26979
rect 19901 26945 19935 26979
rect 20729 26945 20763 26979
rect 22385 26945 22419 26979
rect 3893 26877 3927 26911
rect 4445 26877 4479 26911
rect 6837 26877 6871 26911
rect 9229 26877 9263 26911
rect 9413 26877 9447 26911
rect 12817 26877 12851 26911
rect 15301 26877 15335 26911
rect 18061 26877 18095 26911
rect 18245 26877 18279 26911
rect 20177 26877 20211 26911
rect 22845 26877 22879 26911
rect 23121 26877 23155 26911
rect 25329 26877 25363 26911
rect 8309 26809 8343 26843
rect 10701 26809 10735 26843
rect 8769 26741 8803 26775
rect 11897 26741 11931 26775
rect 14289 26741 14323 26775
rect 14749 26741 14783 26775
rect 17325 26741 17359 26775
rect 19533 26741 19567 26775
rect 22201 26741 22235 26775
rect 24593 26741 24627 26775
rect 4077 26537 4111 26571
rect 11713 26537 11747 26571
rect 17141 26537 17175 26571
rect 22385 26537 22419 26571
rect 17509 26469 17543 26503
rect 19441 26469 19475 26503
rect 22845 26469 22879 26503
rect 23857 26469 23891 26503
rect 25145 26469 25179 26503
rect 6469 26401 6503 26435
rect 6745 26401 6779 26435
rect 9137 26401 9171 26435
rect 10241 26401 10275 26435
rect 12725 26401 12759 26435
rect 15669 26401 15703 26435
rect 19901 26401 19935 26435
rect 20085 26401 20119 26435
rect 20637 26401 20671 26435
rect 23305 26401 23339 26435
rect 23397 26401 23431 26435
rect 1777 26333 1811 26367
rect 9965 26333 9999 26367
rect 12633 26333 12667 26367
rect 15393 26333 15427 26367
rect 19809 26333 19843 26367
rect 24869 26333 24903 26367
rect 2789 26265 2823 26299
rect 8677 26265 8711 26299
rect 17693 26265 17727 26299
rect 20913 26265 20947 26299
rect 23213 26265 23247 26299
rect 24685 26265 24719 26299
rect 8217 26197 8251 26231
rect 12173 26197 12207 26231
rect 12541 26197 12575 26231
rect 14473 26197 14507 26231
rect 2145 25993 2179 26027
rect 8585 25993 8619 26027
rect 9229 25993 9263 26027
rect 10793 25993 10827 26027
rect 10885 25993 10919 26027
rect 15853 25993 15887 26027
rect 19349 25993 19383 26027
rect 20269 25993 20303 26027
rect 20361 25993 20395 26027
rect 21005 25993 21039 26027
rect 22477 25993 22511 26027
rect 14841 25925 14875 25959
rect 23305 25925 23339 25959
rect 2329 25857 2363 25891
rect 3065 25857 3099 25891
rect 4169 25857 4203 25891
rect 8861 25857 8895 25891
rect 9597 25857 9631 25891
rect 12725 25857 12759 25891
rect 15761 25857 15795 25891
rect 17601 25857 17635 25891
rect 22385 25857 22419 25891
rect 23949 25857 23983 25891
rect 3249 25789 3283 25823
rect 8033 25789 8067 25823
rect 9689 25789 9723 25823
rect 9781 25789 9815 25823
rect 10977 25789 11011 25823
rect 11989 25789 12023 25823
rect 13001 25789 13035 25823
rect 14473 25789 14507 25823
rect 16037 25789 16071 25823
rect 17877 25789 17911 25823
rect 20545 25789 20579 25823
rect 21281 25789 21315 25823
rect 22569 25789 22603 25823
rect 25145 25789 25179 25823
rect 3433 25721 3467 25755
rect 4629 25721 4663 25755
rect 19901 25721 19935 25755
rect 23489 25721 23523 25755
rect 4261 25653 4295 25687
rect 10425 25653 10459 25687
rect 15393 25653 15427 25687
rect 22017 25653 22051 25687
rect 7100 25449 7134 25483
rect 8953 25449 8987 25483
rect 11437 25449 11471 25483
rect 14749 25449 14783 25483
rect 18061 25449 18095 25483
rect 23121 25449 23155 25483
rect 23397 25449 23431 25483
rect 25237 25449 25271 25483
rect 25513 25449 25547 25483
rect 10057 25381 10091 25415
rect 22109 25381 22143 25415
rect 6837 25313 6871 25347
rect 9413 25313 9447 25347
rect 10609 25313 10643 25347
rect 11989 25313 12023 25347
rect 13185 25313 13219 25347
rect 15301 25313 15335 25347
rect 15945 25313 15979 25347
rect 16221 25313 16255 25347
rect 19901 25313 19935 25347
rect 20085 25313 20119 25347
rect 22569 25313 22603 25347
rect 22753 25313 22787 25347
rect 4052 25245 4086 25279
rect 10425 25245 10459 25279
rect 10517 25245 10551 25279
rect 11805 25245 11839 25279
rect 13093 25245 13127 25279
rect 19809 25245 19843 25279
rect 22477 25245 22511 25279
rect 24685 25245 24719 25279
rect 23857 25177 23891 25211
rect 4123 25109 4157 25143
rect 8585 25109 8619 25143
rect 11069 25109 11103 25143
rect 11897 25109 11931 25143
rect 12633 25109 12667 25143
rect 13001 25109 13035 25143
rect 15117 25109 15151 25143
rect 15209 25109 15243 25143
rect 17693 25109 17727 25143
rect 18245 25109 18279 25143
rect 19441 25109 19475 25143
rect 23949 25109 23983 25143
rect 24777 25109 24811 25143
rect 5457 24905 5491 24939
rect 8033 24905 8067 24939
rect 15209 24905 15243 24939
rect 16865 24905 16899 24939
rect 18521 24905 18555 24939
rect 19901 24905 19935 24939
rect 20637 24905 20671 24939
rect 9229 24837 9263 24871
rect 12081 24837 12115 24871
rect 12817 24837 12851 24871
rect 17233 24837 17267 24871
rect 23213 24837 23247 24871
rect 7389 24769 7423 24803
rect 10057 24769 10091 24803
rect 12173 24769 12207 24803
rect 13185 24769 13219 24803
rect 13829 24769 13863 24803
rect 14565 24769 14599 24803
rect 15301 24769 15335 24803
rect 17325 24769 17359 24803
rect 18429 24769 18463 24803
rect 22937 24769 22971 24803
rect 25329 24769 25363 24803
rect 3709 24701 3743 24735
rect 3985 24701 4019 24735
rect 8125 24701 8159 24735
rect 8217 24701 8251 24735
rect 9321 24701 9355 24735
rect 9413 24701 9447 24735
rect 12265 24701 12299 24735
rect 13001 24701 13035 24735
rect 13921 24701 13955 24735
rect 14105 24701 14139 24735
rect 15393 24701 15427 24735
rect 17509 24701 17543 24735
rect 18613 24701 18647 24735
rect 20729 24701 20763 24735
rect 20821 24701 20855 24735
rect 24685 24701 24719 24735
rect 7665 24633 7699 24667
rect 11713 24633 11747 24667
rect 13461 24633 13495 24667
rect 25145 24633 25179 24667
rect 5825 24565 5859 24599
rect 8861 24565 8895 24599
rect 14841 24565 14875 24599
rect 16405 24565 16439 24599
rect 18061 24565 18095 24599
rect 20269 24565 20303 24599
rect 3249 24361 3283 24395
rect 3433 24361 3467 24395
rect 5733 24361 5767 24395
rect 6193 24361 6227 24395
rect 8769 24361 8803 24395
rect 13645 24361 13679 24395
rect 17601 24361 17635 24395
rect 4261 24225 4295 24259
rect 10057 24225 10091 24259
rect 11345 24225 11379 24259
rect 12541 24225 12575 24259
rect 13185 24225 13219 24259
rect 16865 24225 16899 24259
rect 17049 24225 17083 24259
rect 18245 24225 18279 24259
rect 19717 24225 19751 24259
rect 23857 24225 23891 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 2973 24157 3007 24191
rect 3985 24157 4019 24191
rect 6377 24157 6411 24191
rect 11161 24157 11195 24191
rect 11253 24157 11287 24191
rect 16773 24157 16807 24191
rect 17785 24157 17819 24191
rect 22017 24157 22051 24191
rect 22753 24157 22787 24191
rect 25053 24157 25087 24191
rect 2697 24089 2731 24123
rect 6745 24089 6779 24123
rect 9873 24089 9907 24123
rect 12357 24089 12391 24123
rect 14289 24089 14323 24123
rect 19993 24089 20027 24123
rect 24961 24089 24995 24123
rect 2053 24021 2087 24055
rect 9413 24021 9447 24055
rect 9781 24021 9815 24055
rect 10425 24021 10459 24055
rect 10793 24021 10827 24055
rect 11989 24021 12023 24055
rect 12449 24021 12483 24055
rect 16405 24021 16439 24055
rect 18061 24021 18095 24055
rect 21465 24021 21499 24055
rect 22109 24021 22143 24055
rect 24593 24021 24627 24055
rect 6009 23817 6043 23851
rect 6469 23817 6503 23851
rect 11805 23817 11839 23851
rect 12449 23817 12483 23851
rect 13921 23817 13955 23851
rect 25145 23817 25179 23851
rect 9873 23749 9907 23783
rect 23213 23749 23247 23783
rect 1777 23681 1811 23715
rect 7665 23681 7699 23715
rect 10333 23681 10367 23715
rect 21189 23681 21223 23715
rect 21557 23681 21591 23715
rect 22937 23681 22971 23715
rect 25329 23681 25363 23715
rect 2053 23613 2087 23647
rect 4261 23613 4295 23647
rect 4537 23613 4571 23647
rect 7941 23613 7975 23647
rect 10885 23613 10919 23647
rect 12173 23613 12207 23647
rect 12541 23613 12575 23647
rect 17049 23613 17083 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 20821 23613 20855 23647
rect 11621 23545 11655 23579
rect 9413 23477 9447 23511
rect 24685 23477 24719 23511
rect 2053 23273 2087 23307
rect 3157 23273 3191 23307
rect 7573 23273 7607 23307
rect 7941 23273 7975 23307
rect 16037 23273 16071 23307
rect 21189 23273 21223 23307
rect 21465 23273 21499 23307
rect 18245 23205 18279 23239
rect 2973 23137 3007 23171
rect 5825 23137 5859 23171
rect 11989 23137 12023 23171
rect 12725 23137 12759 23171
rect 13553 23137 13587 23171
rect 14289 23137 14323 23171
rect 16497 23137 16531 23171
rect 19441 23137 19475 23171
rect 22017 23137 22051 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 2789 23069 2823 23103
rect 4112 23069 4146 23103
rect 4215 23069 4249 23103
rect 9965 23069 9999 23103
rect 11713 23069 11747 23103
rect 12541 23069 12575 23103
rect 13461 23069 13495 23103
rect 22753 23069 22787 23103
rect 23857 23069 23891 23103
rect 24961 23069 24995 23103
rect 6101 23001 6135 23035
rect 10701 23001 10735 23035
rect 13369 23001 13403 23035
rect 14565 23001 14599 23035
rect 16773 23001 16807 23035
rect 19717 23001 19751 23035
rect 25053 23001 25087 23035
rect 11345 22933 11379 22967
rect 11805 22933 11839 22967
rect 13001 22933 13035 22967
rect 18613 22933 18647 22967
rect 24593 22933 24627 22967
rect 2053 22729 2087 22763
rect 5641 22729 5675 22763
rect 6837 22729 6871 22763
rect 7205 22729 7239 22763
rect 9321 22729 9355 22763
rect 10793 22729 10827 22763
rect 15209 22729 15243 22763
rect 16221 22729 16255 22763
rect 17509 22729 17543 22763
rect 23765 22729 23799 22763
rect 24225 22729 24259 22763
rect 24317 22729 24351 22763
rect 24777 22729 24811 22763
rect 25421 22729 25455 22763
rect 8033 22661 8067 22695
rect 10149 22661 10183 22695
rect 10885 22661 10919 22695
rect 13277 22661 13311 22695
rect 16405 22661 16439 22695
rect 17877 22661 17911 22695
rect 18613 22661 18647 22695
rect 19717 22661 19751 22695
rect 20545 22661 20579 22695
rect 2237 22593 2271 22627
rect 5733 22593 5767 22627
rect 11621 22593 11655 22627
rect 12357 22593 12391 22627
rect 13093 22593 13127 22627
rect 15117 22593 15151 22627
rect 19625 22593 19659 22627
rect 21373 22593 21407 22627
rect 22017 22593 22051 22627
rect 5917 22525 5951 22559
rect 7297 22525 7331 22559
rect 7481 22525 7515 22559
rect 8861 22525 8895 22559
rect 10977 22525 11011 22559
rect 12449 22525 12483 22559
rect 12633 22525 12667 22559
rect 13921 22525 13955 22559
rect 15393 22525 15427 22559
rect 19809 22525 19843 22559
rect 22293 22525 22327 22559
rect 10425 22457 10459 22491
rect 5273 22389 5307 22423
rect 11989 22389 12023 22423
rect 14749 22389 14783 22423
rect 19257 22389 19291 22423
rect 16405 22185 16439 22219
rect 19698 22185 19732 22219
rect 21465 22185 21499 22219
rect 11437 22117 11471 22151
rect 18061 22117 18095 22151
rect 11989 22049 12023 22083
rect 14289 22049 14323 22083
rect 16037 22049 16071 22083
rect 17509 22049 17543 22083
rect 18521 22049 18555 22083
rect 18705 22049 18739 22083
rect 22017 22049 22051 22083
rect 24041 22049 24075 22083
rect 11805 21981 11839 22015
rect 13277 21981 13311 22015
rect 16589 21981 16623 22015
rect 17233 21981 17267 22015
rect 19441 21981 19475 22015
rect 24869 21981 24903 22015
rect 11897 21913 11931 21947
rect 12541 21913 12575 21947
rect 14565 21913 14599 21947
rect 18429 21913 18463 21947
rect 22293 21913 22327 21947
rect 24685 21913 24719 21947
rect 4445 21845 4479 21879
rect 10885 21845 10919 21879
rect 11161 21845 11195 21879
rect 13093 21845 13127 21879
rect 16865 21845 16899 21879
rect 17325 21845 17359 21879
rect 21189 21845 21223 21879
rect 7113 21641 7147 21675
rect 7481 21641 7515 21675
rect 8309 21641 8343 21675
rect 8677 21641 8711 21675
rect 9873 21641 9907 21675
rect 11713 21641 11747 21675
rect 12081 21641 12115 21675
rect 13553 21641 13587 21675
rect 13921 21641 13955 21675
rect 18521 21641 18555 21675
rect 22569 21641 22603 21675
rect 25421 21641 25455 21675
rect 14013 21573 14047 21607
rect 23673 21573 23707 21607
rect 1777 21505 1811 21539
rect 3433 21505 3467 21539
rect 4537 21505 4571 21539
rect 7573 21505 7607 21539
rect 12173 21505 12207 21539
rect 15209 21505 15243 21539
rect 16221 21505 16255 21539
rect 17049 21505 17083 21539
rect 18705 21505 18739 21539
rect 22477 21505 22511 21539
rect 23397 21505 23431 21539
rect 2053 21437 2087 21471
rect 3617 21437 3651 21471
rect 4997 21437 5031 21471
rect 7665 21437 7699 21471
rect 8769 21437 8803 21471
rect 8861 21437 8895 21471
rect 9965 21437 9999 21471
rect 10057 21437 10091 21471
rect 12357 21437 12391 21471
rect 14197 21437 14231 21471
rect 15301 21437 15335 21471
rect 15393 21437 15427 21471
rect 17693 21437 17727 21471
rect 22753 21437 22787 21471
rect 25145 21437 25179 21471
rect 3801 21369 3835 21403
rect 9505 21369 9539 21403
rect 16865 21369 16899 21403
rect 4813 21301 4847 21335
rect 14841 21301 14875 21335
rect 16037 21301 16071 21335
rect 20453 21301 20487 21335
rect 22109 21301 22143 21335
rect 3157 21097 3191 21131
rect 7849 21097 7883 21131
rect 16313 21097 16347 21131
rect 16957 21097 16991 21131
rect 21925 21097 21959 21131
rect 4077 21029 4111 21063
rect 14381 21029 14415 21063
rect 16129 21029 16163 21063
rect 2789 20961 2823 20995
rect 8401 20961 8435 20995
rect 9781 20961 9815 20995
rect 13829 20961 13863 20995
rect 14933 20961 14967 20995
rect 17693 20961 17727 20995
rect 17877 20961 17911 20995
rect 19901 20961 19935 20995
rect 20177 20961 20211 20995
rect 23857 20961 23891 20995
rect 2237 20893 2271 20927
rect 2973 20893 3007 20927
rect 4261 20893 4295 20927
rect 11897 20893 11931 20927
rect 13737 20893 13771 20927
rect 14841 20893 14875 20927
rect 15761 20893 15795 20927
rect 17601 20893 17635 20927
rect 18889 20893 18923 20927
rect 22845 20893 22879 20927
rect 10057 20825 10091 20859
rect 14749 20825 14783 20859
rect 2053 20757 2087 20791
rect 7481 20757 7515 20791
rect 8217 20757 8251 20791
rect 8309 20757 8343 20791
rect 11529 20757 11563 20791
rect 15577 20757 15611 20791
rect 17233 20757 17267 20791
rect 18705 20757 18739 20791
rect 21649 20757 21683 20791
rect 9965 20553 9999 20587
rect 17325 20553 17359 20587
rect 19441 20553 19475 20587
rect 4261 20485 4295 20519
rect 6009 20485 6043 20519
rect 10425 20485 10459 20519
rect 17693 20485 17727 20519
rect 23305 20485 23339 20519
rect 3985 20417 4019 20451
rect 6561 20417 6595 20451
rect 9137 20417 9171 20451
rect 10333 20417 10367 20451
rect 12449 20417 12483 20451
rect 13277 20417 13311 20451
rect 15669 20417 15703 20451
rect 18521 20417 18555 20451
rect 19349 20417 19383 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 6837 20349 6871 20383
rect 9229 20349 9263 20383
rect 9321 20349 9355 20383
rect 10517 20349 10551 20383
rect 12541 20349 12575 20383
rect 12725 20349 12759 20383
rect 19625 20349 19659 20383
rect 24409 20349 24443 20383
rect 8769 20281 8803 20315
rect 14657 20281 14691 20315
rect 15485 20281 15519 20315
rect 5733 20213 5767 20247
rect 8309 20213 8343 20247
rect 12081 20213 12115 20247
rect 13737 20213 13771 20247
rect 17785 20213 17819 20247
rect 18337 20213 18371 20247
rect 18981 20213 19015 20247
rect 5089 20009 5123 20043
rect 11713 20009 11747 20043
rect 14289 20009 14323 20043
rect 20269 20009 20303 20043
rect 15393 19941 15427 19975
rect 5733 19873 5767 19907
rect 6009 19873 6043 19907
rect 9137 19873 9171 19907
rect 11161 19873 11195 19907
rect 12265 19873 12299 19907
rect 14841 19873 14875 19907
rect 23857 19873 23891 19907
rect 5273 19805 5307 19839
rect 7757 19805 7791 19839
rect 8401 19805 8435 19839
rect 12081 19805 12115 19839
rect 14657 19805 14691 19839
rect 17233 19805 17267 19839
rect 17785 19805 17819 19839
rect 18705 19805 18739 19839
rect 22017 19805 22051 19839
rect 22845 19805 22879 19839
rect 9413 19737 9447 19771
rect 12173 19737 12207 19771
rect 17325 19737 17359 19771
rect 17969 19737 18003 19771
rect 22201 19737 22235 19771
rect 7481 19669 7515 19703
rect 8677 19669 8711 19703
rect 13921 19669 13955 19703
rect 14749 19669 14783 19703
rect 18521 19669 18555 19703
rect 19349 19669 19383 19703
rect 2053 19465 2087 19499
rect 4261 19465 4295 19499
rect 8769 19465 8803 19499
rect 9229 19465 9263 19499
rect 11713 19465 11747 19499
rect 12081 19465 12115 19499
rect 13277 19465 13311 19499
rect 14013 19465 14047 19499
rect 16865 19465 16899 19499
rect 17509 19465 17543 19499
rect 19901 19465 19935 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 23765 19465 23799 19499
rect 17877 19397 17911 19431
rect 18797 19397 18831 19431
rect 2237 19329 2271 19363
rect 4445 19329 4479 19363
rect 6561 19329 6595 19363
rect 9137 19329 9171 19363
rect 12173 19329 12207 19363
rect 13921 19329 13955 19363
rect 17049 19329 17083 19363
rect 19809 19329 19843 19363
rect 21097 19329 21131 19363
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 11253 19261 11287 19295
rect 12265 19261 12299 19295
rect 14105 19261 14139 19295
rect 17969 19261 18003 19295
rect 18153 19261 18187 19295
rect 20085 19261 20119 19295
rect 21373 19261 21407 19295
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 14749 19193 14783 19227
rect 18981 19193 19015 19227
rect 8309 19125 8343 19159
rect 10885 19125 10919 19159
rect 11069 19125 11103 19159
rect 13553 19125 13587 19159
rect 14657 19125 14691 19159
rect 19441 19125 19475 19159
rect 24133 19125 24167 19159
rect 11897 18921 11931 18955
rect 12173 18921 12207 18955
rect 14289 18921 14323 18955
rect 18337 18921 18371 18955
rect 19073 18921 19107 18955
rect 24041 18921 24075 18955
rect 24409 18921 24443 18955
rect 8953 18853 8987 18887
rect 2053 18785 2087 18819
rect 9413 18785 9447 18819
rect 10057 18785 10091 18819
rect 13553 18785 13587 18819
rect 14841 18785 14875 18819
rect 17969 18785 18003 18819
rect 1777 18717 1811 18751
rect 9781 18717 9815 18751
rect 13461 18717 13495 18751
rect 14657 18717 14691 18751
rect 16221 18717 16255 18751
rect 19625 18717 19659 18751
rect 20361 18717 20395 18751
rect 21557 18717 21591 18751
rect 22293 18717 22327 18751
rect 9229 18649 9263 18683
rect 16497 18649 16531 18683
rect 18521 18649 18555 18683
rect 21097 18649 21131 18683
rect 22569 18649 22603 18683
rect 8493 18581 8527 18615
rect 8677 18581 8711 18615
rect 11529 18581 11563 18615
rect 13001 18581 13035 18615
rect 13369 18581 13403 18615
rect 14749 18581 14783 18615
rect 19717 18581 19751 18615
rect 7757 18377 7791 18411
rect 9781 18377 9815 18411
rect 10425 18377 10459 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 14657 18377 14691 18411
rect 15393 18377 15427 18411
rect 8493 18309 8527 18343
rect 12081 18309 12115 18343
rect 13645 18309 13679 18343
rect 17233 18309 17267 18343
rect 17509 18309 17543 18343
rect 19165 18309 19199 18343
rect 21281 18309 21315 18343
rect 7665 18241 7699 18275
rect 13921 18241 13955 18275
rect 22109 18241 22143 18275
rect 23949 18241 23983 18275
rect 7849 18173 7883 18207
rect 9229 18173 9263 18207
rect 10149 18173 10183 18207
rect 10885 18173 10919 18207
rect 10977 18173 11011 18207
rect 12173 18173 12207 18207
rect 12357 18173 12391 18207
rect 14749 18173 14783 18207
rect 14933 18173 14967 18207
rect 18337 18173 18371 18207
rect 18889 18173 18923 18207
rect 23305 18173 23339 18207
rect 24777 18173 24811 18207
rect 11713 18105 11747 18139
rect 21465 18105 21499 18139
rect 6929 18037 6963 18071
rect 7297 18037 7331 18071
rect 13829 18037 13863 18071
rect 20637 18037 20671 18071
rect 6285 17833 6319 17867
rect 9137 17833 9171 17867
rect 12541 17833 12575 17867
rect 21649 17833 21683 17867
rect 23857 17833 23891 17867
rect 24225 17833 24259 17867
rect 16221 17765 16255 17799
rect 6837 17697 6871 17731
rect 7941 17697 7975 17731
rect 8125 17697 8159 17731
rect 9689 17697 9723 17731
rect 11897 17697 11931 17731
rect 12725 17697 12759 17731
rect 13553 17697 13587 17731
rect 14841 17697 14875 17731
rect 16681 17697 16715 17731
rect 16865 17697 16899 17731
rect 19901 17697 19935 17731
rect 22109 17697 22143 17731
rect 22385 17697 22419 17731
rect 10517 17629 10551 17663
rect 13461 17629 13495 17663
rect 15577 17629 15611 17663
rect 17233 17629 17267 17663
rect 24869 17629 24903 17663
rect 6653 17561 6687 17595
rect 11345 17561 11379 17595
rect 13369 17561 13403 17595
rect 20177 17561 20211 17595
rect 6745 17493 6779 17527
rect 7481 17493 7515 17527
rect 7849 17493 7883 17527
rect 8769 17493 8803 17527
rect 9505 17493 9539 17527
rect 9597 17493 9631 17527
rect 13001 17493 13035 17527
rect 14289 17493 14323 17527
rect 14657 17493 14691 17527
rect 14749 17493 14783 17527
rect 15669 17493 15703 17527
rect 16589 17493 16623 17527
rect 24685 17493 24719 17527
rect 10057 17289 10091 17323
rect 11529 17289 11563 17323
rect 16037 17289 16071 17323
rect 8585 17221 8619 17255
rect 10425 17221 10459 17255
rect 12909 17221 12943 17255
rect 14933 17221 14967 17255
rect 19717 17221 19751 17255
rect 21005 17221 21039 17255
rect 21557 17221 21591 17255
rect 22845 17221 22879 17255
rect 9045 17153 9079 17187
rect 14841 17153 14875 17187
rect 17049 17153 17083 17187
rect 17693 17153 17727 17187
rect 22109 17153 22143 17187
rect 23949 17153 23983 17187
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 9505 17085 9539 17119
rect 10517 17085 10551 17119
rect 10701 17085 10735 17119
rect 12633 17085 12667 17119
rect 14381 17085 14415 17119
rect 17969 17085 18003 17119
rect 19441 17085 19475 17119
rect 20453 17085 20487 17119
rect 24685 17085 24719 17119
rect 15209 17017 15243 17051
rect 22293 17017 22327 17051
rect 23029 17017 23063 17051
rect 9321 16949 9355 16983
rect 16865 16949 16899 16983
rect 5628 16745 5662 16779
rect 7113 16745 7147 16779
rect 7481 16745 7515 16779
rect 9137 16745 9171 16779
rect 10517 16745 10551 16779
rect 23857 16745 23891 16779
rect 8677 16677 8711 16711
rect 10241 16677 10275 16711
rect 19349 16677 19383 16711
rect 5365 16609 5399 16643
rect 7665 16609 7699 16643
rect 9689 16609 9723 16643
rect 10977 16609 11011 16643
rect 11069 16609 11103 16643
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 15025 16609 15059 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 20637 16609 20671 16643
rect 21741 16609 21775 16643
rect 22017 16609 22051 16643
rect 1593 16541 1627 16575
rect 9505 16541 9539 16575
rect 10885 16541 10919 16575
rect 12173 16541 12207 16575
rect 20453 16541 20487 16575
rect 20545 16541 20579 16575
rect 2513 16473 2547 16507
rect 8493 16405 8527 16439
rect 9597 16405 9631 16439
rect 11805 16405 11839 16439
rect 15301 16405 15335 16439
rect 15669 16405 15703 16439
rect 16405 16405 16439 16439
rect 20085 16405 20119 16439
rect 23489 16405 23523 16439
rect 8953 16201 8987 16235
rect 10149 16201 10183 16235
rect 10609 16201 10643 16235
rect 11713 16201 11747 16235
rect 13093 16201 13127 16235
rect 13737 16201 13771 16235
rect 14749 16201 14783 16235
rect 18613 16201 18647 16235
rect 19257 16201 19291 16235
rect 22477 16201 22511 16235
rect 23213 16201 23247 16235
rect 2513 16133 2547 16167
rect 9321 16133 9355 16167
rect 12081 16133 12115 16167
rect 14197 16133 14231 16167
rect 15945 16133 15979 16167
rect 16405 16133 16439 16167
rect 17141 16133 17175 16167
rect 18889 16133 18923 16167
rect 19717 16133 19751 16167
rect 21281 16133 21315 16167
rect 6653 16065 6687 16099
rect 10517 16065 10551 16099
rect 12173 16065 12207 16099
rect 16865 16065 16899 16099
rect 19625 16065 19659 16099
rect 20453 16065 20487 16099
rect 22385 16065 22419 16099
rect 23397 16065 23431 16099
rect 24133 16065 24167 16099
rect 6929 15997 6963 16031
rect 8401 15997 8435 16031
rect 9413 15997 9447 16031
rect 9505 15997 9539 16031
rect 10701 15997 10735 16031
rect 12265 15997 12299 16031
rect 19901 15997 19935 16031
rect 22569 15997 22603 16031
rect 24777 15997 24811 16031
rect 21465 15929 21499 15963
rect 2605 15861 2639 15895
rect 14289 15861 14323 15895
rect 16037 15861 16071 15895
rect 22017 15861 22051 15895
rect 8769 15657 8803 15691
rect 9965 15657 9999 15691
rect 13553 15657 13587 15691
rect 14289 15657 14323 15691
rect 17325 15589 17359 15623
rect 11069 15521 11103 15555
rect 14841 15521 14875 15555
rect 17877 15521 17911 15555
rect 20085 15521 20119 15555
rect 13461 15453 13495 15487
rect 14657 15453 14691 15487
rect 17785 15453 17819 15487
rect 18337 15453 18371 15487
rect 19809 15453 19843 15487
rect 20821 15453 20855 15487
rect 22845 15453 22879 15487
rect 11345 15385 11379 15419
rect 21097 15385 21131 15419
rect 21833 15385 21867 15419
rect 23857 15385 23891 15419
rect 8493 15317 8527 15351
rect 10241 15317 10275 15351
rect 10793 15317 10827 15351
rect 12817 15317 12851 15351
rect 14749 15317 14783 15351
rect 17049 15317 17083 15351
rect 17693 15317 17727 15351
rect 18705 15317 18739 15351
rect 19441 15317 19475 15351
rect 19901 15317 19935 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 13001 15113 13035 15147
rect 14197 15113 14231 15147
rect 18797 15113 18831 15147
rect 18889 15113 18923 15147
rect 22293 15113 22327 15147
rect 9413 15045 9447 15079
rect 12725 15045 12759 15079
rect 13461 15045 13495 15079
rect 17233 15045 17267 15079
rect 17693 15045 17727 15079
rect 13369 14977 13403 15011
rect 14565 14977 14599 15011
rect 14657 14977 14691 15011
rect 15669 14977 15703 15011
rect 16129 14977 16163 15011
rect 19809 14977 19843 15011
rect 23949 14977 23983 15011
rect 9137 14909 9171 14943
rect 11161 14909 11195 14943
rect 13645 14909 13679 14943
rect 14841 14909 14875 14943
rect 15301 14909 15335 14943
rect 18981 14909 19015 14943
rect 24685 14909 24719 14943
rect 15853 14841 15887 14875
rect 17417 14841 17451 14875
rect 11529 14773 11563 14807
rect 18429 14773 18463 14807
rect 19625 14773 19659 14807
rect 20085 14773 20119 14807
rect 13001 14569 13035 14603
rect 17141 14569 17175 14603
rect 23029 14569 23063 14603
rect 11989 14501 12023 14535
rect 14105 14501 14139 14535
rect 9965 14433 9999 14467
rect 12541 14433 12575 14467
rect 13461 14433 13495 14467
rect 13645 14433 13679 14467
rect 15393 14433 15427 14467
rect 21189 14433 21223 14467
rect 12725 14365 12759 14399
rect 18245 14365 18279 14399
rect 18613 14365 18647 14399
rect 19441 14365 19475 14399
rect 20913 14365 20947 14399
rect 10241 14297 10275 14331
rect 13369 14297 13403 14331
rect 15669 14297 15703 14331
rect 18797 14297 18831 14331
rect 11713 14229 11747 14263
rect 14381 14229 14415 14263
rect 14565 14229 14599 14263
rect 17509 14229 17543 14263
rect 19993 14229 20027 14263
rect 22661 14229 22695 14263
rect 12265 14025 12299 14059
rect 13645 14025 13679 14059
rect 18889 14025 18923 14059
rect 21833 14025 21867 14059
rect 23029 14025 23063 14059
rect 17417 13957 17451 13991
rect 19901 13957 19935 13991
rect 21373 13957 21407 13991
rect 25145 13957 25179 13991
rect 1777 13889 1811 13923
rect 8033 13889 8067 13923
rect 10057 13889 10091 13923
rect 12633 13889 12667 13923
rect 13553 13889 13587 13923
rect 14013 13889 14047 13923
rect 17141 13889 17175 13923
rect 19717 13889 19751 13923
rect 20453 13889 20487 13923
rect 21189 13889 21223 13923
rect 23213 13889 23247 13923
rect 23949 13889 23983 13923
rect 2053 13821 2087 13855
rect 9781 13821 9815 13855
rect 11897 13821 11931 13855
rect 12725 13821 12759 13855
rect 12909 13821 12943 13855
rect 19257 13821 19291 13855
rect 20637 13821 20671 13855
rect 8296 13685 8330 13719
rect 7100 13481 7134 13515
rect 8953 13481 8987 13515
rect 11621 13481 11655 13515
rect 12357 13481 12391 13515
rect 13369 13481 13403 13515
rect 16313 13481 16347 13515
rect 20729 13481 20763 13515
rect 18797 13413 18831 13447
rect 19441 13413 19475 13447
rect 9137 13345 9171 13379
rect 9873 13345 9907 13379
rect 12909 13345 12943 13379
rect 14565 13345 14599 13379
rect 18245 13345 18279 13379
rect 18429 13345 18463 13379
rect 20085 13345 20119 13379
rect 6837 13277 6871 13311
rect 12725 13277 12759 13311
rect 17509 13277 17543 13311
rect 18153 13277 18187 13311
rect 19809 13277 19843 13311
rect 22661 13277 22695 13311
rect 10149 13209 10183 13243
rect 12817 13209 12851 13243
rect 14841 13209 14875 13243
rect 23857 13209 23891 13243
rect 8585 13141 8619 13175
rect 11989 13141 12023 13175
rect 16865 13141 16899 13175
rect 17785 13141 17819 13175
rect 19901 13141 19935 13175
rect 21649 13141 21683 13175
rect 8677 12937 8711 12971
rect 11161 12937 11195 12971
rect 13277 12937 13311 12971
rect 14933 12937 14967 12971
rect 16129 12937 16163 12971
rect 16497 12937 16531 12971
rect 17233 12937 17267 12971
rect 17325 12937 17359 12971
rect 19073 12937 19107 12971
rect 21465 12937 21499 12971
rect 11529 12869 11563 12903
rect 14473 12869 14507 12903
rect 15393 12869 15427 12903
rect 15853 12869 15887 12903
rect 18521 12869 18555 12903
rect 8585 12801 8619 12835
rect 9413 12801 9447 12835
rect 13737 12801 13771 12835
rect 22845 12801 22879 12835
rect 23949 12801 23983 12835
rect 8769 12733 8803 12767
rect 9689 12733 9723 12767
rect 17417 12733 17451 12767
rect 19717 12733 19751 12767
rect 19993 12733 20027 12767
rect 22017 12733 22051 12767
rect 24777 12733 24811 12767
rect 13921 12665 13955 12699
rect 14657 12665 14691 12699
rect 16865 12665 16899 12699
rect 8217 12597 8251 12631
rect 15485 12597 15519 12631
rect 18613 12597 18647 12631
rect 22661 12597 22695 12631
rect 14105 12393 14139 12427
rect 14473 12393 14507 12427
rect 15669 12393 15703 12427
rect 18889 12393 18923 12427
rect 21097 12325 21131 12359
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 13921 12257 13955 12291
rect 15117 12257 15151 12291
rect 16221 12257 16255 12291
rect 17141 12257 17175 12291
rect 17417 12257 17451 12291
rect 21557 12257 21591 12291
rect 21741 12257 21775 12291
rect 13737 12189 13771 12223
rect 14933 12189 14967 12223
rect 16037 12189 16071 12223
rect 20637 12189 20671 12223
rect 21465 12189 21499 12223
rect 23397 12189 23431 12223
rect 14841 12121 14875 12155
rect 13277 12053 13311 12087
rect 16129 12053 16163 12087
rect 19349 12053 19383 12087
rect 20453 12053 20487 12087
rect 23213 12053 23247 12087
rect 14565 11849 14599 11883
rect 15485 11849 15519 11883
rect 16129 11849 16163 11883
rect 17509 11849 17543 11883
rect 19993 11849 20027 11883
rect 20361 11849 20395 11883
rect 24225 11849 24259 11883
rect 16957 11781 16991 11815
rect 18521 11781 18555 11815
rect 20913 11781 20947 11815
rect 21373 11781 21407 11815
rect 12817 11713 12851 11747
rect 15393 11713 15427 11747
rect 18245 11713 18279 11747
rect 22937 11713 22971 11747
rect 13093 11645 13127 11679
rect 15577 11645 15611 11679
rect 21097 11645 21131 11679
rect 15025 11509 15059 11543
rect 17049 11509 17083 11543
rect 15485 11305 15519 11339
rect 14749 11169 14783 11203
rect 16037 11169 16071 11203
rect 15853 11033 15887 11067
rect 20821 11033 20855 11067
rect 21005 11033 21039 11067
rect 15945 10965 15979 10999
rect 19625 10965 19659 10999
rect 14657 10761 14691 10795
rect 19533 10761 19567 10795
rect 20361 10761 20395 10795
rect 12081 10693 12115 10727
rect 12541 10693 12575 10727
rect 15393 10693 15427 10727
rect 14841 10625 14875 10659
rect 18429 10625 18463 10659
rect 19625 10625 19659 10659
rect 20545 10625 20579 10659
rect 23397 10625 23431 10659
rect 23949 10625 23983 10659
rect 19717 10557 19751 10591
rect 24777 10557 24811 10591
rect 12265 10489 12299 10523
rect 15209 10489 15243 10523
rect 18245 10421 18279 10455
rect 19165 10421 19199 10455
rect 23213 10421 23247 10455
rect 21281 10149 21315 10183
rect 14657 10013 14691 10047
rect 14841 10013 14875 10047
rect 21465 10013 21499 10047
rect 22201 10013 22235 10047
rect 22661 10013 22695 10047
rect 23857 10013 23891 10047
rect 16773 9945 16807 9979
rect 16957 9945 16991 9979
rect 24685 9945 24719 9979
rect 22017 9877 22051 9911
rect 24777 9877 24811 9911
rect 16957 9605 16991 9639
rect 5825 9537 5859 9571
rect 6929 9537 6963 9571
rect 19257 9537 19291 9571
rect 22937 9537 22971 9571
rect 23949 9537 23983 9571
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 24685 9469 24719 9503
rect 6561 9401 6595 9435
rect 17141 9401 17175 9435
rect 19073 9333 19107 9367
rect 22753 9333 22787 9367
rect 24685 9061 24719 9095
rect 21741 8925 21775 8959
rect 23949 8925 23983 8959
rect 24869 8925 24903 8959
rect 21557 8789 21591 8823
rect 23765 8789 23799 8823
rect 19165 8517 19199 8551
rect 19625 8517 19659 8551
rect 20729 8517 20763 8551
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 19349 8381 19383 8415
rect 22569 8381 22603 8415
rect 24593 8381 24627 8415
rect 20913 8313 20947 8347
rect 6653 8041 6687 8075
rect 25237 8041 25271 8075
rect 4077 7905 4111 7939
rect 6101 7905 6135 7939
rect 6469 7905 6503 7939
rect 23397 7905 23431 7939
rect 20453 7837 20487 7871
rect 21281 7837 21315 7871
rect 22845 7837 22879 7871
rect 24593 7837 24627 7871
rect 4353 7769 4387 7803
rect 20269 7701 20303 7735
rect 21097 7701 21131 7735
rect 18797 7429 18831 7463
rect 20269 7361 20303 7395
rect 22109 7361 22143 7395
rect 23949 7361 23983 7395
rect 21281 7293 21315 7327
rect 22569 7293 22603 7327
rect 24685 7293 24719 7327
rect 18981 7225 19015 7259
rect 19717 6749 19751 6783
rect 19993 6749 20027 6783
rect 20821 6749 20855 6783
rect 22845 6749 22879 6783
rect 24869 6749 24903 6783
rect 22017 6681 22051 6715
rect 23857 6681 23891 6715
rect 19533 6613 19567 6647
rect 24685 6613 24719 6647
rect 3709 6409 3743 6443
rect 17969 6409 18003 6443
rect 3065 6273 3099 6307
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 23949 6273 23983 6307
rect 19257 6205 19291 6239
rect 21281 6205 21315 6239
rect 22477 6205 22511 6239
rect 24593 6205 24627 6239
rect 24777 5865 24811 5899
rect 21005 5729 21039 5763
rect 22845 5729 22879 5763
rect 17693 5661 17727 5695
rect 20545 5661 20579 5695
rect 22385 5661 22419 5695
rect 24685 5661 24719 5695
rect 18705 5593 18739 5627
rect 1593 5321 1627 5355
rect 18797 5253 18831 5287
rect 1777 5185 1811 5219
rect 17785 5185 17819 5219
rect 19533 5185 19567 5219
rect 22017 5185 22051 5219
rect 24041 5185 24075 5219
rect 19901 5117 19935 5151
rect 22477 5117 22511 5151
rect 24777 5117 24811 5151
rect 23857 4777 23891 4811
rect 2053 4709 2087 4743
rect 24869 4709 24903 4743
rect 19901 4641 19935 4675
rect 21741 4641 21775 4675
rect 17693 4573 17727 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 24041 4573 24075 4607
rect 1869 4505 1903 4539
rect 2329 4505 2363 4539
rect 18705 4505 18739 4539
rect 24685 4505 24719 4539
rect 2421 4233 2455 4267
rect 25145 4165 25179 4199
rect 1777 4097 1811 4131
rect 2881 4097 2915 4131
rect 3433 4097 3467 4131
rect 13645 4097 13679 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 18797 4097 18831 4131
rect 22109 4097 22143 4131
rect 24133 4097 24167 4131
rect 11345 4029 11379 4063
rect 11713 4029 11747 4063
rect 11989 4029 12023 4063
rect 14013 4029 14047 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 3065 3961 3099 3995
rect 9965 3961 9999 3995
rect 6377 3893 6411 3927
rect 9505 3893 9539 3927
rect 9781 3893 9815 3927
rect 11069 3893 11103 3927
rect 16221 3893 16255 3927
rect 1961 3689 1995 3723
rect 2697 3689 2731 3723
rect 3249 3689 3283 3723
rect 6745 3689 6779 3723
rect 8217 3689 8251 3723
rect 9321 3689 9355 3723
rect 10057 3689 10091 3723
rect 18613 3689 18647 3723
rect 5273 3621 5307 3655
rect 5917 3621 5951 3655
rect 11253 3553 11287 3587
rect 12817 3553 12851 3587
rect 15485 3553 15519 3587
rect 17325 3553 17359 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 1501 3485 1535 3519
rect 1777 3485 1811 3519
rect 2513 3485 2547 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 5089 3485 5123 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 7757 3485 7791 3519
rect 8033 3485 8067 3519
rect 9137 3485 9171 3519
rect 9873 3485 9907 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 12449 3485 12483 3519
rect 15117 3485 15151 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 21281 3485 21315 3519
rect 23397 3485 23431 3519
rect 24041 3485 24075 3519
rect 24593 3485 24627 3519
rect 7573 3417 7607 3451
rect 4813 3349 4847 3383
rect 7205 3349 7239 3383
rect 8677 3349 8711 3383
rect 10701 3349 10735 3383
rect 25237 3349 25271 3383
rect 2237 3145 2271 3179
rect 2881 3145 2915 3179
rect 5181 3145 5215 3179
rect 5917 3145 5951 3179
rect 6469 3145 6503 3179
rect 7021 3145 7055 3179
rect 7757 3145 7791 3179
rect 8493 3145 8527 3179
rect 11897 3145 11931 3179
rect 25145 3145 25179 3179
rect 1593 3009 1627 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9045 3009 9079 3043
rect 9321 3009 9355 3043
rect 10333 3009 10367 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 12633 3009 12667 3043
rect 14289 3009 14323 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 25329 3009 25363 3043
rect 2789 2941 2823 2975
rect 3249 2941 3283 2975
rect 3525 2941 3559 2975
rect 13369 2941 13403 2975
rect 14749 2941 14783 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 4353 2805 4387 2839
rect 24133 2805 24167 2839
rect 2237 2601 2271 2635
rect 3341 2601 3375 2635
rect 4169 2601 4203 2635
rect 7113 2601 7147 2635
rect 9781 2601 9815 2635
rect 11713 2601 11747 2635
rect 18613 2601 18647 2635
rect 25237 2601 25271 2635
rect 5825 2465 5859 2499
rect 7941 2465 7975 2499
rect 10609 2465 10643 2499
rect 14105 2465 14139 2499
rect 15209 2465 15243 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 24041 2465 24075 2499
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 3157 2397 3191 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 9137 2397 9171 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 16957 2397 16991 2431
rect 19441 2397 19475 2431
rect 22017 2397 22051 2431
rect 24593 2397 24627 2431
rect 6101 2329 6135 2363
rect 6653 2329 6687 2363
rect 9321 2329 9355 2363
rect 13553 2329 13587 2363
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 3970 54272 3976 54324
rect 4028 54272 4034 54324
rect 9950 54272 9956 54324
rect 10008 54272 10014 54324
rect 14553 54315 14611 54321
rect 14553 54281 14565 54315
rect 14599 54312 14611 54315
rect 14734 54312 14740 54324
rect 14599 54284 14740 54312
rect 14599 54281 14611 54284
rect 14553 54275 14611 54281
rect 14734 54272 14740 54284
rect 14792 54272 14798 54324
rect 16206 54272 16212 54324
rect 16264 54312 16270 54324
rect 16393 54315 16451 54321
rect 16393 54312 16405 54315
rect 16264 54284 16405 54312
rect 16264 54272 16270 54284
rect 16393 54281 16405 54284
rect 16439 54312 16451 54315
rect 16439 54284 16574 54312
rect 16439 54281 16451 54284
rect 16393 54275 16451 54281
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 7834 54244 7840 54256
rect 5859 54216 7840 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 7834 54204 7840 54216
rect 7892 54204 7898 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 9968 54244 9996 54272
rect 8435 54216 9996 54244
rect 10965 54247 11023 54253
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 12894 54244 12900 54256
rect 11900 54216 12900 54244
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 2314 54176 2320 54188
rect 2271 54148 2320 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 2314 54136 2320 54148
rect 2372 54136 2378 54188
rect 4801 54179 4859 54185
rect 4801 54145 4813 54179
rect 4847 54176 4859 54179
rect 5350 54176 5356 54188
rect 4847 54148 5356 54176
rect 4847 54145 4859 54148
rect 4801 54139 4859 54145
rect 5350 54136 5356 54148
rect 5408 54136 5414 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54145 7435 54179
rect 7377 54139 7435 54145
rect 3237 54111 3295 54117
rect 3237 54077 3249 54111
rect 3283 54108 3295 54111
rect 5902 54108 5908 54120
rect 3283 54080 5908 54108
rect 3283 54077 3295 54080
rect 3237 54071 3295 54077
rect 5902 54068 5908 54080
rect 5960 54068 5966 54120
rect 7392 54108 7420 54139
rect 9950 54136 9956 54188
rect 10008 54136 10014 54188
rect 11900 54185 11928 54216
rect 12894 54204 12900 54216
rect 12952 54244 12958 54256
rect 14093 54247 14151 54253
rect 14093 54244 14105 54247
rect 12952 54216 14105 54244
rect 12952 54204 12958 54216
rect 14093 54213 14105 54216
rect 14139 54213 14151 54247
rect 14093 54207 14151 54213
rect 11885 54179 11943 54185
rect 11885 54145 11897 54179
rect 11931 54145 11943 54179
rect 11885 54139 11943 54145
rect 12342 54136 12348 54188
rect 12400 54136 12406 54188
rect 14752 54176 14780 54272
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14752 54148 14841 54176
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 15194 54136 15200 54188
rect 15252 54176 15258 54188
rect 15565 54179 15623 54185
rect 15565 54176 15577 54179
rect 15252 54148 15577 54176
rect 15252 54136 15258 54148
rect 15565 54145 15577 54148
rect 15611 54176 15623 54179
rect 16117 54179 16175 54185
rect 16117 54176 16129 54179
rect 15611 54148 16129 54176
rect 15611 54145 15623 54148
rect 15565 54139 15623 54145
rect 16117 54145 16129 54148
rect 16163 54145 16175 54179
rect 16546 54176 16574 54284
rect 24486 54272 24492 54324
rect 24544 54272 24550 54324
rect 17678 54204 17684 54256
rect 17736 54244 17742 54256
rect 18417 54247 18475 54253
rect 18417 54244 18429 54247
rect 17736 54216 18429 54244
rect 17736 54204 17742 54216
rect 18417 54213 18429 54216
rect 18463 54244 18475 54247
rect 18874 54244 18880 54256
rect 18463 54216 18880 54244
rect 18463 54213 18475 54216
rect 18417 54207 18475 54213
rect 18874 54204 18880 54216
rect 18932 54204 18938 54256
rect 21453 54247 21511 54253
rect 21453 54244 21465 54247
rect 20180 54216 21465 54244
rect 16853 54179 16911 54185
rect 16853 54176 16865 54179
rect 16546 54148 16865 54176
rect 16117 54139 16175 54145
rect 16853 54145 16865 54148
rect 16899 54145 16911 54179
rect 16853 54139 16911 54145
rect 16942 54136 16948 54188
rect 17000 54176 17006 54188
rect 17589 54179 17647 54185
rect 17589 54176 17601 54179
rect 17000 54148 17601 54176
rect 17000 54136 17006 54148
rect 17589 54145 17601 54148
rect 17635 54176 17647 54179
rect 18969 54179 19027 54185
rect 18969 54176 18981 54179
rect 17635 54148 18981 54176
rect 17635 54145 17647 54148
rect 17589 54139 17647 54145
rect 18969 54145 18981 54148
rect 19015 54145 19027 54179
rect 18969 54139 19027 54145
rect 19429 54179 19487 54185
rect 19429 54145 19441 54179
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 11238 54108 11244 54120
rect 7392 54080 11244 54108
rect 11238 54068 11244 54080
rect 11296 54068 11302 54120
rect 12526 54068 12532 54120
rect 12584 54108 12590 54120
rect 12805 54111 12863 54117
rect 12805 54108 12817 54111
rect 12584 54080 12817 54108
rect 12584 54068 12590 54080
rect 12805 54077 12817 54080
rect 12851 54077 12863 54111
rect 12805 54071 12863 54077
rect 18414 54068 18420 54120
rect 18472 54108 18478 54120
rect 19444 54108 19472 54139
rect 19518 54136 19524 54188
rect 19576 54176 19582 54188
rect 20180 54185 20208 54216
rect 21453 54213 21465 54216
rect 21499 54213 21511 54247
rect 23293 54247 23351 54253
rect 23293 54244 23305 54247
rect 21453 54207 21511 54213
rect 22020 54216 23305 54244
rect 20165 54179 20223 54185
rect 20165 54176 20177 54179
rect 19576 54148 20177 54176
rect 19576 54136 19582 54148
rect 20165 54145 20177 54148
rect 20211 54145 20223 54179
rect 20165 54139 20223 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 20901 54179 20959 54185
rect 20901 54176 20913 54179
rect 20772 54148 20913 54176
rect 20772 54136 20778 54148
rect 20901 54145 20913 54148
rect 20947 54145 20959 54179
rect 20901 54139 20959 54145
rect 21358 54136 21364 54188
rect 21416 54176 21422 54188
rect 22020 54185 22048 54216
rect 23293 54213 23305 54216
rect 23339 54213 23351 54247
rect 23293 54207 23351 54213
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21416 54148 22017 54176
rect 21416 54136 21422 54148
rect 22005 54145 22017 54148
rect 22051 54145 22063 54179
rect 22005 54139 22063 54145
rect 22462 54136 22468 54188
rect 22520 54176 22526 54188
rect 22741 54179 22799 54185
rect 22741 54176 22753 54179
rect 22520 54148 22753 54176
rect 22520 54136 22526 54148
rect 22741 54145 22753 54148
rect 22787 54145 22799 54179
rect 22741 54139 22799 54145
rect 23753 54179 23811 54185
rect 23753 54145 23765 54179
rect 23799 54176 23811 54179
rect 24504 54176 24532 54272
rect 23799 54148 24532 54176
rect 23799 54145 23811 54148
rect 23753 54139 23811 54145
rect 24946 54136 24952 54188
rect 25004 54136 25010 54188
rect 19702 54108 19708 54120
rect 18472 54080 19708 54108
rect 18472 54068 18478 54080
rect 19702 54068 19708 54080
rect 19760 54068 19766 54120
rect 15562 54000 15568 54052
rect 15620 54040 15626 54052
rect 17773 54043 17831 54049
rect 17773 54040 17785 54043
rect 15620 54012 17785 54040
rect 15620 54000 15626 54012
rect 17773 54009 17785 54012
rect 17819 54009 17831 54043
rect 17773 54003 17831 54009
rect 3786 53932 3792 53984
rect 3844 53932 3850 53984
rect 11701 53975 11759 53981
rect 11701 53941 11713 53975
rect 11747 53972 11759 53975
rect 12250 53972 12256 53984
rect 11747 53944 12256 53972
rect 11747 53941 11759 53944
rect 11701 53935 11759 53941
rect 12250 53932 12256 53944
rect 12308 53932 12314 53984
rect 14918 53932 14924 53984
rect 14976 53972 14982 53984
rect 15013 53975 15071 53981
rect 15013 53972 15025 53975
rect 14976 53944 15025 53972
rect 14976 53932 14982 53944
rect 15013 53941 15025 53944
rect 15059 53941 15071 53975
rect 15013 53935 15071 53941
rect 15194 53932 15200 53984
rect 15252 53972 15258 53984
rect 15749 53975 15807 53981
rect 15749 53972 15761 53975
rect 15252 53944 15761 53972
rect 15252 53932 15258 53944
rect 15749 53941 15761 53944
rect 15795 53941 15807 53975
rect 15749 53935 15807 53941
rect 17034 53932 17040 53984
rect 17092 53932 17098 53984
rect 18414 53932 18420 53984
rect 18472 53972 18478 53984
rect 18509 53975 18567 53981
rect 18509 53972 18521 53975
rect 18472 53944 18521 53972
rect 18472 53932 18478 53944
rect 18509 53941 18521 53944
rect 18555 53941 18567 53975
rect 18509 53935 18567 53941
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 19613 53975 19671 53981
rect 19613 53972 19625 53975
rect 19392 53944 19625 53972
rect 19392 53932 19398 53944
rect 19613 53941 19625 53944
rect 19659 53941 19671 53975
rect 19613 53935 19671 53941
rect 20349 53975 20407 53981
rect 20349 53941 20361 53975
rect 20395 53972 20407 53975
rect 20898 53972 20904 53984
rect 20395 53944 20904 53972
rect 20395 53941 20407 53944
rect 20349 53935 20407 53941
rect 20898 53932 20904 53944
rect 20956 53932 20962 53984
rect 21085 53975 21143 53981
rect 21085 53941 21097 53975
rect 21131 53972 21143 53975
rect 21634 53972 21640 53984
rect 21131 53944 21640 53972
rect 21131 53941 21143 53944
rect 21085 53935 21143 53941
rect 21634 53932 21640 53944
rect 21692 53932 21698 53984
rect 22186 53932 22192 53984
rect 22244 53932 22250 53984
rect 22278 53932 22284 53984
rect 22336 53972 22342 53984
rect 22925 53975 22983 53981
rect 22925 53972 22937 53975
rect 22336 53944 22937 53972
rect 22336 53932 22342 53944
rect 22925 53941 22937 53944
rect 22971 53941 22983 53975
rect 22925 53935 22983 53941
rect 23934 53932 23940 53984
rect 23992 53932 23998 53984
rect 25225 53975 25283 53981
rect 25225 53941 25237 53975
rect 25271 53972 25283 53975
rect 25774 53972 25780 53984
rect 25271 53944 25780 53972
rect 25271 53941 25283 53944
rect 25225 53935 25283 53941
rect 25774 53932 25780 53944
rect 25832 53932 25838 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 16393 53771 16451 53777
rect 16393 53737 16405 53771
rect 16439 53768 16451 53771
rect 16574 53768 16580 53780
rect 16439 53740 16580 53768
rect 16439 53737 16451 53740
rect 16393 53731 16451 53737
rect 16574 53728 16580 53740
rect 16632 53728 16638 53780
rect 18874 53728 18880 53780
rect 18932 53728 18938 53780
rect 5534 53660 5540 53712
rect 5592 53660 5598 53712
rect 21269 53703 21327 53709
rect 21269 53669 21281 53703
rect 21315 53700 21327 53703
rect 21542 53700 21548 53712
rect 21315 53672 21548 53700
rect 21315 53669 21327 53672
rect 21269 53663 21327 53669
rect 21542 53660 21548 53672
rect 21600 53660 21606 53712
rect 22370 53660 22376 53712
rect 22428 53700 22434 53712
rect 23109 53703 23167 53709
rect 23109 53700 23121 53703
rect 22428 53672 23121 53700
rect 22428 53660 22434 53672
rect 23109 53669 23121 53672
rect 23155 53669 23167 53703
rect 23109 53663 23167 53669
rect 3237 53635 3295 53641
rect 3237 53601 3249 53635
rect 3283 53632 3295 53635
rect 5552 53632 5580 53660
rect 3283 53604 5580 53632
rect 6549 53635 6607 53641
rect 3283 53601 3295 53604
rect 3237 53595 3295 53601
rect 6549 53601 6561 53635
rect 6595 53632 6607 53635
rect 7374 53632 7380 53644
rect 6595 53604 7380 53632
rect 6595 53601 6607 53604
rect 6549 53595 6607 53601
rect 7374 53592 7380 53604
rect 7432 53592 7438 53644
rect 8389 53635 8447 53641
rect 8389 53601 8401 53635
rect 8435 53632 8447 53635
rect 8846 53632 8852 53644
rect 8435 53604 8852 53632
rect 8435 53601 8447 53604
rect 8389 53595 8447 53601
rect 8846 53592 8852 53604
rect 8904 53592 8910 53644
rect 11054 53592 11060 53644
rect 11112 53592 11118 53644
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 24397 53635 24455 53641
rect 24397 53632 24409 53635
rect 12713 53595 12771 53601
rect 23308 53604 24409 53632
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53564 2283 53567
rect 2271 53536 3924 53564
rect 2271 53533 2283 53536
rect 2225 53527 2283 53533
rect 3896 53496 3924 53536
rect 3970 53524 3976 53576
rect 4028 53524 4034 53576
rect 5534 53524 5540 53576
rect 5592 53524 5598 53576
rect 7285 53567 7343 53573
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 9122 53564 9128 53576
rect 7331 53536 9128 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 9122 53524 9128 53536
rect 9180 53524 9186 53576
rect 10597 53567 10655 53573
rect 10597 53533 10609 53567
rect 10643 53564 10655 53567
rect 12066 53564 12072 53576
rect 10643 53536 12072 53564
rect 10643 53533 10655 53536
rect 10597 53527 10655 53533
rect 12066 53524 12072 53536
rect 12124 53524 12130 53576
rect 12437 53567 12495 53573
rect 12437 53533 12449 53567
rect 12483 53564 12495 53567
rect 12618 53564 12624 53576
rect 12483 53536 12624 53564
rect 12483 53533 12495 53536
rect 12437 53527 12495 53533
rect 12618 53524 12624 53536
rect 12676 53524 12682 53576
rect 13998 53524 14004 53576
rect 14056 53564 14062 53576
rect 14277 53567 14335 53573
rect 14277 53564 14289 53567
rect 14056 53536 14289 53564
rect 14056 53524 14062 53536
rect 14277 53533 14289 53536
rect 14323 53564 14335 53567
rect 14829 53567 14887 53573
rect 14829 53564 14841 53567
rect 14323 53536 14841 53564
rect 14323 53533 14335 53536
rect 14277 53527 14335 53533
rect 14829 53533 14841 53536
rect 14875 53533 14887 53567
rect 14829 53527 14887 53533
rect 15470 53524 15476 53576
rect 15528 53564 15534 53576
rect 15657 53567 15715 53573
rect 15657 53564 15669 53567
rect 15528 53536 15669 53564
rect 15528 53524 15534 53536
rect 15657 53533 15669 53536
rect 15703 53564 15715 53567
rect 16117 53567 16175 53573
rect 16117 53564 16129 53567
rect 15703 53536 16129 53564
rect 15703 53533 15715 53536
rect 15657 53527 15715 53533
rect 16117 53533 16129 53536
rect 16163 53533 16175 53567
rect 16117 53527 16175 53533
rect 16574 53524 16580 53576
rect 16632 53564 16638 53576
rect 16669 53567 16727 53573
rect 16669 53564 16681 53567
rect 16632 53536 16681 53564
rect 16632 53524 16638 53536
rect 16669 53533 16681 53536
rect 16715 53533 16727 53567
rect 16669 53527 16727 53533
rect 17310 53524 17316 53576
rect 17368 53564 17374 53576
rect 17589 53567 17647 53573
rect 17589 53564 17601 53567
rect 17368 53536 17601 53564
rect 17368 53524 17374 53536
rect 17589 53533 17601 53536
rect 17635 53533 17647 53567
rect 17589 53527 17647 53533
rect 18233 53567 18291 53573
rect 18233 53533 18245 53567
rect 18279 53564 18291 53567
rect 18322 53564 18328 53576
rect 18279 53536 18328 53564
rect 18279 53533 18291 53536
rect 18233 53527 18291 53533
rect 18322 53524 18328 53536
rect 18380 53564 18386 53576
rect 18693 53567 18751 53573
rect 18693 53564 18705 53567
rect 18380 53536 18705 53564
rect 18380 53524 18386 53536
rect 18693 53533 18705 53536
rect 18739 53533 18751 53567
rect 18693 53527 18751 53533
rect 19150 53524 19156 53576
rect 19208 53564 19214 53576
rect 19429 53567 19487 53573
rect 19429 53564 19441 53567
rect 19208 53536 19441 53564
rect 19208 53524 19214 53536
rect 19429 53533 19441 53536
rect 19475 53533 19487 53567
rect 19429 53527 19487 53533
rect 19886 53524 19892 53576
rect 19944 53564 19950 53576
rect 20257 53567 20315 53573
rect 20257 53564 20269 53567
rect 19944 53536 20269 53564
rect 19944 53524 19950 53536
rect 20257 53533 20269 53536
rect 20303 53564 20315 53567
rect 20717 53567 20775 53573
rect 20717 53564 20729 53567
rect 20303 53536 20729 53564
rect 20303 53533 20315 53536
rect 20257 53527 20315 53533
rect 20717 53533 20729 53536
rect 20763 53533 20775 53567
rect 20717 53527 20775 53533
rect 20990 53524 20996 53576
rect 21048 53564 21054 53576
rect 21085 53567 21143 53573
rect 21085 53564 21097 53567
rect 21048 53536 21097 53564
rect 21048 53524 21054 53536
rect 21085 53533 21097 53536
rect 21131 53533 21143 53567
rect 21085 53527 21143 53533
rect 21726 53524 21732 53576
rect 21784 53564 21790 53576
rect 22005 53567 22063 53573
rect 22005 53564 22017 53567
rect 21784 53536 22017 53564
rect 21784 53524 21790 53536
rect 22005 53533 22017 53536
rect 22051 53533 22063 53567
rect 22005 53527 22063 53533
rect 22094 53524 22100 53576
rect 22152 53564 22158 53576
rect 22649 53567 22707 53573
rect 22649 53564 22661 53567
rect 22152 53536 22661 53564
rect 22152 53524 22158 53536
rect 22649 53533 22661 53536
rect 22695 53533 22707 53567
rect 22649 53527 22707 53533
rect 22830 53524 22836 53576
rect 22888 53564 22894 53576
rect 23308 53573 23336 53604
rect 24397 53601 24409 53604
rect 24443 53601 24455 53635
rect 24397 53595 24455 53601
rect 23293 53567 23351 53573
rect 23293 53564 23305 53567
rect 22888 53536 23305 53564
rect 22888 53524 22894 53536
rect 23293 53533 23305 53536
rect 23339 53533 23351 53567
rect 23293 53527 23351 53533
rect 23382 53524 23388 53576
rect 23440 53564 23446 53576
rect 23845 53567 23903 53573
rect 23845 53564 23857 53567
rect 23440 53536 23857 53564
rect 23440 53524 23446 53536
rect 23845 53533 23857 53536
rect 23891 53564 23903 53567
rect 24581 53567 24639 53573
rect 24581 53564 24593 53567
rect 23891 53536 24593 53564
rect 23891 53533 23903 53536
rect 23845 53527 23903 53533
rect 24581 53533 24593 53536
rect 24627 53533 24639 53567
rect 24581 53527 24639 53533
rect 24762 53524 24768 53576
rect 24820 53564 24826 53576
rect 25041 53567 25099 53573
rect 25041 53564 25053 53567
rect 24820 53536 25053 53564
rect 24820 53524 24826 53536
rect 25041 53533 25053 53536
rect 25087 53533 25099 53567
rect 25041 53527 25099 53533
rect 7558 53496 7564 53508
rect 3896 53468 7564 53496
rect 7558 53456 7564 53468
rect 7616 53456 7622 53508
rect 15841 53499 15899 53505
rect 15841 53465 15853 53499
rect 15887 53496 15899 53499
rect 16390 53496 16396 53508
rect 15887 53468 16396 53496
rect 15887 53465 15899 53468
rect 15841 53459 15899 53465
rect 16390 53456 16396 53468
rect 16448 53456 16454 53508
rect 18417 53499 18475 53505
rect 18417 53465 18429 53499
rect 18463 53496 18475 53499
rect 18506 53496 18512 53508
rect 18463 53468 18512 53496
rect 18463 53465 18475 53468
rect 18417 53459 18475 53465
rect 18506 53456 18512 53468
rect 18564 53456 18570 53508
rect 20441 53499 20499 53505
rect 20441 53465 20453 53499
rect 20487 53496 20499 53499
rect 20622 53496 20628 53508
rect 20487 53468 20628 53496
rect 20487 53465 20499 53468
rect 20441 53459 20499 53465
rect 20622 53456 20628 53468
rect 20680 53456 20686 53508
rect 24026 53456 24032 53508
rect 24084 53456 24090 53508
rect 4614 53388 4620 53440
rect 4672 53388 4678 53440
rect 14458 53388 14464 53440
rect 14516 53388 14522 53440
rect 16850 53388 16856 53440
rect 16908 53388 16914 53440
rect 17402 53388 17408 53440
rect 17460 53388 17466 53440
rect 19610 53388 19616 53440
rect 19668 53388 19674 53440
rect 21358 53388 21364 53440
rect 21416 53428 21422 53440
rect 21821 53431 21879 53437
rect 21821 53428 21833 53431
rect 21416 53400 21833 53428
rect 21416 53388 21422 53400
rect 21821 53397 21833 53400
rect 21867 53397 21879 53431
rect 21821 53391 21879 53397
rect 22462 53388 22468 53440
rect 22520 53388 22526 53440
rect 25225 53431 25283 53437
rect 25225 53397 25237 53431
rect 25271 53428 25283 53431
rect 25682 53428 25688 53440
rect 25271 53400 25688 53428
rect 25271 53397 25283 53400
rect 25225 53391 25283 53397
rect 25682 53388 25688 53400
rect 25740 53388 25746 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 5166 53184 5172 53236
rect 5224 53224 5230 53236
rect 6178 53224 6184 53236
rect 5224 53196 6184 53224
rect 5224 53184 5230 53196
rect 6178 53184 6184 53196
rect 6236 53184 6242 53236
rect 17310 53184 17316 53236
rect 17368 53184 17374 53236
rect 19150 53184 19156 53236
rect 19208 53224 19214 53236
rect 19521 53227 19579 53233
rect 19521 53224 19533 53227
rect 19208 53196 19533 53224
rect 19208 53184 19214 53196
rect 19521 53193 19533 53196
rect 19567 53193 19579 53227
rect 19521 53187 19579 53193
rect 19702 53184 19708 53236
rect 19760 53184 19766 53236
rect 20990 53184 20996 53236
rect 21048 53184 21054 53236
rect 21726 53184 21732 53236
rect 21784 53224 21790 53236
rect 21821 53227 21879 53233
rect 21821 53224 21833 53227
rect 21784 53196 21833 53224
rect 21784 53184 21790 53196
rect 21821 53193 21833 53196
rect 21867 53193 21879 53227
rect 21821 53187 21879 53193
rect 22094 53184 22100 53236
rect 22152 53224 22158 53236
rect 22281 53227 22339 53233
rect 22281 53224 22293 53227
rect 22152 53196 22293 53224
rect 22152 53184 22158 53196
rect 22281 53193 22293 53196
rect 22327 53193 22339 53227
rect 22281 53187 22339 53193
rect 22554 53184 22560 53236
rect 22612 53184 22618 53236
rect 23017 53227 23075 53233
rect 23017 53193 23029 53227
rect 23063 53224 23075 53227
rect 23290 53224 23296 53236
rect 23063 53196 23296 53224
rect 23063 53193 23075 53196
rect 23017 53187 23075 53193
rect 23290 53184 23296 53196
rect 23348 53184 23354 53236
rect 3973 53159 4031 53165
rect 3973 53125 3985 53159
rect 4019 53156 4031 53159
rect 4430 53156 4436 53168
rect 4019 53128 4436 53156
rect 4019 53125 4031 53128
rect 3973 53119 4031 53125
rect 4430 53116 4436 53128
rect 4488 53116 4494 53168
rect 5813 53159 5871 53165
rect 5813 53125 5825 53159
rect 5859 53156 5871 53159
rect 6270 53156 6276 53168
rect 5859 53128 6276 53156
rect 5859 53125 5871 53128
rect 5813 53119 5871 53125
rect 6270 53116 6276 53128
rect 6328 53116 6334 53168
rect 9125 53159 9183 53165
rect 9125 53125 9137 53159
rect 9171 53156 9183 53159
rect 9214 53156 9220 53168
rect 9171 53128 9220 53156
rect 9171 53125 9183 53128
rect 9125 53119 9183 53125
rect 9214 53116 9220 53128
rect 9272 53116 9278 53168
rect 13630 53116 13636 53168
rect 13688 53156 13694 53168
rect 13817 53159 13875 53165
rect 13817 53156 13829 53159
rect 13688 53128 13829 53156
rect 13688 53116 13694 53128
rect 13817 53125 13829 53128
rect 13863 53125 13875 53159
rect 13817 53119 13875 53125
rect 20714 53116 20720 53168
rect 20772 53156 20778 53168
rect 21177 53159 21235 53165
rect 21177 53156 21189 53159
rect 20772 53128 21189 53156
rect 20772 53116 20778 53128
rect 21177 53125 21189 53128
rect 21223 53125 21235 53159
rect 21177 53119 21235 53125
rect 1670 53048 1676 53100
rect 1728 53048 1734 53100
rect 2961 53091 3019 53097
rect 2961 53057 2973 53091
rect 3007 53088 3019 53091
rect 4154 53088 4160 53100
rect 3007 53060 4160 53088
rect 3007 53057 3019 53060
rect 2961 53051 3019 53057
rect 4154 53048 4160 53060
rect 4212 53048 4218 53100
rect 4706 53048 4712 53100
rect 4764 53048 4770 53100
rect 7282 53048 7288 53100
rect 7340 53088 7346 53100
rect 7929 53091 7987 53097
rect 7929 53088 7941 53091
rect 7340 53060 7941 53088
rect 7340 53048 7346 53060
rect 7929 53057 7941 53060
rect 7975 53057 7987 53091
rect 7929 53051 7987 53057
rect 9306 53048 9312 53100
rect 9364 53088 9370 53100
rect 9769 53091 9827 53097
rect 9769 53088 9781 53091
rect 9364 53060 9781 53088
rect 9364 53048 9370 53060
rect 9769 53057 9781 53060
rect 9815 53057 9827 53091
rect 9769 53051 9827 53057
rect 11882 53048 11888 53100
rect 11940 53048 11946 53100
rect 14366 53048 14372 53100
rect 14424 53088 14430 53100
rect 14645 53091 14703 53097
rect 14645 53088 14657 53091
rect 14424 53060 14657 53088
rect 14424 53048 14430 53060
rect 14645 53057 14657 53060
rect 14691 53088 14703 53091
rect 14921 53091 14979 53097
rect 14921 53088 14933 53091
rect 14691 53060 14933 53088
rect 14691 53057 14703 53060
rect 14645 53051 14703 53057
rect 14921 53057 14933 53060
rect 14967 53057 14979 53091
rect 14921 53051 14979 53057
rect 15838 53048 15844 53100
rect 15896 53088 15902 53100
rect 16117 53091 16175 53097
rect 16117 53088 16129 53091
rect 15896 53060 16129 53088
rect 15896 53048 15902 53060
rect 16117 53057 16129 53060
rect 16163 53088 16175 53091
rect 16393 53091 16451 53097
rect 16393 53088 16405 53091
rect 16163 53060 16405 53088
rect 16163 53057 16175 53060
rect 16117 53051 16175 53057
rect 16393 53057 16405 53060
rect 16439 53057 16451 53091
rect 16393 53051 16451 53057
rect 18782 53048 18788 53100
rect 18840 53088 18846 53100
rect 19061 53091 19119 53097
rect 19061 53088 19073 53091
rect 18840 53060 19073 53088
rect 18840 53048 18846 53060
rect 19061 53057 19073 53060
rect 19107 53088 19119 53091
rect 19337 53091 19395 53097
rect 19337 53088 19349 53091
rect 19107 53060 19349 53088
rect 19107 53057 19119 53060
rect 19061 53051 19119 53057
rect 19337 53057 19349 53060
rect 19383 53057 19395 53091
rect 19337 53051 19395 53057
rect 20254 53048 20260 53100
rect 20312 53088 20318 53100
rect 20533 53091 20591 53097
rect 20533 53088 20545 53091
rect 20312 53060 20545 53088
rect 20312 53048 20318 53060
rect 20533 53057 20545 53060
rect 20579 53088 20591 53091
rect 20809 53091 20867 53097
rect 20809 53088 20821 53091
rect 20579 53060 20821 53088
rect 20579 53057 20591 53060
rect 20533 53051 20591 53057
rect 20809 53057 20821 53060
rect 20855 53057 20867 53091
rect 23308 53088 23336 53184
rect 23477 53091 23535 53097
rect 23477 53088 23489 53091
rect 23308 53060 23489 53088
rect 20809 53051 20867 53057
rect 23477 53057 23489 53060
rect 23523 53057 23535 53091
rect 23477 53051 23535 53057
rect 23566 53048 23572 53100
rect 23624 53088 23630 53100
rect 24121 53091 24179 53097
rect 24121 53088 24133 53091
rect 23624 53060 24133 53088
rect 23624 53048 23630 53060
rect 24121 53057 24133 53060
rect 24167 53088 24179 53091
rect 24397 53091 24455 53097
rect 24397 53088 24409 53091
rect 24167 53060 24409 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 24397 53057 24409 53060
rect 24443 53057 24455 53091
rect 24397 53051 24455 53057
rect 24765 53091 24823 53097
rect 24765 53057 24777 53091
rect 24811 53088 24823 53091
rect 25038 53088 25044 53100
rect 24811 53060 25044 53088
rect 24811 53057 24823 53060
rect 24765 53051 24823 53057
rect 25038 53048 25044 53060
rect 25096 53048 25102 53100
rect 10318 52980 10324 53032
rect 10376 52980 10382 53032
rect 11790 52980 11796 53032
rect 11848 53020 11854 53032
rect 12345 53023 12403 53029
rect 12345 53020 12357 53023
rect 11848 52992 12357 53020
rect 11848 52980 11854 52992
rect 12345 52989 12357 52992
rect 12391 52989 12403 53023
rect 12345 52983 12403 52989
rect 1854 52912 1860 52964
rect 1912 52952 1918 52964
rect 3510 52952 3516 52964
rect 1912 52924 3516 52952
rect 1912 52912 1918 52924
rect 3510 52912 3516 52924
rect 3568 52912 3574 52964
rect 13998 52912 14004 52964
rect 14056 52912 14062 52964
rect 1762 52844 1768 52896
rect 1820 52884 1826 52896
rect 2317 52887 2375 52893
rect 2317 52884 2329 52887
rect 1820 52856 2329 52884
rect 1820 52844 1826 52856
rect 2317 52853 2329 52856
rect 2363 52853 2375 52887
rect 2317 52847 2375 52853
rect 14461 52887 14519 52893
rect 14461 52853 14473 52887
rect 14507 52884 14519 52887
rect 14734 52884 14740 52896
rect 14507 52856 14740 52884
rect 14507 52853 14519 52856
rect 14461 52847 14519 52853
rect 14734 52844 14740 52856
rect 14792 52844 14798 52896
rect 15930 52844 15936 52896
rect 15988 52844 15994 52896
rect 18598 52844 18604 52896
rect 18656 52884 18662 52896
rect 18877 52887 18935 52893
rect 18877 52884 18889 52887
rect 18656 52856 18889 52884
rect 18656 52844 18662 52856
rect 18877 52853 18889 52856
rect 18923 52853 18935 52887
rect 18877 52847 18935 52853
rect 20162 52844 20168 52896
rect 20220 52884 20226 52896
rect 20349 52887 20407 52893
rect 20349 52884 20361 52887
rect 20220 52856 20361 52884
rect 20220 52844 20226 52856
rect 20349 52853 20361 52856
rect 20395 52853 20407 52887
rect 20349 52847 20407 52853
rect 22186 52844 22192 52896
rect 22244 52884 22250 52896
rect 23293 52887 23351 52893
rect 23293 52884 23305 52887
rect 22244 52856 23305 52884
rect 22244 52844 22250 52856
rect 23293 52853 23305 52856
rect 23339 52853 23351 52887
rect 23293 52847 23351 52853
rect 23382 52844 23388 52896
rect 23440 52884 23446 52896
rect 23937 52887 23995 52893
rect 23937 52884 23949 52887
rect 23440 52856 23949 52884
rect 23440 52844 23446 52856
rect 23937 52853 23949 52856
rect 23983 52853 23995 52887
rect 23937 52847 23995 52853
rect 24946 52844 24952 52896
rect 25004 52884 25010 52896
rect 25225 52887 25283 52893
rect 25225 52884 25237 52887
rect 25004 52856 25237 52884
rect 25004 52844 25010 52856
rect 25225 52853 25237 52856
rect 25271 52853 25283 52887
rect 25225 52847 25283 52853
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 2222 52640 2228 52692
rect 2280 52680 2286 52692
rect 3418 52680 3424 52692
rect 2280 52652 3424 52680
rect 2280 52640 2286 52652
rect 3418 52640 3424 52652
rect 3476 52640 3482 52692
rect 12618 52640 12624 52692
rect 12676 52640 12682 52692
rect 13630 52640 13636 52692
rect 13688 52680 13694 52692
rect 14093 52683 14151 52689
rect 14093 52680 14105 52683
rect 13688 52652 14105 52680
rect 13688 52640 13694 52652
rect 14093 52649 14105 52652
rect 14139 52649 14151 52683
rect 14093 52643 14151 52649
rect 24581 52683 24639 52689
rect 24581 52649 24593 52683
rect 24627 52680 24639 52683
rect 24762 52680 24768 52692
rect 24627 52652 24768 52680
rect 24627 52649 24639 52652
rect 24581 52643 24639 52649
rect 24762 52640 24768 52652
rect 24820 52640 24826 52692
rect 1302 52572 1308 52624
rect 1360 52612 1366 52624
rect 3786 52612 3792 52624
rect 1360 52584 3792 52612
rect 1360 52572 1366 52584
rect 3786 52572 3792 52584
rect 3844 52612 3850 52624
rect 25225 52615 25283 52621
rect 3844 52584 4016 52612
rect 3844 52572 3850 52584
rect 3237 52547 3295 52553
rect 3237 52513 3249 52547
rect 3283 52544 3295 52547
rect 3694 52544 3700 52556
rect 3283 52516 3700 52544
rect 3283 52513 3295 52516
rect 3237 52507 3295 52513
rect 3694 52504 3700 52516
rect 3752 52504 3758 52556
rect 3988 52553 4016 52584
rect 25225 52581 25237 52615
rect 25271 52612 25283 52615
rect 25958 52612 25964 52624
rect 25271 52584 25964 52612
rect 25271 52581 25283 52584
rect 25225 52575 25283 52581
rect 25958 52572 25964 52584
rect 26016 52572 26022 52624
rect 3973 52547 4031 52553
rect 3973 52513 3985 52547
rect 4019 52513 4031 52547
rect 3973 52507 4031 52513
rect 4249 52547 4307 52553
rect 4249 52513 4261 52547
rect 4295 52544 4307 52547
rect 4295 52516 7696 52544
rect 4295 52513 4307 52516
rect 4249 52507 4307 52513
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52476 2283 52479
rect 5166 52476 5172 52488
rect 2271 52448 5172 52476
rect 2271 52445 2283 52448
rect 2225 52439 2283 52445
rect 5166 52436 5172 52448
rect 5224 52436 5230 52488
rect 5445 52479 5503 52485
rect 5445 52445 5457 52479
rect 5491 52476 5503 52479
rect 5994 52476 6000 52488
rect 5491 52448 6000 52476
rect 5491 52445 5503 52448
rect 5445 52439 5503 52445
rect 5994 52436 6000 52448
rect 6052 52436 6058 52488
rect 6549 52479 6607 52485
rect 6549 52445 6561 52479
rect 6595 52476 6607 52479
rect 6638 52476 6644 52488
rect 6595 52448 6644 52476
rect 6595 52445 6607 52448
rect 6549 52439 6607 52445
rect 6638 52436 6644 52448
rect 6696 52436 6702 52488
rect 7374 52436 7380 52488
rect 7432 52436 7438 52488
rect 7668 52476 7696 52516
rect 7742 52504 7748 52556
rect 7800 52504 7806 52556
rect 10686 52504 10692 52556
rect 10744 52544 10750 52556
rect 11241 52547 11299 52553
rect 11241 52544 11253 52547
rect 10744 52516 11253 52544
rect 10744 52504 10750 52516
rect 11241 52513 11253 52516
rect 11287 52513 11299 52547
rect 11241 52507 11299 52513
rect 8662 52476 8668 52488
rect 7668 52448 8668 52476
rect 8662 52436 8668 52448
rect 8720 52436 8726 52488
rect 9582 52436 9588 52488
rect 9640 52476 9646 52488
rect 10781 52479 10839 52485
rect 10781 52476 10793 52479
rect 9640 52448 10793 52476
rect 9640 52436 9646 52448
rect 10781 52445 10793 52448
rect 10827 52445 10839 52479
rect 10781 52439 10839 52445
rect 12802 52436 12808 52488
rect 12860 52436 12866 52488
rect 13538 52436 13544 52488
rect 13596 52476 13602 52488
rect 13633 52479 13691 52485
rect 13633 52476 13645 52479
rect 13596 52448 13645 52476
rect 13596 52436 13602 52448
rect 13633 52445 13645 52448
rect 13679 52445 13691 52479
rect 13633 52439 13691 52445
rect 24762 52436 24768 52488
rect 24820 52476 24826 52488
rect 25041 52479 25099 52485
rect 25041 52476 25053 52479
rect 24820 52448 25053 52476
rect 24820 52436 24826 52448
rect 25041 52445 25053 52448
rect 25087 52445 25099 52479
rect 25041 52439 25099 52445
rect 13354 52368 13360 52420
rect 13412 52408 13418 52420
rect 13449 52411 13507 52417
rect 13449 52408 13461 52411
rect 13412 52380 13461 52408
rect 13412 52368 13418 52380
rect 13449 52377 13461 52380
rect 13495 52377 13507 52411
rect 13449 52371 13507 52377
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 1670 52096 1676 52148
rect 1728 52136 1734 52148
rect 2225 52139 2283 52145
rect 2225 52136 2237 52139
rect 1728 52108 2237 52136
rect 1728 52096 1734 52108
rect 2225 52105 2237 52108
rect 2271 52105 2283 52139
rect 2225 52099 2283 52105
rect 4154 52096 4160 52148
rect 4212 52136 4218 52148
rect 7009 52139 7067 52145
rect 7009 52136 7021 52139
rect 4212 52108 7021 52136
rect 4212 52096 4218 52108
rect 7009 52105 7021 52108
rect 7055 52105 7067 52139
rect 7009 52099 7067 52105
rect 11701 52139 11759 52145
rect 11701 52105 11713 52139
rect 11747 52136 11759 52139
rect 11882 52136 11888 52148
rect 11747 52108 11888 52136
rect 11747 52105 11759 52108
rect 11701 52099 11759 52105
rect 11882 52096 11888 52108
rect 11940 52096 11946 52148
rect 12342 52096 12348 52148
rect 12400 52096 12406 52148
rect 13265 52139 13323 52145
rect 13265 52105 13277 52139
rect 13311 52136 13323 52139
rect 13354 52136 13360 52148
rect 13311 52108 13360 52136
rect 13311 52105 13323 52108
rect 13265 52099 13323 52105
rect 13354 52096 13360 52108
rect 13412 52096 13418 52148
rect 25314 52096 25320 52148
rect 25372 52096 25378 52148
rect 4614 52068 4620 52080
rect 1596 52040 4620 52068
rect 1596 52009 1624 52040
rect 4614 52028 4620 52040
rect 4672 52028 4678 52080
rect 6917 52071 6975 52077
rect 6917 52037 6929 52071
rect 6963 52068 6975 52071
rect 9030 52068 9036 52080
rect 6963 52040 9036 52068
rect 6963 52037 6975 52040
rect 6917 52031 6975 52037
rect 9030 52028 9036 52040
rect 9088 52028 9094 52080
rect 1581 52003 1639 52009
rect 1581 51969 1593 52003
rect 1627 51969 1639 52003
rect 1581 51963 1639 51969
rect 2961 52003 3019 52009
rect 2961 51969 2973 52003
rect 3007 51969 3019 52003
rect 2961 51963 3019 51969
rect 4801 52003 4859 52009
rect 4801 51969 4813 52003
rect 4847 52000 4859 52003
rect 7190 52000 7196 52012
rect 4847 51972 7196 52000
rect 4847 51969 4859 51972
rect 4801 51963 4859 51969
rect 2976 51796 3004 51963
rect 7190 51960 7196 51972
rect 7248 51960 7254 52012
rect 8021 52003 8079 52009
rect 8021 51969 8033 52003
rect 8067 51969 8079 52003
rect 8021 51963 8079 51969
rect 3326 51892 3332 51944
rect 3384 51892 3390 51944
rect 4890 51892 4896 51944
rect 4948 51932 4954 51944
rect 5077 51935 5135 51941
rect 5077 51932 5089 51935
rect 4948 51904 5089 51932
rect 4948 51892 4954 51904
rect 5077 51901 5089 51904
rect 5123 51901 5135 51935
rect 5077 51895 5135 51901
rect 8036 51864 8064 51963
rect 9674 51960 9680 52012
rect 9732 51960 9738 52012
rect 10870 51960 10876 52012
rect 10928 52000 10934 52012
rect 11885 52003 11943 52009
rect 11885 52000 11897 52003
rect 10928 51972 11897 52000
rect 10928 51960 10934 51972
rect 11885 51969 11897 51972
rect 11931 51969 11943 52003
rect 11885 51963 11943 51969
rect 11974 51960 11980 52012
rect 12032 52000 12038 52012
rect 12529 52003 12587 52009
rect 12529 52000 12541 52003
rect 12032 51972 12541 52000
rect 12032 51960 12038 51972
rect 12529 51969 12541 51972
rect 12575 51969 12587 52003
rect 12529 51963 12587 51969
rect 8478 51892 8484 51944
rect 8536 51892 8542 51944
rect 9766 51892 9772 51944
rect 9824 51932 9830 51944
rect 10137 51935 10195 51941
rect 10137 51932 10149 51935
rect 9824 51904 10149 51932
rect 9824 51892 9830 51904
rect 10137 51901 10149 51904
rect 10183 51901 10195 51935
rect 10137 51895 10195 51901
rect 10410 51864 10416 51876
rect 8036 51836 10416 51864
rect 10410 51824 10416 51836
rect 10468 51824 10474 51876
rect 4890 51796 4896 51808
rect 2976 51768 4896 51796
rect 4890 51756 4896 51768
rect 4948 51756 4954 51808
rect 25498 51756 25504 51808
rect 25556 51756 25562 51808
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 9950 51552 9956 51604
rect 10008 51592 10014 51604
rect 10229 51595 10287 51601
rect 10229 51592 10241 51595
rect 10008 51564 10241 51592
rect 10008 51552 10014 51564
rect 10229 51561 10241 51564
rect 10275 51561 10287 51595
rect 10229 51555 10287 51561
rect 2866 51416 2872 51468
rect 2924 51416 2930 51468
rect 6914 51456 6920 51468
rect 3896 51428 6920 51456
rect 2225 51391 2283 51397
rect 2225 51357 2237 51391
rect 2271 51388 2283 51391
rect 3896 51388 3924 51428
rect 6914 51416 6920 51428
rect 6972 51416 6978 51468
rect 7006 51416 7012 51468
rect 7064 51456 7070 51468
rect 7561 51459 7619 51465
rect 7561 51456 7573 51459
rect 7064 51428 7573 51456
rect 7064 51416 7070 51428
rect 7561 51425 7573 51428
rect 7607 51425 7619 51459
rect 7561 51419 7619 51425
rect 2271 51360 3924 51388
rect 2271 51357 2283 51360
rect 2225 51351 2283 51357
rect 3970 51348 3976 51400
rect 4028 51348 4034 51400
rect 5445 51391 5503 51397
rect 5445 51357 5457 51391
rect 5491 51388 5503 51391
rect 6730 51388 6736 51400
rect 5491 51360 6736 51388
rect 5491 51357 5503 51360
rect 5445 51351 5503 51357
rect 6730 51348 6736 51360
rect 6788 51348 6794 51400
rect 7098 51348 7104 51400
rect 7156 51348 7162 51400
rect 9214 51348 9220 51400
rect 9272 51388 9278 51400
rect 10413 51391 10471 51397
rect 10413 51388 10425 51391
rect 9272 51360 10425 51388
rect 9272 51348 9278 51360
rect 10413 51357 10425 51360
rect 10459 51357 10471 51391
rect 10413 51351 10471 51357
rect 25041 51391 25099 51397
rect 25041 51357 25053 51391
rect 25087 51388 25099 51391
rect 25498 51388 25504 51400
rect 25087 51360 25504 51388
rect 25087 51357 25099 51360
rect 25041 51351 25099 51357
rect 25498 51348 25504 51360
rect 25556 51348 25562 51400
rect 6178 51280 6184 51332
rect 6236 51280 6242 51332
rect 7006 51280 7012 51332
rect 7064 51320 7070 51332
rect 7190 51320 7196 51332
rect 7064 51292 7196 51320
rect 7064 51280 7070 51292
rect 7190 51280 7196 51292
rect 7248 51280 7254 51332
rect 4246 51212 4252 51264
rect 4304 51252 4310 51264
rect 4617 51255 4675 51261
rect 4617 51252 4629 51255
rect 4304 51224 4629 51252
rect 4304 51212 4310 51224
rect 4617 51221 4629 51224
rect 4663 51221 4675 51255
rect 4617 51215 4675 51221
rect 25222 51212 25228 51264
rect 25280 51212 25286 51264
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 1581 51051 1639 51057
rect 1581 51017 1593 51051
rect 1627 51048 1639 51051
rect 3970 51048 3976 51060
rect 1627 51020 3976 51048
rect 1627 51017 1639 51020
rect 1581 51011 1639 51017
rect 3970 51008 3976 51020
rect 4028 51008 4034 51060
rect 6914 51008 6920 51060
rect 6972 51008 6978 51060
rect 2314 50940 2320 50992
rect 2372 50980 2378 50992
rect 2372 50952 7788 50980
rect 2372 50940 2378 50952
rect 1762 50872 1768 50924
rect 1820 50872 1826 50924
rect 2501 50915 2559 50921
rect 2501 50881 2513 50915
rect 2547 50912 2559 50915
rect 4249 50915 4307 50921
rect 2547 50884 2912 50912
rect 2547 50881 2559 50884
rect 2501 50875 2559 50881
rect 2774 50804 2780 50856
rect 2832 50804 2838 50856
rect 2884 50776 2912 50884
rect 4249 50881 4261 50915
rect 4295 50912 4307 50915
rect 5442 50912 5448 50924
rect 4295 50884 5448 50912
rect 4295 50881 4307 50884
rect 4249 50875 4307 50881
rect 5442 50872 5448 50884
rect 5500 50872 5506 50924
rect 6825 50915 6883 50921
rect 6825 50881 6837 50915
rect 6871 50912 6883 50915
rect 7650 50912 7656 50924
rect 6871 50884 7656 50912
rect 6871 50881 6883 50884
rect 6825 50875 6883 50881
rect 7650 50872 7656 50884
rect 7708 50872 7714 50924
rect 7760 50921 7788 50952
rect 9582 50940 9588 50992
rect 9640 50940 9646 50992
rect 7745 50915 7803 50921
rect 7745 50881 7757 50915
rect 7791 50881 7803 50915
rect 7745 50875 7803 50881
rect 7834 50872 7840 50924
rect 7892 50912 7898 50924
rect 9401 50915 9459 50921
rect 9401 50912 9413 50915
rect 7892 50884 9413 50912
rect 7892 50872 7898 50884
rect 9401 50881 9413 50884
rect 9447 50881 9459 50915
rect 9401 50875 9459 50881
rect 24765 50915 24823 50921
rect 24765 50881 24777 50915
rect 24811 50912 24823 50915
rect 25038 50912 25044 50924
rect 24811 50884 25044 50912
rect 24811 50881 24823 50884
rect 24765 50875 24823 50881
rect 25038 50872 25044 50884
rect 25096 50872 25102 50924
rect 4338 50804 4344 50856
rect 4396 50844 4402 50856
rect 4617 50847 4675 50853
rect 4617 50844 4629 50847
rect 4396 50816 4629 50844
rect 4396 50804 4402 50816
rect 4617 50813 4629 50816
rect 4663 50813 4675 50847
rect 4617 50807 4675 50813
rect 7466 50804 7472 50856
rect 7524 50804 7530 50856
rect 4154 50776 4160 50788
rect 2884 50748 4160 50776
rect 4154 50736 4160 50748
rect 4212 50736 4218 50788
rect 25225 50711 25283 50717
rect 25225 50677 25237 50711
rect 25271 50708 25283 50711
rect 25866 50708 25872 50720
rect 25271 50680 25872 50708
rect 25271 50677 25283 50680
rect 25225 50671 25283 50677
rect 25866 50668 25872 50680
rect 25924 50668 25930 50720
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 6825 50507 6883 50513
rect 6825 50504 6837 50507
rect 5592 50476 6837 50504
rect 5592 50464 5598 50476
rect 6825 50473 6837 50476
rect 6871 50473 6883 50507
rect 6825 50467 6883 50473
rect 9122 50464 9128 50516
rect 9180 50504 9186 50516
rect 9217 50507 9275 50513
rect 9217 50504 9229 50507
rect 9180 50476 9229 50504
rect 9180 50464 9186 50476
rect 9217 50473 9229 50476
rect 9263 50473 9275 50507
rect 9217 50467 9275 50473
rect 2746 50408 4016 50436
rect 1302 50328 1308 50380
rect 1360 50368 1366 50380
rect 2746 50368 2774 50408
rect 1360 50340 2774 50368
rect 3237 50371 3295 50377
rect 1360 50328 1366 50340
rect 3237 50337 3249 50371
rect 3283 50368 3295 50371
rect 3418 50368 3424 50380
rect 3283 50340 3424 50368
rect 3283 50337 3295 50340
rect 3237 50331 3295 50337
rect 3418 50328 3424 50340
rect 3476 50328 3482 50380
rect 3988 50377 4016 50408
rect 3973 50371 4031 50377
rect 3973 50337 3985 50371
rect 4019 50368 4031 50371
rect 5077 50371 5135 50377
rect 5077 50368 5089 50371
rect 4019 50340 5089 50368
rect 4019 50337 4031 50340
rect 3973 50331 4031 50337
rect 5077 50337 5089 50340
rect 5123 50337 5135 50371
rect 5077 50331 5135 50337
rect 2225 50303 2283 50309
rect 2225 50269 2237 50303
rect 2271 50269 2283 50303
rect 2225 50263 2283 50269
rect 4249 50303 4307 50309
rect 4249 50269 4261 50303
rect 4295 50269 4307 50303
rect 4249 50263 4307 50269
rect 2240 50164 2268 50263
rect 4264 50232 4292 50263
rect 5810 50260 5816 50312
rect 5868 50300 5874 50312
rect 7009 50303 7067 50309
rect 7009 50300 7021 50303
rect 5868 50272 7021 50300
rect 5868 50260 5874 50272
rect 7009 50269 7021 50272
rect 7055 50269 7067 50303
rect 7009 50263 7067 50269
rect 9398 50260 9404 50312
rect 9456 50260 9462 50312
rect 8570 50232 8576 50244
rect 4264 50204 8576 50232
rect 8570 50192 8576 50204
rect 8628 50192 8634 50244
rect 5074 50164 5080 50176
rect 2240 50136 5080 50164
rect 5074 50124 5080 50136
rect 5132 50124 5138 50176
rect 25314 50124 25320 50176
rect 25372 50164 25378 50176
rect 25409 50167 25467 50173
rect 25409 50164 25421 50167
rect 25372 50136 25421 50164
rect 25372 50124 25378 50136
rect 25409 50133 25421 50136
rect 25455 50133 25467 50167
rect 25409 50127 25467 50133
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 6549 49963 6607 49969
rect 6549 49960 6561 49963
rect 3988 49932 6561 49960
rect 3145 49895 3203 49901
rect 3145 49861 3157 49895
rect 3191 49892 3203 49895
rect 3510 49892 3516 49904
rect 3191 49864 3516 49892
rect 3191 49861 3203 49864
rect 3145 49855 3203 49861
rect 3510 49852 3516 49864
rect 3568 49852 3574 49904
rect 1946 49784 1952 49836
rect 2004 49784 2010 49836
rect 3988 49833 4016 49932
rect 6549 49929 6561 49932
rect 6595 49960 6607 49963
rect 9858 49960 9864 49972
rect 6595 49932 9864 49960
rect 6595 49929 6607 49932
rect 6549 49923 6607 49929
rect 9858 49920 9864 49932
rect 9916 49920 9922 49972
rect 20806 49920 20812 49972
rect 20864 49960 20870 49972
rect 25133 49963 25191 49969
rect 25133 49960 25145 49963
rect 20864 49932 25145 49960
rect 20864 49920 20870 49932
rect 25133 49929 25145 49932
rect 25179 49929 25191 49963
rect 25133 49923 25191 49929
rect 4246 49852 4252 49904
rect 4304 49852 4310 49904
rect 6365 49895 6423 49901
rect 6365 49892 6377 49895
rect 5474 49864 6377 49892
rect 6365 49861 6377 49864
rect 6411 49892 6423 49895
rect 8938 49892 8944 49904
rect 6411 49864 8944 49892
rect 6411 49861 6423 49864
rect 6365 49855 6423 49861
rect 8938 49852 8944 49864
rect 8996 49852 9002 49904
rect 9306 49852 9312 49904
rect 9364 49852 9370 49904
rect 3973 49827 4031 49833
rect 3973 49793 3985 49827
rect 4019 49793 4031 49827
rect 3973 49787 4031 49793
rect 7742 49784 7748 49836
rect 7800 49824 7806 49836
rect 9125 49827 9183 49833
rect 9125 49824 9137 49827
rect 7800 49796 9137 49824
rect 7800 49784 7806 49796
rect 9125 49793 9137 49796
rect 9171 49793 9183 49827
rect 9125 49787 9183 49793
rect 25314 49784 25320 49836
rect 25372 49784 25378 49836
rect 5997 49759 6055 49765
rect 5997 49725 6009 49759
rect 6043 49756 6055 49759
rect 8846 49756 8852 49768
rect 6043 49728 8852 49756
rect 6043 49725 6055 49728
rect 5997 49719 6055 49725
rect 8846 49716 8852 49728
rect 8904 49716 8910 49768
rect 16022 49716 16028 49768
rect 16080 49756 16086 49768
rect 16850 49756 16856 49768
rect 16080 49728 16856 49756
rect 16080 49716 16086 49728
rect 16850 49716 16856 49728
rect 16908 49716 16914 49768
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 11609 49419 11667 49425
rect 11609 49385 11621 49419
rect 11655 49416 11667 49419
rect 11974 49416 11980 49428
rect 11655 49388 11980 49416
rect 11655 49385 11667 49388
rect 11609 49379 11667 49385
rect 11974 49376 11980 49388
rect 12032 49376 12038 49428
rect 1486 49240 1492 49292
rect 1544 49280 1550 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1544 49252 2053 49280
rect 1544 49240 1550 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49212 1823 49215
rect 1811 49184 2774 49212
rect 1811 49181 1823 49184
rect 1765 49175 1823 49181
rect 2746 49076 2774 49184
rect 10686 49172 10692 49224
rect 10744 49212 10750 49224
rect 11793 49215 11851 49221
rect 11793 49212 11805 49215
rect 10744 49184 11805 49212
rect 10744 49172 10750 49184
rect 11793 49181 11805 49184
rect 11839 49181 11851 49215
rect 11793 49175 11851 49181
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 25314 49212 25320 49224
rect 24903 49184 25320 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 25314 49172 25320 49184
rect 25372 49172 25378 49224
rect 3329 49079 3387 49085
rect 3329 49076 3341 49079
rect 2746 49048 3341 49076
rect 3329 49045 3341 49048
rect 3375 49076 3387 49079
rect 10778 49076 10784 49088
rect 3375 49048 10784 49076
rect 3375 49045 3387 49048
rect 3329 49039 3387 49045
rect 10778 49036 10784 49048
rect 10836 49036 10842 49088
rect 19058 49036 19064 49088
rect 19116 49076 19122 49088
rect 25133 49079 25191 49085
rect 25133 49076 25145 49079
rect 19116 49048 25145 49076
rect 19116 49036 19122 49048
rect 25133 49045 25145 49048
rect 25179 49045 25191 49079
rect 25133 49039 25191 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 12713 48875 12771 48881
rect 12713 48841 12725 48875
rect 12759 48872 12771 48875
rect 12802 48872 12808 48884
rect 12759 48844 12808 48872
rect 12759 48841 12771 48844
rect 12713 48835 12771 48841
rect 12802 48832 12808 48844
rect 12860 48832 12866 48884
rect 12802 48696 12808 48748
rect 12860 48736 12866 48748
rect 12897 48739 12955 48745
rect 12897 48736 12909 48739
rect 12860 48708 12909 48736
rect 12860 48696 12866 48708
rect 12897 48705 12909 48708
rect 12943 48705 12955 48739
rect 12897 48699 12955 48705
rect 25498 48492 25504 48544
rect 25556 48492 25562 48544
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 7282 48084 7288 48136
rect 7340 48124 7346 48136
rect 9950 48124 9956 48136
rect 7340 48096 9956 48124
rect 7340 48084 7346 48096
rect 9950 48084 9956 48096
rect 10008 48084 10014 48136
rect 24857 48127 24915 48133
rect 24857 48093 24869 48127
rect 24903 48124 24915 48127
rect 25314 48124 25320 48136
rect 24903 48096 25320 48124
rect 24903 48093 24915 48096
rect 24857 48087 24915 48093
rect 25314 48084 25320 48096
rect 25372 48084 25378 48136
rect 1302 48016 1308 48068
rect 1360 48056 1366 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 1360 48028 1685 48056
rect 1360 48016 1366 48028
rect 1673 48025 1685 48028
rect 1719 48056 1731 48059
rect 2133 48059 2191 48065
rect 2133 48056 2145 48059
rect 1719 48028 2145 48056
rect 1719 48025 1731 48028
rect 1673 48019 1731 48025
rect 2133 48025 2145 48028
rect 2179 48025 2191 48059
rect 2133 48019 2191 48025
rect 1765 47991 1823 47997
rect 1765 47957 1777 47991
rect 1811 47988 1823 47991
rect 4062 47988 4068 48000
rect 1811 47960 4068 47988
rect 1811 47957 1823 47960
rect 1765 47951 1823 47957
rect 4062 47948 4068 47960
rect 4120 47948 4126 48000
rect 17586 47948 17592 48000
rect 17644 47988 17650 48000
rect 17681 47991 17739 47997
rect 17681 47988 17693 47991
rect 17644 47960 17693 47988
rect 17644 47948 17650 47960
rect 17681 47957 17693 47960
rect 17727 47988 17739 47991
rect 18414 47988 18420 48000
rect 17727 47960 18420 47988
rect 17727 47957 17739 47960
rect 17681 47951 17739 47957
rect 18414 47948 18420 47960
rect 18472 47948 18478 48000
rect 20530 47948 20536 48000
rect 20588 47988 20594 48000
rect 25133 47991 25191 47997
rect 25133 47988 25145 47991
rect 20588 47960 25145 47988
rect 20588 47948 20594 47960
rect 25133 47957 25145 47960
rect 25179 47957 25191 47991
rect 25133 47951 25191 47957
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9030 47744 9036 47796
rect 9088 47784 9094 47796
rect 9125 47787 9183 47793
rect 9125 47784 9137 47787
rect 9088 47756 9137 47784
rect 9088 47744 9094 47756
rect 9125 47753 9137 47756
rect 9171 47753 9183 47787
rect 9125 47747 9183 47753
rect 15930 47744 15936 47796
rect 15988 47784 15994 47796
rect 17221 47787 17279 47793
rect 17221 47784 17233 47787
rect 15988 47756 17233 47784
rect 15988 47744 15994 47756
rect 17221 47753 17233 47756
rect 17267 47753 17279 47787
rect 17221 47747 17279 47753
rect 17402 47744 17408 47796
rect 17460 47784 17466 47796
rect 18417 47787 18475 47793
rect 18417 47784 18429 47787
rect 17460 47756 18429 47784
rect 17460 47744 17466 47756
rect 18417 47753 18429 47756
rect 18463 47753 18475 47787
rect 18417 47747 18475 47753
rect 9309 47651 9367 47657
rect 9309 47617 9321 47651
rect 9355 47648 9367 47651
rect 11790 47648 11796 47660
rect 9355 47620 11796 47648
rect 9355 47617 9367 47620
rect 9309 47611 9367 47617
rect 11790 47608 11796 47620
rect 11848 47608 11854 47660
rect 17313 47651 17371 47657
rect 17313 47617 17325 47651
rect 17359 47648 17371 47651
rect 17586 47648 17592 47660
rect 17359 47620 17592 47648
rect 17359 47617 17371 47620
rect 17313 47611 17371 47617
rect 17586 47608 17592 47620
rect 17644 47608 17650 47660
rect 18506 47608 18512 47660
rect 18564 47648 18570 47660
rect 18690 47648 18696 47660
rect 18564 47620 18696 47648
rect 18564 47608 18570 47620
rect 18690 47608 18696 47620
rect 18748 47648 18754 47660
rect 19061 47651 19119 47657
rect 19061 47648 19073 47651
rect 18748 47620 19073 47648
rect 18748 47608 18754 47620
rect 19061 47617 19073 47620
rect 19107 47617 19119 47651
rect 19061 47611 19119 47617
rect 24489 47651 24547 47657
rect 24489 47617 24501 47651
rect 24535 47648 24547 47651
rect 25498 47648 25504 47660
rect 24535 47620 25504 47648
rect 24535 47617 24547 47620
rect 24489 47611 24547 47617
rect 25498 47608 25504 47620
rect 25556 47608 25562 47660
rect 17405 47583 17463 47589
rect 17405 47549 17417 47583
rect 17451 47549 17463 47583
rect 17405 47543 17463 47549
rect 18601 47583 18659 47589
rect 18601 47549 18613 47583
rect 18647 47549 18659 47583
rect 18601 47543 18659 47549
rect 16298 47472 16304 47524
rect 16356 47512 16362 47524
rect 17420 47512 17448 47543
rect 16356 47484 17448 47512
rect 16356 47472 16362 47484
rect 18414 47472 18420 47524
rect 18472 47512 18478 47524
rect 18616 47512 18644 47543
rect 22738 47540 22744 47592
rect 22796 47580 22802 47592
rect 24765 47583 24823 47589
rect 24765 47580 24777 47583
rect 22796 47552 24777 47580
rect 22796 47540 22802 47552
rect 24765 47549 24777 47552
rect 24811 47549 24823 47583
rect 24765 47543 24823 47549
rect 18472 47484 18644 47512
rect 18472 47472 18478 47484
rect 16574 47404 16580 47456
rect 16632 47444 16638 47456
rect 16853 47447 16911 47453
rect 16853 47444 16865 47447
rect 16632 47416 16865 47444
rect 16632 47404 16638 47416
rect 16853 47413 16865 47416
rect 16899 47413 16911 47447
rect 16853 47407 16911 47413
rect 17494 47404 17500 47456
rect 17552 47444 17558 47456
rect 18049 47447 18107 47453
rect 18049 47444 18061 47447
rect 17552 47416 18061 47444
rect 17552 47404 17558 47416
rect 18049 47413 18061 47416
rect 18095 47413 18107 47447
rect 18049 47407 18107 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9858 47200 9864 47252
rect 9916 47200 9922 47252
rect 15920 47243 15978 47249
rect 15920 47209 15932 47243
rect 15966 47240 15978 47243
rect 18414 47240 18420 47252
rect 15966 47212 18420 47240
rect 15966 47209 15978 47212
rect 15920 47203 15978 47209
rect 18414 47200 18420 47212
rect 18472 47200 18478 47252
rect 21450 47200 21456 47252
rect 21508 47240 21514 47252
rect 21508 47212 22416 47240
rect 21508 47200 21514 47212
rect 9876 47104 9904 47200
rect 18141 47175 18199 47181
rect 18141 47141 18153 47175
rect 18187 47172 18199 47175
rect 18506 47172 18512 47184
rect 18187 47144 18512 47172
rect 18187 47141 18199 47144
rect 18141 47135 18199 47141
rect 18506 47132 18512 47144
rect 18564 47132 18570 47184
rect 10229 47107 10287 47113
rect 10229 47104 10241 47107
rect 9876 47076 10241 47104
rect 10229 47073 10241 47076
rect 10275 47073 10287 47107
rect 10229 47067 10287 47073
rect 15657 47107 15715 47113
rect 15657 47073 15669 47107
rect 15703 47104 15715 47107
rect 16666 47104 16672 47116
rect 15703 47076 16672 47104
rect 15703 47073 15715 47076
rect 15657 47067 15715 47073
rect 16666 47064 16672 47076
rect 16724 47064 16730 47116
rect 17405 47107 17463 47113
rect 17405 47073 17417 47107
rect 17451 47104 17463 47107
rect 17678 47104 17684 47116
rect 17451 47076 17684 47104
rect 17451 47073 17463 47076
rect 17405 47067 17463 47073
rect 17678 47064 17684 47076
rect 17736 47064 17742 47116
rect 18598 47064 18604 47116
rect 18656 47064 18662 47116
rect 18785 47107 18843 47113
rect 18785 47073 18797 47107
rect 18831 47104 18843 47107
rect 19334 47104 19340 47116
rect 18831 47076 19340 47104
rect 18831 47073 18843 47076
rect 18785 47067 18843 47073
rect 19334 47064 19340 47076
rect 19392 47064 19398 47116
rect 22388 47045 22416 47212
rect 25133 47175 25191 47181
rect 25133 47141 25145 47175
rect 25179 47172 25191 47175
rect 25590 47172 25596 47184
rect 25179 47144 25596 47172
rect 25179 47141 25191 47144
rect 25133 47135 25191 47141
rect 25590 47132 25596 47144
rect 25648 47132 25654 47184
rect 22462 47064 22468 47116
rect 22520 47064 22526 47116
rect 22649 47107 22707 47113
rect 22649 47073 22661 47107
rect 22695 47104 22707 47107
rect 22830 47104 22836 47116
rect 22695 47076 22836 47104
rect 22695 47073 22707 47076
rect 22649 47067 22707 47073
rect 22830 47064 22836 47076
rect 22888 47064 22894 47116
rect 22373 47039 22431 47045
rect 22373 47005 22385 47039
rect 22419 47005 22431 47039
rect 25317 47039 25375 47045
rect 25317 47036 25329 47039
rect 22373 46999 22431 47005
rect 24872 47008 25329 47036
rect 8938 46928 8944 46980
rect 8996 46968 9002 46980
rect 8996 46940 9674 46968
rect 8996 46928 9002 46940
rect 9646 46900 9674 46940
rect 10502 46928 10508 46980
rect 10560 46928 10566 46980
rect 12253 46971 12311 46977
rect 12253 46968 12265 46971
rect 10888 46940 10994 46968
rect 11900 46940 12265 46968
rect 10594 46900 10600 46912
rect 9646 46872 10600 46900
rect 10594 46860 10600 46872
rect 10652 46900 10658 46912
rect 10888 46900 10916 46940
rect 11900 46900 11928 46940
rect 12253 46937 12265 46940
rect 12299 46968 12311 46971
rect 12618 46968 12624 46980
rect 12299 46940 12624 46968
rect 12299 46937 12311 46940
rect 12253 46931 12311 46937
rect 12618 46928 12624 46940
rect 12676 46968 12682 46980
rect 14185 46971 14243 46977
rect 14185 46968 14197 46971
rect 12676 46940 14197 46968
rect 12676 46928 12682 46940
rect 14185 46937 14197 46940
rect 14231 46937 14243 46971
rect 14185 46931 14243 46937
rect 16390 46928 16396 46980
rect 16448 46928 16454 46980
rect 18322 46928 18328 46980
rect 18380 46968 18386 46980
rect 18509 46971 18567 46977
rect 18509 46968 18521 46971
rect 18380 46940 18521 46968
rect 18380 46928 18386 46940
rect 18509 46937 18521 46940
rect 18555 46968 18567 46971
rect 19242 46968 19248 46980
rect 18555 46940 19248 46968
rect 18555 46937 18567 46940
rect 18509 46931 18567 46937
rect 19242 46928 19248 46940
rect 19300 46928 19306 46980
rect 21450 46928 21456 46980
rect 21508 46968 21514 46980
rect 21637 46971 21695 46977
rect 21637 46968 21649 46971
rect 21508 46940 21649 46968
rect 21508 46928 21514 46940
rect 21637 46937 21649 46940
rect 21683 46937 21695 46971
rect 21637 46931 21695 46937
rect 24762 46928 24768 46980
rect 24820 46968 24826 46980
rect 24872 46977 24900 47008
rect 25317 47005 25329 47008
rect 25363 47005 25375 47039
rect 25317 46999 25375 47005
rect 24857 46971 24915 46977
rect 24857 46968 24869 46971
rect 24820 46940 24869 46968
rect 24820 46928 24826 46940
rect 24857 46937 24869 46940
rect 24903 46937 24915 46971
rect 24857 46931 24915 46937
rect 10652 46872 11928 46900
rect 11977 46903 12035 46909
rect 10652 46860 10658 46872
rect 11977 46869 11989 46903
rect 12023 46900 12035 46903
rect 12158 46900 12164 46912
rect 12023 46872 12164 46900
rect 12023 46869 12035 46872
rect 11977 46863 12035 46869
rect 12158 46860 12164 46872
rect 12216 46860 12222 46912
rect 17402 46860 17408 46912
rect 17460 46900 17466 46912
rect 17681 46903 17739 46909
rect 17681 46900 17693 46903
rect 17460 46872 17693 46900
rect 17460 46860 17466 46872
rect 17681 46869 17693 46872
rect 17727 46869 17739 46903
rect 17681 46863 17739 46869
rect 22002 46860 22008 46912
rect 22060 46860 22066 46912
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 7193 46699 7251 46705
rect 7193 46665 7205 46699
rect 7239 46696 7251 46699
rect 7466 46696 7472 46708
rect 7239 46668 7472 46696
rect 7239 46665 7251 46668
rect 7193 46659 7251 46665
rect 7466 46656 7472 46668
rect 7524 46656 7530 46708
rect 10870 46656 10876 46708
rect 10928 46656 10934 46708
rect 14458 46696 14464 46708
rect 12636 46668 14464 46696
rect 12636 46637 12664 46668
rect 14458 46656 14464 46668
rect 14516 46656 14522 46708
rect 18414 46656 18420 46708
rect 18472 46696 18478 46708
rect 18601 46699 18659 46705
rect 18601 46696 18613 46699
rect 18472 46668 18613 46696
rect 18472 46656 18478 46668
rect 18601 46665 18613 46668
rect 18647 46665 18659 46699
rect 18601 46659 18659 46665
rect 18966 46656 18972 46708
rect 19024 46696 19030 46708
rect 20809 46699 20867 46705
rect 20809 46696 20821 46699
rect 19024 46668 20821 46696
rect 19024 46656 19030 46668
rect 20809 46665 20821 46668
rect 20855 46665 20867 46699
rect 20809 46659 20867 46665
rect 21910 46656 21916 46708
rect 21968 46696 21974 46708
rect 22094 46696 22100 46708
rect 21968 46668 22100 46696
rect 21968 46656 21974 46668
rect 22094 46656 22100 46668
rect 22152 46696 22158 46708
rect 22649 46699 22707 46705
rect 22649 46696 22661 46699
rect 22152 46668 22661 46696
rect 22152 46656 22158 46668
rect 22649 46665 22661 46668
rect 22695 46665 22707 46699
rect 22649 46659 22707 46665
rect 22741 46699 22799 46705
rect 22741 46665 22753 46699
rect 22787 46696 22799 46699
rect 23382 46696 23388 46708
rect 22787 46668 23388 46696
rect 22787 46665 22799 46668
rect 22741 46659 22799 46665
rect 23382 46656 23388 46668
rect 23440 46656 23446 46708
rect 12621 46631 12679 46637
rect 12621 46597 12633 46631
rect 12667 46597 12679 46631
rect 12621 46591 12679 46597
rect 12710 46588 12716 46640
rect 12768 46628 12774 46640
rect 12768 46600 13110 46628
rect 12768 46588 12774 46600
rect 15102 46588 15108 46640
rect 15160 46628 15166 46640
rect 15160 46600 15318 46628
rect 15160 46588 15166 46600
rect 16390 46588 16396 46640
rect 16448 46628 16454 46640
rect 17402 46628 17408 46640
rect 16448 46600 17408 46628
rect 16448 46588 16454 46600
rect 17402 46588 17408 46600
rect 17460 46628 17466 46640
rect 17460 46600 17618 46628
rect 17460 46588 17466 46600
rect 19242 46588 19248 46640
rect 19300 46628 19306 46640
rect 19300 46600 19826 46628
rect 19300 46588 19306 46600
rect 7377 46563 7435 46569
rect 7377 46529 7389 46563
rect 7423 46560 7435 46563
rect 9582 46560 9588 46572
rect 7423 46532 9588 46560
rect 7423 46529 7435 46532
rect 7377 46523 7435 46529
rect 9582 46520 9588 46532
rect 9640 46520 9646 46572
rect 11054 46520 11060 46572
rect 11112 46520 11118 46572
rect 12345 46495 12403 46501
rect 12345 46461 12357 46495
rect 12391 46461 12403 46495
rect 14553 46495 14611 46501
rect 14553 46492 14565 46495
rect 12345 46455 12403 46461
rect 13648 46464 14565 46492
rect 11882 46316 11888 46368
rect 11940 46356 11946 46368
rect 12360 46356 12388 46455
rect 12710 46356 12716 46368
rect 11940 46328 12716 46356
rect 11940 46316 11946 46328
rect 12710 46316 12716 46328
rect 12768 46356 12774 46368
rect 13648 46356 13676 46464
rect 14553 46461 14565 46464
rect 14599 46461 14611 46495
rect 14553 46455 14611 46461
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 14875 46464 16712 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 16684 46368 16712 46464
rect 16758 46452 16764 46504
rect 16816 46492 16822 46504
rect 16853 46495 16911 46501
rect 16853 46492 16865 46495
rect 16816 46464 16865 46492
rect 16816 46452 16822 46464
rect 16853 46461 16865 46464
rect 16899 46461 16911 46495
rect 16853 46455 16911 46461
rect 17129 46495 17187 46501
rect 17129 46461 17141 46495
rect 17175 46492 17187 46495
rect 18598 46492 18604 46504
rect 17175 46464 18604 46492
rect 17175 46461 17187 46464
rect 17129 46455 17187 46461
rect 18598 46452 18604 46464
rect 18656 46452 18662 46504
rect 19061 46495 19119 46501
rect 19061 46461 19073 46495
rect 19107 46461 19119 46495
rect 19061 46455 19119 46461
rect 12768 46328 13676 46356
rect 12768 46316 12774 46328
rect 13722 46316 13728 46368
rect 13780 46356 13786 46368
rect 14093 46359 14151 46365
rect 14093 46356 14105 46359
rect 13780 46328 14105 46356
rect 13780 46316 13786 46328
rect 14093 46325 14105 46328
rect 14139 46325 14151 46359
rect 14093 46319 14151 46325
rect 16298 46316 16304 46368
rect 16356 46316 16362 46368
rect 16666 46316 16672 46368
rect 16724 46316 16730 46368
rect 19076 46356 19104 46455
rect 19334 46452 19340 46504
rect 19392 46452 19398 46504
rect 22462 46452 22468 46504
rect 22520 46492 22526 46504
rect 22833 46495 22891 46501
rect 22833 46492 22845 46495
rect 22520 46464 22845 46492
rect 22520 46452 22526 46464
rect 22833 46461 22845 46464
rect 22879 46492 22891 46495
rect 23293 46495 23351 46501
rect 23293 46492 23305 46495
rect 22879 46464 23305 46492
rect 22879 46461 22891 46464
rect 22833 46455 22891 46461
rect 23293 46461 23305 46464
rect 23339 46461 23351 46495
rect 23293 46455 23351 46461
rect 24486 46452 24492 46504
rect 24544 46452 24550 46504
rect 24578 46452 24584 46504
rect 24636 46492 24642 46504
rect 24765 46495 24823 46501
rect 24765 46492 24777 46495
rect 24636 46464 24777 46492
rect 24636 46452 24642 46464
rect 24765 46461 24777 46464
rect 24811 46461 24823 46495
rect 24765 46455 24823 46461
rect 19518 46356 19524 46368
rect 19076 46328 19524 46356
rect 19518 46316 19524 46328
rect 19576 46316 19582 46368
rect 21082 46316 21088 46368
rect 21140 46316 21146 46368
rect 21910 46316 21916 46368
rect 21968 46316 21974 46368
rect 22281 46359 22339 46365
rect 22281 46325 22293 46359
rect 22327 46356 22339 46359
rect 22646 46356 22652 46368
rect 22327 46328 22652 46356
rect 22327 46325 22339 46328
rect 22281 46319 22339 46325
rect 22646 46316 22652 46328
rect 22704 46316 22710 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 5994 46112 6000 46164
rect 6052 46152 6058 46164
rect 8113 46155 8171 46161
rect 8113 46152 8125 46155
rect 6052 46124 8125 46152
rect 6052 46112 6058 46124
rect 8113 46121 8125 46124
rect 8159 46121 8171 46155
rect 8113 46115 8171 46121
rect 9125 46155 9183 46161
rect 9125 46121 9137 46155
rect 9171 46152 9183 46155
rect 9214 46152 9220 46164
rect 9171 46124 9220 46152
rect 9171 46121 9183 46124
rect 9125 46115 9183 46121
rect 9214 46112 9220 46124
rect 9272 46112 9278 46164
rect 10686 46112 10692 46164
rect 10744 46112 10750 46164
rect 17402 46112 17408 46164
rect 17460 46152 17466 46164
rect 18693 46155 18751 46161
rect 18693 46152 18705 46155
rect 17460 46124 18705 46152
rect 17460 46112 17466 46124
rect 18693 46121 18705 46124
rect 18739 46152 18751 46155
rect 19150 46152 19156 46164
rect 18739 46124 19156 46152
rect 18739 46121 18751 46124
rect 18693 46115 18751 46121
rect 19150 46112 19156 46124
rect 19208 46112 19214 46164
rect 24486 46112 24492 46164
rect 24544 46152 24550 46164
rect 25409 46155 25467 46161
rect 25409 46152 25421 46155
rect 24544 46124 25421 46152
rect 24544 46112 24550 46124
rect 25409 46121 25421 46124
rect 25455 46152 25467 46155
rect 25498 46152 25504 46164
rect 25455 46124 25504 46152
rect 25455 46121 25467 46124
rect 25409 46115 25467 46121
rect 25498 46112 25504 46124
rect 25556 46112 25562 46164
rect 7650 46044 7656 46096
rect 7708 46084 7714 46096
rect 10045 46087 10103 46093
rect 10045 46084 10057 46087
rect 7708 46056 10057 46084
rect 7708 46044 7714 46056
rect 10045 46053 10057 46056
rect 10091 46053 10103 46087
rect 10045 46047 10103 46053
rect 11348 46056 12020 46084
rect 1857 46019 1915 46025
rect 1857 45985 1869 46019
rect 1903 46016 1915 46019
rect 9122 46016 9128 46028
rect 1903 45988 9128 46016
rect 1903 45985 1915 45988
rect 1857 45979 1915 45985
rect 9122 45976 9128 45988
rect 9180 45976 9186 46028
rect 11348 46025 11376 46056
rect 11333 46019 11391 46025
rect 11333 45985 11345 46019
rect 11379 45985 11391 46019
rect 11333 45979 11391 45985
rect 11882 45976 11888 46028
rect 11940 45976 11946 46028
rect 11992 46016 12020 46056
rect 12158 46016 12164 46028
rect 11992 45988 12164 46016
rect 12158 45976 12164 45988
rect 12216 45976 12222 46028
rect 12618 45976 12624 46028
rect 12676 46016 12682 46028
rect 14090 46016 14096 46028
rect 12676 45988 14096 46016
rect 12676 45976 12682 45988
rect 14090 45976 14096 45988
rect 14148 45976 14154 46028
rect 20162 45976 20168 46028
rect 20220 45976 20226 46028
rect 20349 46019 20407 46025
rect 20349 45985 20361 46019
rect 20395 46016 20407 46019
rect 20438 46016 20444 46028
rect 20395 45988 20444 46016
rect 20395 45985 20407 45988
rect 20349 45979 20407 45985
rect 20438 45976 20444 45988
rect 20496 45976 20502 46028
rect 21358 45976 21364 46028
rect 21416 45976 21422 46028
rect 21450 45976 21456 46028
rect 21508 45976 21514 46028
rect 1302 45908 1308 45960
rect 1360 45948 1366 45960
rect 1581 45951 1639 45957
rect 1581 45948 1593 45951
rect 1360 45920 1593 45948
rect 1360 45908 1366 45920
rect 1581 45917 1593 45920
rect 1627 45917 1639 45951
rect 1581 45911 1639 45917
rect 7466 45908 7472 45960
rect 7524 45948 7530 45960
rect 9309 45951 9367 45957
rect 9309 45948 9321 45951
rect 7524 45920 9321 45948
rect 7524 45908 7530 45920
rect 9309 45917 9321 45920
rect 9355 45917 9367 45951
rect 9309 45911 9367 45917
rect 10042 45908 10048 45960
rect 10100 45948 10106 45960
rect 10229 45951 10287 45957
rect 10229 45948 10241 45951
rect 10100 45920 10241 45948
rect 10100 45908 10106 45920
rect 10229 45917 10241 45920
rect 10275 45917 10287 45951
rect 10229 45911 10287 45917
rect 23201 45951 23259 45957
rect 23201 45917 23213 45951
rect 23247 45917 23259 45951
rect 23201 45911 23259 45917
rect 23477 45951 23535 45957
rect 23477 45917 23489 45951
rect 23523 45948 23535 45951
rect 23658 45948 23664 45960
rect 23523 45920 23664 45948
rect 23523 45917 23535 45920
rect 23477 45911 23535 45917
rect 6914 45840 6920 45892
rect 6972 45880 6978 45892
rect 8021 45883 8079 45889
rect 8021 45880 8033 45883
rect 6972 45852 8033 45880
rect 6972 45840 6978 45852
rect 8021 45849 8033 45852
rect 8067 45880 8079 45883
rect 8481 45883 8539 45889
rect 8481 45880 8493 45883
rect 8067 45852 8493 45880
rect 8067 45849 8079 45852
rect 8021 45843 8079 45849
rect 8481 45849 8493 45852
rect 8527 45849 8539 45883
rect 8481 45843 8539 45849
rect 11057 45883 11115 45889
rect 11057 45849 11069 45883
rect 11103 45880 11115 45883
rect 11698 45880 11704 45892
rect 11103 45852 11704 45880
rect 11103 45849 11115 45852
rect 11057 45843 11115 45849
rect 11698 45840 11704 45852
rect 11756 45840 11762 45892
rect 12618 45840 12624 45892
rect 12676 45840 12682 45892
rect 19429 45883 19487 45889
rect 19429 45849 19441 45883
rect 19475 45880 19487 45883
rect 19610 45880 19616 45892
rect 19475 45852 19616 45880
rect 19475 45849 19487 45852
rect 19429 45843 19487 45849
rect 19610 45840 19616 45852
rect 19668 45880 19674 45892
rect 19668 45852 20116 45880
rect 19668 45840 19674 45852
rect 20088 45824 20116 45852
rect 11146 45772 11152 45824
rect 11204 45772 11210 45824
rect 13446 45772 13452 45824
rect 13504 45812 13510 45824
rect 13633 45815 13691 45821
rect 13633 45812 13645 45815
rect 13504 45784 13645 45812
rect 13504 45772 13510 45784
rect 13633 45781 13645 45784
rect 13679 45781 13691 45815
rect 13633 45775 13691 45781
rect 16390 45772 16396 45824
rect 16448 45772 16454 45824
rect 19705 45815 19763 45821
rect 19705 45781 19717 45815
rect 19751 45812 19763 45815
rect 19886 45812 19892 45824
rect 19751 45784 19892 45812
rect 19751 45781 19763 45784
rect 19705 45775 19763 45781
rect 19886 45772 19892 45784
rect 19944 45772 19950 45824
rect 20070 45772 20076 45824
rect 20128 45772 20134 45824
rect 20901 45815 20959 45821
rect 20901 45781 20913 45815
rect 20947 45812 20959 45815
rect 20990 45812 20996 45824
rect 20947 45784 20996 45812
rect 20947 45781 20959 45784
rect 20901 45775 20959 45781
rect 20990 45772 20996 45784
rect 21048 45772 21054 45824
rect 21266 45772 21272 45824
rect 21324 45772 21330 45824
rect 23216 45812 23244 45911
rect 23658 45908 23664 45920
rect 23716 45908 23722 45960
rect 24489 45815 24547 45821
rect 24489 45812 24501 45815
rect 23216 45784 24501 45812
rect 24489 45781 24501 45784
rect 24535 45812 24547 45815
rect 24854 45812 24860 45824
rect 24535 45784 24860 45812
rect 24535 45781 24547 45784
rect 24489 45775 24547 45781
rect 24854 45772 24860 45784
rect 24912 45772 24918 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 1302 45568 1308 45620
rect 1360 45608 1366 45620
rect 1397 45611 1455 45617
rect 1397 45608 1409 45611
rect 1360 45580 1409 45608
rect 1360 45568 1366 45580
rect 1397 45577 1409 45580
rect 1443 45577 1455 45611
rect 16390 45608 16396 45620
rect 1397 45571 1455 45577
rect 15028 45580 16396 45608
rect 8846 45500 8852 45552
rect 8904 45500 8910 45552
rect 9766 45540 9772 45552
rect 9232 45512 9772 45540
rect 8864 45404 8892 45500
rect 9232 45484 9260 45512
rect 9766 45500 9772 45512
rect 9824 45500 9830 45552
rect 14090 45500 14096 45552
rect 14148 45540 14154 45552
rect 15028 45540 15056 45580
rect 16390 45568 16396 45580
rect 16448 45568 16454 45620
rect 19334 45568 19340 45620
rect 19392 45608 19398 45620
rect 20165 45611 20223 45617
rect 20165 45608 20177 45611
rect 19392 45580 20177 45608
rect 19392 45568 19398 45580
rect 20165 45577 20177 45580
rect 20211 45577 20223 45611
rect 23753 45611 23811 45617
rect 23753 45608 23765 45611
rect 20165 45571 20223 45577
rect 22664 45580 23765 45608
rect 15102 45540 15108 45552
rect 14148 45512 15108 45540
rect 14148 45500 14154 45512
rect 15102 45500 15108 45512
rect 15160 45500 15166 45552
rect 19150 45500 19156 45552
rect 19208 45500 19214 45552
rect 21450 45500 21456 45552
rect 21508 45540 21514 45552
rect 22664 45540 22692 45580
rect 23753 45577 23765 45580
rect 23799 45577 23811 45611
rect 23753 45571 23811 45577
rect 21508 45512 22692 45540
rect 21508 45500 21514 45512
rect 9214 45432 9220 45484
rect 9272 45432 9278 45484
rect 10594 45432 10600 45484
rect 10652 45472 10658 45484
rect 11241 45475 11299 45481
rect 11241 45472 11253 45475
rect 10652 45444 11253 45472
rect 10652 45432 10658 45444
rect 11241 45441 11253 45444
rect 11287 45441 11299 45475
rect 23566 45472 23572 45484
rect 23414 45444 23572 45472
rect 11241 45435 11299 45441
rect 23566 45432 23572 45444
rect 23624 45472 23630 45484
rect 24029 45475 24087 45481
rect 24029 45472 24041 45475
rect 23624 45444 24041 45472
rect 23624 45432 23630 45444
rect 24029 45441 24041 45444
rect 24075 45441 24087 45475
rect 24029 45435 24087 45441
rect 24118 45432 24124 45484
rect 24176 45472 24182 45484
rect 24765 45475 24823 45481
rect 24765 45472 24777 45475
rect 24176 45444 24777 45472
rect 24176 45432 24182 45444
rect 24765 45441 24777 45444
rect 24811 45441 24823 45475
rect 24765 45435 24823 45441
rect 9493 45407 9551 45413
rect 9493 45404 9505 45407
rect 8864 45376 9505 45404
rect 9493 45373 9505 45376
rect 9539 45373 9551 45407
rect 9493 45367 9551 45373
rect 9858 45364 9864 45416
rect 9916 45404 9922 45416
rect 11517 45407 11575 45413
rect 11517 45404 11529 45407
rect 9916 45376 11529 45404
rect 9916 45364 9922 45376
rect 11517 45373 11529 45376
rect 11563 45373 11575 45407
rect 11517 45367 11575 45373
rect 12158 45364 12164 45416
rect 12216 45364 12222 45416
rect 14366 45364 14372 45416
rect 14424 45364 14430 45416
rect 14645 45407 14703 45413
rect 14645 45373 14657 45407
rect 14691 45404 14703 45407
rect 16298 45404 16304 45416
rect 14691 45376 16304 45404
rect 14691 45373 14703 45376
rect 14645 45367 14703 45373
rect 16298 45364 16304 45376
rect 16356 45364 16362 45416
rect 18322 45364 18328 45416
rect 18380 45404 18386 45416
rect 18417 45407 18475 45413
rect 18417 45404 18429 45407
rect 18380 45376 18429 45404
rect 18380 45364 18386 45376
rect 18417 45373 18429 45376
rect 18463 45373 18475 45407
rect 18417 45367 18475 45373
rect 18693 45407 18751 45413
rect 18693 45373 18705 45407
rect 18739 45404 18751 45407
rect 20070 45404 20076 45416
rect 18739 45376 20076 45404
rect 18739 45373 18751 45376
rect 18693 45367 18751 45373
rect 20070 45364 20076 45376
rect 20128 45364 20134 45416
rect 20254 45364 20260 45416
rect 20312 45404 20318 45416
rect 20441 45407 20499 45413
rect 20441 45404 20453 45407
rect 20312 45376 20453 45404
rect 20312 45364 20318 45376
rect 20441 45373 20453 45376
rect 20487 45404 20499 45407
rect 21082 45404 21088 45416
rect 20487 45376 21088 45404
rect 20487 45373 20499 45376
rect 20441 45367 20499 45373
rect 21082 45364 21088 45376
rect 21140 45364 21146 45416
rect 22005 45407 22063 45413
rect 22005 45373 22017 45407
rect 22051 45373 22063 45407
rect 22005 45367 22063 45373
rect 22281 45407 22339 45413
rect 22281 45373 22293 45407
rect 22327 45404 22339 45407
rect 22327 45376 23428 45404
rect 22327 45373 22339 45376
rect 22281 45367 22339 45373
rect 10502 45296 10508 45348
rect 10560 45336 10566 45348
rect 10965 45339 11023 45345
rect 10965 45336 10977 45339
rect 10560 45308 10977 45336
rect 10560 45296 10566 45308
rect 10965 45305 10977 45308
rect 11011 45336 11023 45339
rect 12176 45336 12204 45364
rect 20717 45339 20775 45345
rect 20717 45336 20729 45339
rect 11011 45308 12204 45336
rect 20364 45308 20729 45336
rect 11011 45305 11023 45308
rect 10965 45299 11023 45305
rect 12161 45271 12219 45277
rect 12161 45237 12173 45271
rect 12207 45268 12219 45271
rect 12342 45268 12348 45280
rect 12207 45240 12348 45268
rect 12207 45237 12219 45240
rect 12161 45231 12219 45237
rect 12342 45228 12348 45240
rect 12400 45228 12406 45280
rect 16114 45228 16120 45280
rect 16172 45228 16178 45280
rect 18874 45228 18880 45280
rect 18932 45268 18938 45280
rect 20364 45268 20392 45308
rect 20717 45305 20729 45308
rect 20763 45336 20775 45339
rect 20898 45336 20904 45348
rect 20763 45308 20904 45336
rect 20763 45305 20775 45308
rect 20717 45299 20775 45305
rect 20898 45296 20904 45308
rect 20956 45336 20962 45348
rect 21266 45336 21272 45348
rect 20956 45308 21272 45336
rect 20956 45296 20962 45308
rect 21266 45296 21272 45308
rect 21324 45296 21330 45348
rect 18932 45240 20392 45268
rect 22020 45268 22048 45367
rect 23400 45348 23428 45376
rect 24486 45364 24492 45416
rect 24544 45364 24550 45416
rect 23382 45296 23388 45348
rect 23440 45296 23446 45348
rect 22278 45268 22284 45280
rect 22020 45240 22284 45268
rect 18932 45228 18938 45240
rect 22278 45228 22284 45240
rect 22336 45228 22342 45280
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 7374 45024 7380 45076
rect 7432 45064 7438 45076
rect 9309 45067 9367 45073
rect 9309 45064 9321 45067
rect 7432 45036 9321 45064
rect 7432 45024 7438 45036
rect 9309 45033 9321 45036
rect 9355 45033 9367 45067
rect 9309 45027 9367 45033
rect 11238 45024 11244 45076
rect 11296 45064 11302 45076
rect 11609 45067 11667 45073
rect 11609 45064 11621 45067
rect 11296 45036 11621 45064
rect 11296 45024 11302 45036
rect 11609 45033 11621 45036
rect 11655 45033 11667 45067
rect 11609 45027 11667 45033
rect 12066 45024 12072 45076
rect 12124 45064 12130 45076
rect 12437 45067 12495 45073
rect 12437 45064 12449 45067
rect 12124 45036 12449 45064
rect 12124 45024 12130 45036
rect 12437 45033 12449 45036
rect 12483 45033 12495 45067
rect 12437 45027 12495 45033
rect 12802 45024 12808 45076
rect 12860 45064 12866 45076
rect 12989 45067 13047 45073
rect 12989 45064 13001 45067
rect 12860 45036 13001 45064
rect 12860 45024 12866 45036
rect 12989 45033 13001 45036
rect 13035 45033 13047 45067
rect 12989 45027 13047 45033
rect 15368 45067 15426 45073
rect 15368 45033 15380 45067
rect 15414 45064 15426 45067
rect 15414 45036 16528 45064
rect 15414 45033 15426 45036
rect 15368 45027 15426 45033
rect 4706 44956 4712 45008
rect 4764 44996 4770 45008
rect 7929 44999 7987 45005
rect 7929 44996 7941 44999
rect 4764 44968 7941 44996
rect 4764 44956 4770 44968
rect 7929 44965 7941 44968
rect 7975 44965 7987 44999
rect 7929 44959 7987 44965
rect 14366 44956 14372 45008
rect 14424 44996 14430 45008
rect 16500 44996 16528 45036
rect 16666 45024 16672 45076
rect 16724 45064 16730 45076
rect 16853 45067 16911 45073
rect 16853 45064 16865 45067
rect 16724 45036 16865 45064
rect 16724 45024 16730 45036
rect 16853 45033 16865 45036
rect 16899 45064 16911 45067
rect 16942 45064 16948 45076
rect 16899 45036 16948 45064
rect 16899 45033 16911 45036
rect 16853 45027 16911 45033
rect 16942 45024 16948 45036
rect 17000 45024 17006 45076
rect 17678 44996 17684 45008
rect 14424 44968 15148 44996
rect 16500 44968 17684 44996
rect 14424 44956 14430 44968
rect 12618 44888 12624 44940
rect 12676 44928 12682 44940
rect 13541 44931 13599 44937
rect 13541 44928 13553 44931
rect 12676 44900 13553 44928
rect 12676 44888 12682 44900
rect 13541 44897 13553 44900
rect 13587 44928 13599 44931
rect 13722 44928 13728 44940
rect 13587 44900 13728 44928
rect 13587 44897 13599 44900
rect 13541 44891 13599 44897
rect 13722 44888 13728 44900
rect 13780 44888 13786 44940
rect 15120 44937 15148 44968
rect 17678 44956 17684 44968
rect 17736 44956 17742 45008
rect 15105 44931 15163 44937
rect 15105 44897 15117 44931
rect 15151 44928 15163 44931
rect 16758 44928 16764 44940
rect 15151 44900 16764 44928
rect 15151 44897 15163 44900
rect 15105 44891 15163 44897
rect 16758 44888 16764 44900
rect 16816 44888 16822 44940
rect 23014 44888 23020 44940
rect 23072 44928 23078 44940
rect 23566 44928 23572 44940
rect 23072 44900 23572 44928
rect 23072 44888 23078 44900
rect 23566 44888 23572 44900
rect 23624 44928 23630 44940
rect 24397 44931 24455 44937
rect 24397 44928 24409 44931
rect 23624 44900 24409 44928
rect 23624 44888 23630 44900
rect 24397 44897 24409 44900
rect 24443 44897 24455 44931
rect 24397 44891 24455 44897
rect 12342 44820 12348 44872
rect 12400 44860 12406 44872
rect 14366 44860 14372 44872
rect 12400 44832 14372 44860
rect 12400 44820 12406 44832
rect 14366 44820 14372 44832
rect 14424 44820 14430 44872
rect 19518 44820 19524 44872
rect 19576 44820 19582 44872
rect 21082 44820 21088 44872
rect 21140 44860 21146 44872
rect 21545 44863 21603 44869
rect 21545 44860 21557 44863
rect 21140 44832 21557 44860
rect 21140 44820 21146 44832
rect 21545 44829 21557 44832
rect 21591 44860 21603 44863
rect 21591 44832 22094 44860
rect 21591 44829 21603 44832
rect 21545 44823 21603 44829
rect 7745 44795 7803 44801
rect 7745 44761 7757 44795
rect 7791 44792 7803 44795
rect 9217 44795 9275 44801
rect 7791 44764 8340 44792
rect 7791 44761 7803 44764
rect 7745 44755 7803 44761
rect 6457 44727 6515 44733
rect 6457 44693 6469 44727
rect 6503 44724 6515 44727
rect 6638 44724 6644 44736
rect 6503 44696 6644 44724
rect 6503 44693 6515 44696
rect 6457 44687 6515 44693
rect 6638 44684 6644 44696
rect 6696 44684 6702 44736
rect 7098 44684 7104 44736
rect 7156 44684 7162 44736
rect 8312 44733 8340 44764
rect 9217 44761 9229 44795
rect 9263 44792 9275 44795
rect 11149 44795 11207 44801
rect 9263 44764 9812 44792
rect 9263 44761 9275 44764
rect 9217 44755 9275 44761
rect 9784 44736 9812 44764
rect 11149 44761 11161 44795
rect 11195 44792 11207 44795
rect 11517 44795 11575 44801
rect 11517 44792 11529 44795
rect 11195 44764 11529 44792
rect 11195 44761 11207 44764
rect 11149 44755 11207 44761
rect 11517 44761 11529 44764
rect 11563 44792 11575 44795
rect 12526 44792 12532 44804
rect 11563 44764 12532 44792
rect 11563 44761 11575 44764
rect 11517 44755 11575 44761
rect 12526 44752 12532 44764
rect 12584 44752 12590 44804
rect 15102 44752 15108 44804
rect 15160 44792 15166 44804
rect 15160 44764 15870 44792
rect 15160 44752 15166 44764
rect 8297 44727 8355 44733
rect 8297 44693 8309 44727
rect 8343 44724 8355 44727
rect 8478 44724 8484 44736
rect 8343 44696 8484 44724
rect 8343 44693 8355 44696
rect 8297 44687 8355 44693
rect 8478 44684 8484 44696
rect 8536 44684 8542 44736
rect 9766 44684 9772 44736
rect 9824 44684 9830 44736
rect 13354 44684 13360 44736
rect 13412 44684 13418 44736
rect 13449 44727 13507 44733
rect 13449 44693 13461 44727
rect 13495 44724 13507 44727
rect 15286 44724 15292 44736
rect 13495 44696 15292 44724
rect 13495 44693 13507 44696
rect 13449 44687 13507 44693
rect 15286 44684 15292 44696
rect 15344 44684 15350 44736
rect 15764 44724 15792 44764
rect 19794 44752 19800 44804
rect 19852 44752 19858 44804
rect 20254 44752 20260 44804
rect 20312 44752 20318 44804
rect 17126 44724 17132 44736
rect 15764 44696 17132 44724
rect 17126 44684 17132 44696
rect 17184 44684 17190 44736
rect 21266 44684 21272 44736
rect 21324 44684 21330 44736
rect 22066 44724 22094 44832
rect 22278 44820 22284 44872
rect 22336 44820 22342 44872
rect 22554 44752 22560 44804
rect 22612 44752 22618 44804
rect 23014 44792 23020 44804
rect 22940 44764 23020 44792
rect 22940 44724 22968 44764
rect 23014 44752 23020 44764
rect 23072 44752 23078 44804
rect 22066 44696 22968 44724
rect 23382 44684 23388 44736
rect 23440 44724 23446 44736
rect 24029 44727 24087 44733
rect 24029 44724 24041 44727
rect 23440 44696 24041 44724
rect 23440 44684 23446 44696
rect 24029 44693 24041 44696
rect 24075 44693 24087 44727
rect 24029 44687 24087 44693
rect 24486 44684 24492 44736
rect 24544 44724 24550 44736
rect 25498 44724 25504 44736
rect 24544 44696 25504 44724
rect 24544 44684 24550 44696
rect 25498 44684 25504 44696
rect 25556 44684 25562 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 5810 44480 5816 44532
rect 5868 44480 5874 44532
rect 6730 44480 6736 44532
rect 6788 44480 6794 44532
rect 7834 44480 7840 44532
rect 7892 44520 7898 44532
rect 8021 44523 8079 44529
rect 8021 44520 8033 44523
rect 7892 44492 8033 44520
rect 7892 44480 7898 44492
rect 8021 44489 8033 44492
rect 8067 44489 8079 44523
rect 8021 44483 8079 44489
rect 9674 44480 9680 44532
rect 9732 44520 9738 44532
rect 11057 44523 11115 44529
rect 11057 44520 11069 44523
rect 9732 44492 11069 44520
rect 9732 44480 9738 44492
rect 11057 44489 11069 44492
rect 11103 44489 11115 44523
rect 11057 44483 11115 44489
rect 11146 44480 11152 44532
rect 11204 44520 11210 44532
rect 11885 44523 11943 44529
rect 11885 44520 11897 44523
rect 11204 44492 11897 44520
rect 11204 44480 11210 44492
rect 11885 44489 11897 44492
rect 11931 44489 11943 44523
rect 11885 44483 11943 44489
rect 14458 44480 14464 44532
rect 14516 44520 14522 44532
rect 14921 44523 14979 44529
rect 14921 44520 14933 44523
rect 14516 44492 14933 44520
rect 14516 44480 14522 44492
rect 14921 44489 14933 44492
rect 14967 44489 14979 44523
rect 14921 44483 14979 44489
rect 15102 44480 15108 44532
rect 15160 44520 15166 44532
rect 15381 44523 15439 44529
rect 15381 44520 15393 44523
rect 15160 44492 15393 44520
rect 15160 44480 15166 44492
rect 15381 44489 15393 44492
rect 15427 44489 15439 44523
rect 15381 44483 15439 44489
rect 17512 44492 18460 44520
rect 7558 44412 7564 44464
rect 7616 44412 7622 44464
rect 12342 44412 12348 44464
rect 12400 44452 12406 44464
rect 12710 44452 12716 44464
rect 12400 44424 12716 44452
rect 12400 44412 12406 44424
rect 12710 44412 12716 44424
rect 12768 44412 12774 44464
rect 13446 44412 13452 44464
rect 13504 44412 13510 44464
rect 14090 44412 14096 44464
rect 14148 44412 14154 44464
rect 17126 44412 17132 44464
rect 17184 44452 17190 44464
rect 17512 44452 17540 44492
rect 18432 44452 18460 44492
rect 18598 44480 18604 44532
rect 18656 44520 18662 44532
rect 18782 44520 18788 44532
rect 18656 44492 18788 44520
rect 18656 44480 18662 44492
rect 18782 44480 18788 44492
rect 18840 44480 18846 44532
rect 19794 44480 19800 44532
rect 19852 44520 19858 44532
rect 20438 44520 20444 44532
rect 19852 44492 20444 44520
rect 19852 44480 19858 44492
rect 20438 44480 20444 44492
rect 20496 44520 20502 44532
rect 21269 44523 21327 44529
rect 21269 44520 21281 44523
rect 20496 44492 21281 44520
rect 20496 44480 20502 44492
rect 21269 44489 21281 44492
rect 21315 44489 21327 44523
rect 21269 44483 21327 44489
rect 22554 44480 22560 44532
rect 22612 44520 22618 44532
rect 24029 44523 24087 44529
rect 24029 44520 24041 44523
rect 22612 44492 24041 44520
rect 22612 44480 22618 44492
rect 24029 44489 24041 44492
rect 24075 44489 24087 44523
rect 24029 44483 24087 44489
rect 18877 44455 18935 44461
rect 18877 44452 18889 44455
rect 17184 44424 17618 44452
rect 18432 44424 18889 44452
rect 17184 44412 17190 44424
rect 18877 44421 18889 44424
rect 18923 44452 18935 44455
rect 20254 44452 20260 44464
rect 18923 44424 20260 44452
rect 18923 44421 18935 44424
rect 18877 44415 18935 44421
rect 20254 44412 20260 44424
rect 20312 44412 20318 44464
rect 21082 44412 21088 44464
rect 21140 44452 21146 44464
rect 21545 44455 21603 44461
rect 21545 44452 21557 44455
rect 21140 44424 21557 44452
rect 21140 44412 21146 44424
rect 21545 44421 21557 44424
rect 21591 44421 21603 44455
rect 21545 44415 21603 44421
rect 23014 44412 23020 44464
rect 23072 44412 23078 44464
rect 5258 44344 5264 44396
rect 5316 44384 5322 44396
rect 5997 44387 6055 44393
rect 5997 44384 6009 44387
rect 5316 44356 6009 44384
rect 5316 44344 5322 44356
rect 5997 44353 6009 44356
rect 6043 44353 6055 44387
rect 5997 44347 6055 44353
rect 6641 44387 6699 44393
rect 6641 44353 6653 44387
rect 6687 44384 6699 44387
rect 6730 44384 6736 44396
rect 6687 44356 6736 44384
rect 6687 44353 6699 44356
rect 6641 44347 6699 44353
rect 6730 44344 6736 44356
rect 6788 44344 6794 44396
rect 7098 44344 7104 44396
rect 7156 44384 7162 44396
rect 7377 44387 7435 44393
rect 7377 44384 7389 44387
rect 7156 44356 7389 44384
rect 7156 44344 7162 44356
rect 7377 44353 7389 44356
rect 7423 44353 7435 44387
rect 7377 44347 7435 44353
rect 7466 44344 7472 44396
rect 7524 44384 7530 44396
rect 8205 44387 8263 44393
rect 8205 44384 8217 44387
rect 7524 44356 8217 44384
rect 7524 44344 7530 44356
rect 8205 44353 8217 44356
rect 8251 44353 8263 44387
rect 8205 44347 8263 44353
rect 8941 44387 8999 44393
rect 8941 44353 8953 44387
rect 8987 44384 8999 44387
rect 10965 44387 11023 44393
rect 8987 44356 9536 44384
rect 8987 44353 8999 44356
rect 8941 44347 8999 44353
rect 7190 44276 7196 44328
rect 7248 44316 7254 44328
rect 9125 44319 9183 44325
rect 9125 44316 9137 44319
rect 7248 44288 9137 44316
rect 7248 44276 7254 44288
rect 9125 44285 9137 44288
rect 9171 44285 9183 44319
rect 9125 44279 9183 44285
rect 9508 44260 9536 44356
rect 10965 44353 10977 44387
rect 11011 44384 11023 44387
rect 11606 44384 11612 44396
rect 11011 44356 11612 44384
rect 11011 44353 11023 44356
rect 10965 44347 11023 44353
rect 11606 44344 11612 44356
rect 11664 44344 11670 44396
rect 12253 44387 12311 44393
rect 12253 44353 12265 44387
rect 12299 44384 12311 44387
rect 12728 44384 12756 44412
rect 13173 44387 13231 44393
rect 13173 44384 13185 44387
rect 12299 44356 12664 44384
rect 12728 44356 13185 44384
rect 12299 44353 12311 44356
rect 12253 44347 12311 44353
rect 11146 44276 11152 44328
rect 11204 44316 11210 44328
rect 12345 44319 12403 44325
rect 12345 44316 12357 44319
rect 11204 44288 12357 44316
rect 11204 44276 11210 44288
rect 12345 44285 12357 44288
rect 12391 44285 12403 44319
rect 12345 44279 12403 44285
rect 12437 44319 12495 44325
rect 12437 44285 12449 44319
rect 12483 44285 12495 44319
rect 12437 44279 12495 44285
rect 9490 44208 9496 44260
rect 9548 44208 9554 44260
rect 12158 44208 12164 44260
rect 12216 44248 12222 44260
rect 12452 44248 12480 44279
rect 12216 44220 12480 44248
rect 12216 44208 12222 44220
rect 11606 44140 11612 44192
rect 11664 44140 11670 44192
rect 12636 44180 12664 44356
rect 13173 44353 13185 44356
rect 13219 44353 13231 44387
rect 13173 44347 13231 44353
rect 24489 44387 24547 44393
rect 24489 44353 24501 44387
rect 24535 44384 24547 44387
rect 25314 44384 25320 44396
rect 24535 44356 25320 44384
rect 24535 44353 24547 44356
rect 24489 44347 24547 44353
rect 25314 44344 25320 44356
rect 25372 44344 25378 44396
rect 13446 44276 13452 44328
rect 13504 44316 13510 44328
rect 15197 44319 15255 44325
rect 15197 44316 15209 44319
rect 13504 44288 15209 44316
rect 13504 44276 13510 44288
rect 15197 44285 15209 44288
rect 15243 44316 15255 44319
rect 16666 44316 16672 44328
rect 15243 44288 16672 44316
rect 15243 44285 15255 44288
rect 15197 44279 15255 44285
rect 16666 44276 16672 44288
rect 16724 44276 16730 44328
rect 16758 44276 16764 44328
rect 16816 44316 16822 44328
rect 16853 44319 16911 44325
rect 16853 44316 16865 44319
rect 16816 44288 16865 44316
rect 16816 44276 16822 44288
rect 16853 44285 16865 44288
rect 16899 44285 16911 44319
rect 16853 44279 16911 44285
rect 17129 44319 17187 44325
rect 17129 44285 17141 44319
rect 17175 44316 17187 44319
rect 18966 44316 18972 44328
rect 17175 44288 18972 44316
rect 17175 44285 17187 44288
rect 17129 44279 17187 44285
rect 18966 44276 18972 44288
rect 19024 44276 19030 44328
rect 19518 44276 19524 44328
rect 19576 44276 19582 44328
rect 19797 44319 19855 44325
rect 19797 44285 19809 44319
rect 19843 44316 19855 44319
rect 21174 44316 21180 44328
rect 19843 44288 21180 44316
rect 19843 44285 19855 44288
rect 19797 44279 19855 44285
rect 21174 44276 21180 44288
rect 21232 44276 21238 44328
rect 22278 44276 22284 44328
rect 22336 44276 22342 44328
rect 22557 44319 22615 44325
rect 22557 44285 22569 44319
rect 22603 44316 22615 44319
rect 22922 44316 22928 44328
rect 22603 44288 22928 44316
rect 22603 44285 22615 44288
rect 22557 44279 22615 44285
rect 22922 44276 22928 44288
rect 22980 44276 22986 44328
rect 24762 44276 24768 44328
rect 24820 44276 24826 44328
rect 14550 44180 14556 44192
rect 12636 44152 14556 44180
rect 14550 44140 14556 44152
rect 14608 44140 14614 44192
rect 19536 44180 19564 44276
rect 22296 44248 22324 44276
rect 20824 44220 22324 44248
rect 20824 44180 20852 44220
rect 19536 44152 20852 44180
rect 22296 44180 22324 44220
rect 23290 44180 23296 44192
rect 22296 44152 23296 44180
rect 23290 44140 23296 44152
rect 23348 44140 23354 44192
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 8389 43979 8447 43985
rect 8389 43945 8401 43979
rect 8435 43976 8447 43979
rect 9398 43976 9404 43988
rect 8435 43948 9404 43976
rect 8435 43945 8447 43948
rect 8389 43939 8447 43945
rect 9398 43936 9404 43948
rect 9456 43936 9462 43988
rect 9950 43936 9956 43988
rect 10008 43976 10014 43988
rect 11609 43979 11667 43985
rect 11609 43976 11621 43979
rect 10008 43948 11621 43976
rect 10008 43936 10014 43948
rect 11609 43945 11621 43948
rect 11655 43945 11667 43979
rect 11609 43939 11667 43945
rect 18414 43936 18420 43988
rect 18472 43936 18478 43988
rect 21542 43936 21548 43988
rect 21600 43976 21606 43988
rect 21637 43979 21695 43985
rect 21637 43976 21649 43979
rect 21600 43948 21649 43976
rect 21600 43936 21606 43948
rect 21637 43945 21649 43948
rect 21683 43945 21695 43979
rect 21637 43939 21695 43945
rect 23290 43936 23296 43988
rect 23348 43976 23354 43988
rect 23474 43976 23480 43988
rect 23348 43948 23480 43976
rect 23348 43936 23354 43948
rect 23474 43936 23480 43948
rect 23532 43936 23538 43988
rect 23566 43936 23572 43988
rect 23624 43976 23630 43988
rect 24121 43979 24179 43985
rect 24121 43976 24133 43979
rect 23624 43948 24133 43976
rect 23624 43936 23630 43948
rect 24121 43945 24133 43948
rect 24167 43976 24179 43979
rect 24210 43976 24216 43988
rect 24167 43948 24216 43976
rect 24167 43945 24179 43948
rect 24121 43939 24179 43945
rect 24210 43936 24216 43948
rect 24268 43976 24274 43988
rect 25409 43979 25467 43985
rect 25409 43976 25421 43979
rect 24268 43948 25421 43976
rect 24268 43936 24274 43948
rect 25409 43945 25421 43948
rect 25455 43945 25467 43979
rect 25409 43939 25467 43945
rect 6917 43911 6975 43917
rect 6917 43877 6929 43911
rect 6963 43908 6975 43911
rect 7006 43908 7012 43920
rect 6963 43880 7012 43908
rect 6963 43877 6975 43880
rect 6917 43871 6975 43877
rect 7006 43868 7012 43880
rect 7064 43868 7070 43920
rect 16850 43868 16856 43920
rect 16908 43908 16914 43920
rect 18432 43908 18460 43936
rect 16908 43880 18460 43908
rect 16908 43868 16914 43880
rect 9125 43843 9183 43849
rect 9125 43809 9137 43843
rect 9171 43840 9183 43843
rect 9398 43840 9404 43852
rect 9171 43812 9404 43840
rect 9171 43809 9183 43812
rect 9125 43803 9183 43809
rect 9398 43800 9404 43812
rect 9456 43800 9462 43852
rect 9490 43800 9496 43852
rect 9548 43840 9554 43852
rect 18414 43840 18420 43852
rect 9548 43812 18420 43840
rect 9548 43800 9554 43812
rect 18414 43800 18420 43812
rect 18472 43800 18478 43852
rect 22186 43800 22192 43852
rect 22244 43840 22250 43852
rect 22465 43843 22523 43849
rect 22465 43840 22477 43843
rect 22244 43812 22477 43840
rect 22244 43800 22250 43812
rect 22465 43809 22477 43812
rect 22511 43809 22523 43843
rect 22465 43803 22523 43809
rect 22649 43843 22707 43849
rect 22649 43809 22661 43843
rect 22695 43840 22707 43843
rect 23290 43840 23296 43852
rect 22695 43812 23296 43840
rect 22695 43809 22707 43812
rect 22649 43803 22707 43809
rect 23290 43800 23296 43812
rect 23348 43800 23354 43852
rect 8573 43775 8631 43781
rect 8573 43741 8585 43775
rect 8619 43772 8631 43775
rect 9030 43772 9036 43784
rect 8619 43744 9036 43772
rect 8619 43741 8631 43744
rect 8573 43735 8631 43741
rect 9030 43732 9036 43744
rect 9088 43732 9094 43784
rect 6733 43707 6791 43713
rect 6733 43673 6745 43707
rect 6779 43704 6791 43707
rect 9401 43707 9459 43713
rect 6779 43676 7236 43704
rect 6779 43673 6791 43676
rect 6733 43667 6791 43673
rect 7208 43645 7236 43676
rect 9401 43673 9413 43707
rect 9447 43704 9459 43707
rect 10686 43704 10692 43716
rect 9447 43676 9812 43704
rect 10626 43676 10692 43704
rect 9447 43673 9459 43676
rect 9401 43667 9459 43673
rect 7193 43639 7251 43645
rect 7193 43605 7205 43639
rect 7239 43636 7251 43639
rect 8754 43636 8760 43648
rect 7239 43608 8760 43636
rect 7239 43605 7251 43608
rect 7193 43599 7251 43605
rect 8754 43596 8760 43608
rect 8812 43596 8818 43648
rect 9784 43636 9812 43676
rect 10686 43664 10692 43676
rect 10744 43664 10750 43716
rect 10796 43676 11008 43704
rect 10796 43636 10824 43676
rect 9784 43608 10824 43636
rect 10870 43596 10876 43648
rect 10928 43596 10934 43648
rect 10980 43636 11008 43676
rect 11422 43664 11428 43716
rect 11480 43704 11486 43716
rect 11517 43707 11575 43713
rect 11517 43704 11529 43707
rect 11480 43676 11529 43704
rect 11480 43664 11486 43676
rect 11517 43673 11529 43676
rect 11563 43704 11575 43707
rect 11977 43707 12035 43713
rect 11977 43704 11989 43707
rect 11563 43676 11989 43704
rect 11563 43673 11575 43676
rect 11517 43667 11575 43673
rect 11977 43673 11989 43676
rect 12023 43673 12035 43707
rect 11977 43667 12035 43673
rect 21542 43664 21548 43716
rect 21600 43704 21606 43716
rect 22373 43707 22431 43713
rect 22373 43704 22385 43707
rect 21600 43676 22385 43704
rect 21600 43664 21606 43676
rect 22373 43673 22385 43676
rect 22419 43673 22431 43707
rect 22373 43667 22431 43673
rect 16390 43636 16396 43648
rect 10980 43608 16396 43636
rect 16390 43596 16396 43608
rect 16448 43596 16454 43648
rect 17402 43596 17408 43648
rect 17460 43636 17466 43648
rect 17957 43639 18015 43645
rect 17957 43636 17969 43639
rect 17460 43608 17969 43636
rect 17460 43596 17466 43608
rect 17957 43605 17969 43608
rect 18003 43636 18015 43639
rect 19334 43636 19340 43648
rect 18003 43608 19340 43636
rect 18003 43605 18015 43608
rect 17957 43599 18015 43605
rect 19334 43596 19340 43608
rect 19392 43596 19398 43648
rect 21910 43596 21916 43648
rect 21968 43636 21974 43648
rect 22005 43639 22063 43645
rect 22005 43636 22017 43639
rect 21968 43608 22017 43636
rect 21968 43596 21974 43608
rect 22005 43605 22017 43608
rect 22051 43605 22063 43639
rect 22005 43599 22063 43605
rect 25314 43596 25320 43648
rect 25372 43596 25378 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 7742 43392 7748 43444
rect 7800 43392 7806 43444
rect 8573 43435 8631 43441
rect 8573 43401 8585 43435
rect 8619 43401 8631 43435
rect 8573 43395 8631 43401
rect 5350 43324 5356 43376
rect 5408 43364 5414 43376
rect 8588 43364 8616 43395
rect 8662 43392 8668 43444
rect 8720 43432 8726 43444
rect 9493 43435 9551 43441
rect 9493 43432 9505 43435
rect 8720 43404 9505 43432
rect 8720 43392 8726 43404
rect 9493 43401 9505 43404
rect 9539 43401 9551 43435
rect 9493 43395 9551 43401
rect 10410 43392 10416 43444
rect 10468 43432 10474 43444
rect 10597 43435 10655 43441
rect 10597 43432 10609 43435
rect 10468 43404 10609 43432
rect 10468 43392 10474 43404
rect 10597 43401 10609 43404
rect 10643 43401 10655 43435
rect 10597 43395 10655 43401
rect 14734 43392 14740 43444
rect 14792 43432 14798 43444
rect 15013 43435 15071 43441
rect 15013 43432 15025 43435
rect 14792 43404 15025 43432
rect 14792 43392 14798 43404
rect 15013 43401 15025 43404
rect 15059 43401 15071 43435
rect 15013 43395 15071 43401
rect 15105 43435 15163 43441
rect 15105 43401 15117 43435
rect 15151 43432 15163 43435
rect 15562 43432 15568 43444
rect 15151 43404 15568 43432
rect 15151 43401 15163 43404
rect 15105 43395 15163 43401
rect 15562 43392 15568 43404
rect 15620 43432 15626 43444
rect 15657 43435 15715 43441
rect 15657 43432 15669 43435
rect 15620 43404 15669 43432
rect 15620 43392 15626 43404
rect 15657 43401 15669 43404
rect 15703 43401 15715 43435
rect 15657 43395 15715 43401
rect 17402 43392 17408 43444
rect 17460 43392 17466 43444
rect 17494 43392 17500 43444
rect 17552 43392 17558 43444
rect 20070 43392 20076 43444
rect 20128 43392 20134 43444
rect 20441 43435 20499 43441
rect 20441 43401 20453 43435
rect 20487 43432 20499 43435
rect 20898 43432 20904 43444
rect 20487 43404 20904 43432
rect 20487 43401 20499 43404
rect 20441 43395 20499 43401
rect 5408 43336 8616 43364
rect 5408 43324 5414 43336
rect 9122 43324 9128 43376
rect 9180 43364 9186 43376
rect 9585 43367 9643 43373
rect 9585 43364 9597 43367
rect 9180 43336 9597 43364
rect 9180 43324 9186 43336
rect 9585 43333 9597 43336
rect 9631 43333 9643 43367
rect 9585 43327 9643 43333
rect 10686 43324 10692 43376
rect 10744 43364 10750 43376
rect 10962 43364 10968 43376
rect 10744 43336 10968 43364
rect 10744 43324 10750 43336
rect 10962 43324 10968 43336
rect 11020 43364 11026 43376
rect 11057 43367 11115 43373
rect 11057 43364 11069 43367
rect 11020 43336 11069 43364
rect 11020 43324 11026 43336
rect 11057 43333 11069 43336
rect 11103 43333 11115 43367
rect 11057 43327 11115 43333
rect 12618 43324 12624 43376
rect 12676 43324 12682 43376
rect 14090 43364 14096 43376
rect 13846 43336 14096 43364
rect 14090 43324 14096 43336
rect 14148 43364 14154 43376
rect 16206 43364 16212 43376
rect 14148 43336 16212 43364
rect 14148 43324 14154 43336
rect 16206 43324 16212 43336
rect 16264 43364 16270 43376
rect 16669 43367 16727 43373
rect 16669 43364 16681 43367
rect 16264 43336 16681 43364
rect 16264 43324 16270 43336
rect 16669 43333 16681 43336
rect 16715 43333 16727 43367
rect 20456 43364 20484 43395
rect 20898 43392 20904 43404
rect 20956 43432 20962 43444
rect 21082 43432 21088 43444
rect 20956 43404 21088 43432
rect 20956 43392 20962 43404
rect 21082 43392 21088 43404
rect 21140 43432 21146 43444
rect 21361 43435 21419 43441
rect 21361 43432 21373 43435
rect 21140 43404 21373 43432
rect 21140 43392 21146 43404
rect 21361 43401 21373 43404
rect 21407 43401 21419 43435
rect 21361 43395 21419 43401
rect 21634 43392 21640 43444
rect 21692 43432 21698 43444
rect 21692 43404 22094 43432
rect 21692 43392 21698 43404
rect 19826 43336 20484 43364
rect 16669 43327 16727 43333
rect 1302 43256 1308 43308
rect 1360 43296 1366 43308
rect 1673 43299 1731 43305
rect 1673 43296 1685 43299
rect 1360 43268 1685 43296
rect 1360 43256 1366 43268
rect 1673 43265 1685 43268
rect 1719 43296 1731 43299
rect 2133 43299 2191 43305
rect 2133 43296 2145 43299
rect 1719 43268 2145 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 2133 43265 2145 43268
rect 2179 43265 2191 43299
rect 2133 43259 2191 43265
rect 7650 43256 7656 43308
rect 7708 43296 7714 43308
rect 7929 43299 7987 43305
rect 7929 43296 7941 43299
rect 7708 43268 7941 43296
rect 7708 43256 7714 43268
rect 7929 43265 7941 43268
rect 7975 43265 7987 43299
rect 7929 43259 7987 43265
rect 8386 43256 8392 43308
rect 8444 43296 8450 43308
rect 8481 43299 8539 43305
rect 8481 43296 8493 43299
rect 8444 43268 8493 43296
rect 8444 43256 8450 43268
rect 8481 43265 8493 43268
rect 8527 43265 8539 43299
rect 8481 43259 8539 43265
rect 8754 43256 8760 43308
rect 8812 43296 8818 43308
rect 9766 43296 9772 43308
rect 8812 43268 9772 43296
rect 8812 43256 8818 43268
rect 9766 43256 9772 43268
rect 9824 43256 9830 43308
rect 10318 43256 10324 43308
rect 10376 43296 10382 43308
rect 10505 43299 10563 43305
rect 10505 43296 10517 43299
rect 10376 43268 10517 43296
rect 10376 43256 10382 43268
rect 10505 43265 10517 43268
rect 10551 43265 10563 43299
rect 10505 43259 10563 43265
rect 14642 43256 14648 43308
rect 14700 43296 14706 43308
rect 22066 43296 22094 43404
rect 22370 43392 22376 43444
rect 22428 43432 22434 43444
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 22428 43404 22477 43432
rect 22428 43392 22434 43404
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 24210 43392 24216 43444
rect 24268 43392 24274 43444
rect 22186 43324 22192 43376
rect 22244 43364 22250 43376
rect 22738 43364 22744 43376
rect 22244 43336 22744 43364
rect 22244 43324 22250 43336
rect 22738 43324 22744 43336
rect 22796 43324 22802 43376
rect 23566 43324 23572 43376
rect 23624 43364 23630 43376
rect 23845 43367 23903 43373
rect 23845 43364 23857 43367
rect 23624 43336 23857 43364
rect 23624 43324 23630 43336
rect 23845 43333 23857 43336
rect 23891 43333 23903 43367
rect 24228 43364 24256 43392
rect 24228 43336 24334 43364
rect 23845 43327 23903 43333
rect 22373 43299 22431 43305
rect 22373 43296 22385 43299
rect 14700 43268 15240 43296
rect 22066 43268 22385 43296
rect 14700 43256 14706 43268
rect 8846 43188 8852 43240
rect 8904 43228 8910 43240
rect 9306 43228 9312 43240
rect 8904 43200 9312 43228
rect 8904 43188 8910 43200
rect 9306 43188 9312 43200
rect 9364 43228 9370 43240
rect 9490 43228 9496 43240
rect 9364 43200 9496 43228
rect 9364 43188 9370 43200
rect 9490 43188 9496 43200
rect 9548 43228 9554 43240
rect 9677 43231 9735 43237
rect 9677 43228 9689 43231
rect 9548 43200 9689 43228
rect 9548 43188 9554 43200
rect 9677 43197 9689 43200
rect 9723 43197 9735 43231
rect 9677 43191 9735 43197
rect 12342 43188 12348 43240
rect 12400 43188 12406 43240
rect 15212 43237 15240 43268
rect 22373 43265 22385 43268
rect 22419 43265 22431 43299
rect 22373 43259 22431 43265
rect 15197 43231 15255 43237
rect 15197 43197 15209 43231
rect 15243 43197 15255 43231
rect 15197 43191 15255 43197
rect 15654 43188 15660 43240
rect 15712 43228 15718 43240
rect 17678 43228 17684 43240
rect 15712 43200 17684 43228
rect 15712 43188 15718 43200
rect 17678 43188 17684 43200
rect 17736 43188 17742 43240
rect 18322 43188 18328 43240
rect 18380 43188 18386 43240
rect 18601 43231 18659 43237
rect 18601 43197 18613 43231
rect 18647 43228 18659 43231
rect 19610 43228 19616 43240
rect 18647 43200 19616 43228
rect 18647 43197 18659 43200
rect 18601 43191 18659 43197
rect 19610 43188 19616 43200
rect 19668 43228 19674 43240
rect 21266 43228 21272 43240
rect 19668 43200 21272 43228
rect 19668 43188 19674 43200
rect 21266 43188 21272 43200
rect 21324 43188 21330 43240
rect 22649 43231 22707 43237
rect 22649 43197 22661 43231
rect 22695 43228 22707 43231
rect 22738 43228 22744 43240
rect 22695 43200 22744 43228
rect 22695 43197 22707 43200
rect 22649 43191 22707 43197
rect 22738 43188 22744 43200
rect 22796 43188 22802 43240
rect 23474 43188 23480 43240
rect 23532 43228 23538 43240
rect 23569 43231 23627 43237
rect 23569 43228 23581 43231
rect 23532 43200 23581 43228
rect 23532 43188 23538 43200
rect 23569 43197 23581 43200
rect 23615 43197 23627 43231
rect 23569 43191 23627 43197
rect 1857 43163 1915 43169
rect 1857 43129 1869 43163
rect 1903 43160 1915 43163
rect 3970 43160 3976 43172
rect 1903 43132 3976 43160
rect 1903 43129 1915 43132
rect 1857 43123 1915 43129
rect 3970 43120 3976 43132
rect 4028 43120 4034 43172
rect 9125 43163 9183 43169
rect 9125 43129 9137 43163
rect 9171 43160 9183 43163
rect 11146 43160 11152 43172
rect 9171 43132 11152 43160
rect 9171 43129 9183 43132
rect 9125 43123 9183 43129
rect 11146 43120 11152 43132
rect 11204 43120 11210 43172
rect 13722 43120 13728 43172
rect 13780 43160 13786 43172
rect 14645 43163 14703 43169
rect 14645 43160 14657 43163
rect 13780 43132 14657 43160
rect 13780 43120 13786 43132
rect 14645 43129 14657 43132
rect 14691 43129 14703 43163
rect 14645 43123 14703 43129
rect 16758 43120 16764 43172
rect 16816 43160 16822 43172
rect 18340 43160 18368 43188
rect 16816 43132 18368 43160
rect 16816 43120 16822 43132
rect 13906 43052 13912 43104
rect 13964 43092 13970 43104
rect 14093 43095 14151 43101
rect 14093 43092 14105 43095
rect 13964 43064 14105 43092
rect 13964 43052 13970 43064
rect 14093 43061 14105 43064
rect 14139 43061 14151 43095
rect 14093 43055 14151 43061
rect 17034 43052 17040 43104
rect 17092 43052 17098 43104
rect 18340 43092 18368 43132
rect 19242 43092 19248 43104
rect 18340 43064 19248 43092
rect 19242 43052 19248 43064
rect 19300 43052 19306 43104
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 24946 43092 24952 43104
rect 22051 43064 24952 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 24946 43052 24952 43064
rect 25004 43052 25010 43104
rect 25130 43052 25136 43104
rect 25188 43092 25194 43104
rect 25317 43095 25375 43101
rect 25317 43092 25329 43095
rect 25188 43064 25329 43092
rect 25188 43052 25194 43064
rect 25317 43061 25329 43064
rect 25363 43061 25375 43095
rect 25317 43055 25375 43061
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 8662 42848 8668 42900
rect 8720 42848 8726 42900
rect 8846 42848 8852 42900
rect 8904 42888 8910 42900
rect 8941 42891 8999 42897
rect 8941 42888 8953 42891
rect 8904 42860 8953 42888
rect 8904 42848 8910 42860
rect 8941 42857 8953 42860
rect 8987 42857 8999 42891
rect 8941 42851 8999 42857
rect 9122 42848 9128 42900
rect 9180 42888 9186 42900
rect 9490 42888 9496 42900
rect 9180 42860 9496 42888
rect 9180 42848 9186 42860
rect 9490 42848 9496 42860
rect 9548 42848 9554 42900
rect 9585 42891 9643 42897
rect 9585 42857 9597 42891
rect 9631 42888 9643 42891
rect 10686 42888 10692 42900
rect 9631 42860 10692 42888
rect 9631 42857 9643 42860
rect 9585 42851 9643 42857
rect 9600 42820 9628 42851
rect 10686 42848 10692 42860
rect 10744 42848 10750 42900
rect 12897 42891 12955 42897
rect 12897 42857 12909 42891
rect 12943 42888 12955 42891
rect 14090 42888 14096 42900
rect 12943 42860 14096 42888
rect 12943 42857 12955 42860
rect 12897 42851 12955 42857
rect 9140 42792 9628 42820
rect 9140 42764 9168 42792
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 4985 42755 5043 42761
rect 4985 42752 4997 42755
rect 4948 42724 4997 42752
rect 4948 42712 4954 42724
rect 4985 42721 4997 42724
rect 5031 42721 5043 42755
rect 4985 42715 5043 42721
rect 9122 42712 9128 42764
rect 9180 42712 9186 42764
rect 9214 42712 9220 42764
rect 9272 42752 9278 42764
rect 9309 42755 9367 42761
rect 9309 42752 9321 42755
rect 9272 42724 9321 42752
rect 9272 42712 9278 42724
rect 9309 42721 9321 42724
rect 9355 42721 9367 42755
rect 9309 42715 9367 42721
rect 9398 42712 9404 42764
rect 9456 42752 9462 42764
rect 10781 42755 10839 42761
rect 10781 42752 10793 42755
rect 9456 42724 10793 42752
rect 9456 42712 9462 42724
rect 10781 42721 10793 42724
rect 10827 42752 10839 42755
rect 12342 42752 12348 42764
rect 10827 42724 12348 42752
rect 10827 42721 10839 42724
rect 10781 42715 10839 42721
rect 12342 42712 12348 42724
rect 12400 42712 12406 42764
rect 12912 42684 12940 42851
rect 14090 42848 14096 42860
rect 14148 42888 14154 42900
rect 14277 42891 14335 42897
rect 14277 42888 14289 42891
rect 14148 42860 14289 42888
rect 14148 42848 14154 42860
rect 14277 42857 14289 42860
rect 14323 42857 14335 42891
rect 14277 42851 14335 42857
rect 19784 42891 19842 42897
rect 19784 42857 19796 42891
rect 19830 42888 19842 42891
rect 20346 42888 20352 42900
rect 19830 42860 20352 42888
rect 19830 42857 19842 42860
rect 19784 42851 19842 42857
rect 20346 42848 20352 42860
rect 20404 42888 20410 42900
rect 21450 42888 21456 42900
rect 20404 42860 21456 42888
rect 20404 42848 20410 42860
rect 21450 42848 21456 42860
rect 21508 42848 21514 42900
rect 24210 42848 24216 42900
rect 24268 42888 24274 42900
rect 25317 42891 25375 42897
rect 25317 42888 25329 42891
rect 24268 42860 25329 42888
rect 24268 42848 24274 42860
rect 25317 42857 25329 42860
rect 25363 42857 25375 42891
rect 25317 42851 25375 42857
rect 21634 42780 21640 42832
rect 21692 42820 21698 42832
rect 23431 42823 23489 42829
rect 23431 42820 23443 42823
rect 21692 42792 23443 42820
rect 21692 42780 21698 42792
rect 23431 42789 23443 42792
rect 23477 42789 23489 42823
rect 23431 42783 23489 42789
rect 14829 42755 14887 42761
rect 14829 42721 14841 42755
rect 14875 42752 14887 42755
rect 16758 42752 16764 42764
rect 14875 42724 16764 42752
rect 14875 42721 14887 42724
rect 14829 42715 14887 42721
rect 16758 42712 16764 42724
rect 16816 42712 16822 42764
rect 17773 42755 17831 42761
rect 17773 42721 17785 42755
rect 17819 42752 17831 42755
rect 18141 42755 18199 42761
rect 18141 42752 18153 42755
rect 17819 42724 18153 42752
rect 17819 42721 17831 42724
rect 17773 42715 17831 42721
rect 18141 42721 18153 42724
rect 18187 42752 18199 42755
rect 18414 42752 18420 42764
rect 18187 42724 18420 42752
rect 18187 42721 18199 42724
rect 18141 42715 18199 42721
rect 18414 42712 18420 42724
rect 18472 42712 18478 42764
rect 19521 42755 19579 42761
rect 19521 42721 19533 42755
rect 19567 42752 19579 42755
rect 19567 42724 21864 42752
rect 19567 42721 19579 42724
rect 19521 42715 19579 42721
rect 12190 42656 12940 42684
rect 16206 42644 16212 42696
rect 16264 42644 16270 42696
rect 17589 42687 17647 42693
rect 17589 42653 17601 42687
rect 17635 42684 17647 42687
rect 18325 42687 18383 42693
rect 18325 42684 18337 42687
rect 17635 42656 18337 42684
rect 17635 42653 17647 42656
rect 17589 42647 17647 42653
rect 18325 42653 18337 42656
rect 18371 42684 18383 42687
rect 18598 42684 18604 42696
rect 18371 42656 18604 42684
rect 18371 42653 18383 42656
rect 18325 42647 18383 42653
rect 18598 42644 18604 42656
rect 18656 42684 18662 42696
rect 19058 42684 19064 42696
rect 18656 42656 19064 42684
rect 18656 42644 18662 42656
rect 19058 42644 19064 42656
rect 19116 42644 19122 42696
rect 20898 42644 20904 42696
rect 20956 42644 20962 42696
rect 21836 42684 21864 42724
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22281 42755 22339 42761
rect 22281 42752 22293 42755
rect 22060 42724 22293 42752
rect 22060 42712 22066 42724
rect 22281 42721 22293 42724
rect 22327 42721 22339 42755
rect 22281 42715 22339 42721
rect 22465 42755 22523 42761
rect 22465 42721 22477 42755
rect 22511 42752 22523 42755
rect 22554 42752 22560 42764
rect 22511 42724 22560 42752
rect 22511 42721 22523 42724
rect 22465 42715 22523 42721
rect 22554 42712 22560 42724
rect 22612 42712 22618 42764
rect 23106 42712 23112 42764
rect 23164 42752 23170 42764
rect 24854 42752 24860 42764
rect 23164 42724 24860 42752
rect 23164 42712 23170 42724
rect 24854 42712 24860 42724
rect 24912 42712 24918 42764
rect 22830 42684 22836 42696
rect 21836 42656 22836 42684
rect 22830 42644 22836 42656
rect 22888 42644 22894 42696
rect 23201 42687 23259 42693
rect 23201 42653 23213 42687
rect 23247 42653 23259 42687
rect 23201 42647 23259 42653
rect 4798 42576 4804 42628
rect 4856 42616 4862 42628
rect 5261 42619 5319 42625
rect 5261 42616 5273 42619
rect 4856 42588 5273 42616
rect 4856 42576 4862 42588
rect 5261 42585 5273 42588
rect 5307 42585 5319 42619
rect 5261 42579 5319 42585
rect 9674 42576 9680 42628
rect 9732 42616 9738 42628
rect 11057 42619 11115 42625
rect 11057 42616 11069 42619
rect 9732 42588 11069 42616
rect 9732 42576 9738 42588
rect 11057 42585 11069 42588
rect 11103 42585 11115 42619
rect 15105 42619 15163 42625
rect 15105 42616 15117 42619
rect 11057 42579 11115 42585
rect 12544 42588 15117 42616
rect 8297 42551 8355 42557
rect 8297 42517 8309 42551
rect 8343 42548 8355 42551
rect 8386 42548 8392 42560
rect 8343 42520 8392 42548
rect 8343 42517 8355 42520
rect 8297 42511 8355 42517
rect 8386 42508 8392 42520
rect 8444 42508 8450 42560
rect 10318 42508 10324 42560
rect 10376 42508 10382 42560
rect 12434 42508 12440 42560
rect 12492 42548 12498 42560
rect 12544 42557 12572 42588
rect 15105 42585 15117 42588
rect 15151 42585 15163 42619
rect 17497 42619 17555 42625
rect 15105 42579 15163 42585
rect 16408 42588 17172 42616
rect 12529 42551 12587 42557
rect 12529 42548 12541 42551
rect 12492 42520 12541 42548
rect 12492 42508 12498 42520
rect 12529 42517 12541 42520
rect 12575 42517 12587 42551
rect 12529 42511 12587 42517
rect 14550 42508 14556 42560
rect 14608 42548 14614 42560
rect 16408 42548 16436 42588
rect 14608 42520 16436 42548
rect 16577 42551 16635 42557
rect 14608 42508 14614 42520
rect 16577 42517 16589 42551
rect 16623 42548 16635 42551
rect 16758 42548 16764 42560
rect 16623 42520 16764 42548
rect 16623 42517 16635 42520
rect 16577 42511 16635 42517
rect 16758 42508 16764 42520
rect 16816 42508 16822 42560
rect 17144 42557 17172 42588
rect 17497 42585 17509 42619
rect 17543 42616 17555 42619
rect 17543 42588 19748 42616
rect 17543 42585 17555 42588
rect 17497 42579 17555 42585
rect 17129 42551 17187 42557
rect 17129 42517 17141 42551
rect 17175 42517 17187 42551
rect 19720 42548 19748 42588
rect 21082 42576 21088 42628
rect 21140 42616 21146 42628
rect 22189 42619 22247 42625
rect 22189 42616 22201 42619
rect 21140 42588 22201 42616
rect 21140 42576 21146 42588
rect 22189 42585 22201 42588
rect 22235 42585 22247 42619
rect 23216 42616 23244 42647
rect 23216 42588 24532 42616
rect 22189 42579 22247 42585
rect 20438 42548 20444 42560
rect 19720 42520 20444 42548
rect 17129 42511 17187 42517
rect 20438 42508 20444 42520
rect 20496 42508 20502 42560
rect 21266 42508 21272 42560
rect 21324 42508 21330 42560
rect 21821 42551 21879 42557
rect 21821 42517 21833 42551
rect 21867 42548 21879 42551
rect 22094 42548 22100 42560
rect 21867 42520 22100 42548
rect 21867 42517 21879 42520
rect 21821 42511 21879 42517
rect 22094 42508 22100 42520
rect 22152 42508 22158 42560
rect 24504 42557 24532 42588
rect 24489 42551 24547 42557
rect 24489 42517 24501 42551
rect 24535 42548 24547 42551
rect 24854 42548 24860 42560
rect 24535 42520 24860 42548
rect 24535 42517 24547 42520
rect 24489 42511 24547 42517
rect 24854 42508 24860 42520
rect 24912 42508 24918 42560
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 4154 42304 4160 42356
rect 4212 42344 4218 42356
rect 4341 42347 4399 42353
rect 4341 42344 4353 42347
rect 4212 42316 4353 42344
rect 4212 42304 4218 42316
rect 4341 42313 4353 42316
rect 4387 42313 4399 42347
rect 4341 42307 4399 42313
rect 5074 42304 5080 42356
rect 5132 42304 5138 42356
rect 5442 42304 5448 42356
rect 5500 42344 5506 42356
rect 6733 42347 6791 42353
rect 6733 42344 6745 42347
rect 5500 42316 6745 42344
rect 5500 42304 5506 42316
rect 6733 42313 6745 42316
rect 6779 42313 6791 42347
rect 8110 42344 8116 42356
rect 6733 42307 6791 42313
rect 7576 42316 8116 42344
rect 7576 42276 7604 42316
rect 8110 42304 8116 42316
rect 8168 42344 8174 42356
rect 9214 42344 9220 42356
rect 8168 42316 9220 42344
rect 8168 42304 8174 42316
rect 9214 42304 9220 42316
rect 9272 42304 9278 42356
rect 9582 42304 9588 42356
rect 9640 42344 9646 42356
rect 9677 42347 9735 42353
rect 9677 42344 9689 42347
rect 9640 42316 9689 42344
rect 9640 42304 9646 42316
rect 9677 42313 9689 42316
rect 9723 42313 9735 42347
rect 9677 42307 9735 42313
rect 11790 42304 11796 42356
rect 11848 42304 11854 42356
rect 12989 42347 13047 42353
rect 12989 42313 13001 42347
rect 13035 42344 13047 42347
rect 13354 42344 13360 42356
rect 13035 42316 13360 42344
rect 13035 42313 13047 42316
rect 12989 42307 13047 42313
rect 13354 42304 13360 42316
rect 13412 42304 13418 42356
rect 15286 42304 15292 42356
rect 15344 42344 15350 42356
rect 15381 42347 15439 42353
rect 15381 42344 15393 42347
rect 15344 42316 15393 42344
rect 15344 42304 15350 42316
rect 15381 42313 15393 42316
rect 15427 42313 15439 42347
rect 15381 42307 15439 42313
rect 15841 42347 15899 42353
rect 15841 42313 15853 42347
rect 15887 42344 15899 42347
rect 16853 42347 16911 42353
rect 16853 42344 16865 42347
rect 15887 42316 16865 42344
rect 15887 42313 15899 42316
rect 15841 42307 15899 42313
rect 16853 42313 16865 42316
rect 16899 42313 16911 42347
rect 16853 42307 16911 42313
rect 17221 42347 17279 42353
rect 17221 42313 17233 42347
rect 17267 42344 17279 42347
rect 18141 42347 18199 42353
rect 18141 42344 18153 42347
rect 17267 42316 18153 42344
rect 17267 42313 17279 42316
rect 17221 42307 17279 42313
rect 18141 42313 18153 42316
rect 18187 42344 18199 42347
rect 20530 42344 20536 42356
rect 18187 42316 20536 42344
rect 18187 42313 18199 42316
rect 18141 42307 18199 42313
rect 20530 42304 20536 42316
rect 20588 42304 20594 42356
rect 20898 42304 20904 42356
rect 20956 42344 20962 42356
rect 21269 42347 21327 42353
rect 21269 42344 21281 42347
rect 20956 42316 21281 42344
rect 20956 42304 20962 42316
rect 21269 42313 21281 42316
rect 21315 42313 21327 42347
rect 21269 42307 21327 42313
rect 22370 42304 22376 42356
rect 22428 42344 22434 42356
rect 23290 42344 23296 42356
rect 22428 42316 23296 42344
rect 22428 42304 22434 42316
rect 23290 42304 23296 42316
rect 23348 42344 23354 42356
rect 25225 42347 25283 42353
rect 25225 42344 25237 42347
rect 23348 42316 25237 42344
rect 23348 42304 23354 42316
rect 25225 42313 25237 42316
rect 25271 42313 25283 42347
rect 25225 42307 25283 42313
rect 9122 42276 9128 42288
rect 7484 42248 7604 42276
rect 8970 42248 9128 42276
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42208 3939 42211
rect 4246 42208 4252 42220
rect 3927 42180 4252 42208
rect 3927 42177 3939 42180
rect 3881 42171 3939 42177
rect 4246 42168 4252 42180
rect 4304 42168 4310 42220
rect 4985 42211 5043 42217
rect 4985 42177 4997 42211
rect 5031 42208 5043 42211
rect 6641 42211 6699 42217
rect 5031 42180 5580 42208
rect 5031 42177 5043 42180
rect 4985 42171 5043 42177
rect 5552 42013 5580 42180
rect 6641 42177 6653 42211
rect 6687 42208 6699 42211
rect 7190 42208 7196 42220
rect 6687 42180 7196 42208
rect 6687 42177 6699 42180
rect 6641 42171 6699 42177
rect 7190 42168 7196 42180
rect 7248 42168 7254 42220
rect 7484 42217 7512 42248
rect 9122 42236 9128 42248
rect 9180 42236 9186 42288
rect 10137 42279 10195 42285
rect 10137 42245 10149 42279
rect 10183 42276 10195 42279
rect 11882 42276 11888 42288
rect 10183 42248 11888 42276
rect 10183 42245 10195 42248
rect 10137 42239 10195 42245
rect 11882 42236 11888 42248
rect 11940 42236 11946 42288
rect 12253 42279 12311 42285
rect 12253 42245 12265 42279
rect 12299 42276 12311 42279
rect 15562 42276 15568 42288
rect 12299 42248 15568 42276
rect 12299 42245 12311 42248
rect 12253 42239 12311 42245
rect 15562 42236 15568 42248
rect 15620 42236 15626 42288
rect 15749 42279 15807 42285
rect 15749 42245 15761 42279
rect 15795 42276 15807 42279
rect 17402 42276 17408 42288
rect 15795 42248 17408 42276
rect 15795 42245 15807 42248
rect 15749 42239 15807 42245
rect 17402 42236 17408 42248
rect 17460 42236 17466 42288
rect 20714 42276 20720 42288
rect 18892 42248 20720 42276
rect 7469 42211 7527 42217
rect 7469 42177 7481 42211
rect 7515 42177 7527 42211
rect 9582 42208 9588 42220
rect 7469 42171 7527 42177
rect 8956 42180 9588 42208
rect 7742 42100 7748 42152
rect 7800 42140 7806 42152
rect 8956 42140 8984 42180
rect 9582 42168 9588 42180
rect 9640 42168 9646 42220
rect 10045 42211 10103 42217
rect 10045 42177 10057 42211
rect 10091 42177 10103 42211
rect 10045 42171 10103 42177
rect 10060 42140 10088 42171
rect 11146 42168 11152 42220
rect 11204 42208 11210 42220
rect 12161 42211 12219 42217
rect 12161 42208 12173 42211
rect 11204 42180 12173 42208
rect 11204 42168 11210 42180
rect 12161 42177 12173 42180
rect 12207 42177 12219 42211
rect 12161 42171 12219 42177
rect 13357 42211 13415 42217
rect 13357 42177 13369 42211
rect 13403 42208 13415 42211
rect 14185 42211 14243 42217
rect 14185 42208 14197 42211
rect 13403 42180 14197 42208
rect 13403 42177 13415 42180
rect 13357 42171 13415 42177
rect 14185 42177 14197 42180
rect 14231 42177 14243 42211
rect 14185 42171 14243 42177
rect 16666 42168 16672 42220
rect 16724 42208 16730 42220
rect 18892 42217 18920 42248
rect 20714 42236 20720 42248
rect 20772 42276 20778 42288
rect 21545 42279 21603 42285
rect 21545 42276 21557 42279
rect 20772 42248 21557 42276
rect 20772 42236 20778 42248
rect 21545 42245 21557 42248
rect 21591 42276 21603 42279
rect 22005 42279 22063 42285
rect 22005 42276 22017 42279
rect 21591 42248 22017 42276
rect 21591 42245 21603 42248
rect 21545 42239 21603 42245
rect 22005 42245 22017 42248
rect 22051 42245 22063 42279
rect 22005 42239 22063 42245
rect 24210 42236 24216 42288
rect 24268 42236 24274 42288
rect 17865 42211 17923 42217
rect 17865 42208 17877 42211
rect 16724 42180 17877 42208
rect 16724 42168 16730 42180
rect 7800 42112 8984 42140
rect 9048 42112 10088 42140
rect 10229 42143 10287 42149
rect 7800 42100 7806 42112
rect 5537 42007 5595 42013
rect 5537 41973 5549 42007
rect 5583 42004 5595 42007
rect 6362 42004 6368 42016
rect 5583 41976 6368 42004
rect 5583 41973 5595 41976
rect 5537 41967 5595 41973
rect 6362 41964 6368 41976
rect 6420 41964 6426 42016
rect 7190 41964 7196 42016
rect 7248 41964 7254 42016
rect 7558 41964 7564 42016
rect 7616 42004 7622 42016
rect 9048 42004 9076 42112
rect 10229 42109 10241 42143
rect 10275 42109 10287 42143
rect 10229 42103 10287 42109
rect 9582 42032 9588 42084
rect 9640 42072 9646 42084
rect 10244 42072 10272 42103
rect 12434 42100 12440 42152
rect 12492 42100 12498 42152
rect 13449 42143 13507 42149
rect 13449 42140 13461 42143
rect 13372 42112 13461 42140
rect 13372 42084 13400 42112
rect 13449 42109 13461 42112
rect 13495 42109 13507 42143
rect 13449 42103 13507 42109
rect 13633 42143 13691 42149
rect 13633 42109 13645 42143
rect 13679 42140 13691 42143
rect 14458 42140 14464 42152
rect 13679 42112 14464 42140
rect 13679 42109 13691 42112
rect 13633 42103 13691 42109
rect 14458 42100 14464 42112
rect 14516 42140 14522 42152
rect 17420 42149 17448 42180
rect 17865 42177 17877 42180
rect 17911 42177 17923 42211
rect 17865 42171 17923 42177
rect 18601 42211 18659 42217
rect 18601 42177 18613 42211
rect 18647 42208 18659 42211
rect 18877 42211 18935 42217
rect 18877 42208 18889 42211
rect 18647 42180 18889 42208
rect 18647 42177 18659 42180
rect 18601 42171 18659 42177
rect 18877 42177 18889 42180
rect 18923 42177 18935 42211
rect 18877 42171 18935 42177
rect 15933 42143 15991 42149
rect 15933 42140 15945 42143
rect 14516 42112 15945 42140
rect 14516 42100 14522 42112
rect 15933 42109 15945 42112
rect 15979 42109 15991 42143
rect 15933 42103 15991 42109
rect 17313 42143 17371 42149
rect 17313 42109 17325 42143
rect 17359 42109 17371 42143
rect 17313 42103 17371 42109
rect 17405 42143 17463 42149
rect 17405 42109 17417 42143
rect 17451 42109 17463 42143
rect 17880 42140 17908 42171
rect 20622 42168 20628 42220
rect 20680 42168 20686 42220
rect 20990 42208 20996 42220
rect 20732 42180 20996 42208
rect 19058 42140 19064 42152
rect 17880 42112 19064 42140
rect 17405 42103 17463 42109
rect 9640 42044 10272 42072
rect 9640 42032 9646 42044
rect 13354 42032 13360 42084
rect 13412 42032 13418 42084
rect 7616 41976 9076 42004
rect 9217 42007 9275 42013
rect 7616 41964 7622 41976
rect 9217 41973 9229 42007
rect 9263 42004 9275 42007
rect 9674 42004 9680 42016
rect 9263 41976 9680 42004
rect 9263 41973 9275 41976
rect 9217 41967 9275 41973
rect 9674 41964 9680 41976
rect 9732 41964 9738 42016
rect 10502 41964 10508 42016
rect 10560 42004 10566 42016
rect 10689 42007 10747 42013
rect 10689 42004 10701 42007
rect 10560 41976 10701 42004
rect 10560 41964 10566 41976
rect 10689 41973 10701 41976
rect 10735 41973 10747 42007
rect 10689 41967 10747 41973
rect 14458 41964 14464 42016
rect 14516 42004 14522 42016
rect 16393 42007 16451 42013
rect 16393 42004 16405 42007
rect 14516 41976 16405 42004
rect 14516 41964 14522 41976
rect 16393 41973 16405 41976
rect 16439 42004 16451 42007
rect 17328 42004 17356 42103
rect 19058 42100 19064 42112
rect 19116 42100 19122 42152
rect 19242 42100 19248 42152
rect 19300 42140 19306 42152
rect 20732 42149 20760 42180
rect 20990 42168 20996 42180
rect 21048 42168 21054 42220
rect 19613 42143 19671 42149
rect 19613 42140 19625 42143
rect 19300 42112 19625 42140
rect 19300 42100 19306 42112
rect 19613 42109 19625 42112
rect 19659 42109 19671 42143
rect 19613 42103 19671 42109
rect 20717 42143 20775 42149
rect 20717 42109 20729 42143
rect 20763 42109 20775 42143
rect 20717 42103 20775 42109
rect 20809 42143 20867 42149
rect 20809 42109 20821 42143
rect 20855 42140 20867 42143
rect 21266 42140 21272 42152
rect 20855 42112 21272 42140
rect 20855 42109 20867 42112
rect 20809 42103 20867 42109
rect 19702 42032 19708 42084
rect 19760 42072 19766 42084
rect 20824 42072 20852 42103
rect 21266 42100 21272 42112
rect 21324 42100 21330 42152
rect 22830 42100 22836 42152
rect 22888 42140 22894 42152
rect 23474 42140 23480 42152
rect 22888 42112 23480 42140
rect 22888 42100 22894 42112
rect 23474 42100 23480 42112
rect 23532 42100 23538 42152
rect 23753 42143 23811 42149
rect 23753 42109 23765 42143
rect 23799 42140 23811 42143
rect 25130 42140 25136 42152
rect 23799 42112 25136 42140
rect 23799 42109 23811 42112
rect 23753 42103 23811 42109
rect 25130 42100 25136 42112
rect 25188 42100 25194 42152
rect 19760 42044 20852 42072
rect 19760 42032 19766 42044
rect 16439 41976 17356 42004
rect 16439 41973 16451 41976
rect 16393 41967 16451 41973
rect 20254 41964 20260 42016
rect 20312 41964 20318 42016
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 5166 41760 5172 41812
rect 5224 41760 5230 41812
rect 7653 41803 7711 41809
rect 7653 41769 7665 41803
rect 7699 41800 7711 41803
rect 7742 41800 7748 41812
rect 7699 41772 7748 41800
rect 7699 41769 7711 41772
rect 7653 41763 7711 41769
rect 7742 41760 7748 41772
rect 7800 41760 7806 41812
rect 7834 41760 7840 41812
rect 7892 41800 7898 41812
rect 8110 41800 8116 41812
rect 7892 41772 8116 41800
rect 7892 41760 7898 41772
rect 8110 41760 8116 41772
rect 8168 41760 8174 41812
rect 10689 41803 10747 41809
rect 10689 41769 10701 41803
rect 10735 41800 10747 41803
rect 11054 41800 11060 41812
rect 10735 41772 11060 41800
rect 10735 41769 10747 41772
rect 10689 41763 10747 41769
rect 11054 41760 11060 41772
rect 11112 41760 11118 41812
rect 17313 41803 17371 41809
rect 17313 41769 17325 41803
rect 17359 41800 17371 41803
rect 22922 41800 22928 41812
rect 17359 41772 22928 41800
rect 17359 41769 17371 41772
rect 17313 41763 17371 41769
rect 8021 41735 8079 41741
rect 8021 41701 8033 41735
rect 8067 41732 8079 41735
rect 8294 41732 8300 41744
rect 8067 41704 8300 41732
rect 8067 41701 8079 41704
rect 8021 41695 8079 41701
rect 5905 41667 5963 41673
rect 5905 41633 5917 41667
rect 5951 41664 5963 41667
rect 6178 41664 6184 41676
rect 5951 41636 6184 41664
rect 5951 41633 5963 41636
rect 5905 41627 5963 41633
rect 6178 41624 6184 41636
rect 6236 41624 6242 41676
rect 8036 41596 8064 41695
rect 8294 41692 8300 41704
rect 8352 41732 8358 41744
rect 9122 41732 9128 41744
rect 8352 41704 9128 41732
rect 8352 41692 8358 41704
rect 9122 41692 9128 41704
rect 9180 41692 9186 41744
rect 15286 41692 15292 41744
rect 15344 41732 15350 41744
rect 16114 41732 16120 41744
rect 15344 41704 16120 41732
rect 15344 41692 15350 41704
rect 16114 41692 16120 41704
rect 16172 41732 16178 41744
rect 16172 41704 16804 41732
rect 16172 41692 16178 41704
rect 9214 41624 9220 41676
rect 9272 41664 9278 41676
rect 10045 41667 10103 41673
rect 10045 41664 10057 41667
rect 9272 41636 10057 41664
rect 9272 41624 9278 41636
rect 10045 41633 10057 41636
rect 10091 41664 10103 41667
rect 10594 41664 10600 41676
rect 10091 41636 10600 41664
rect 10091 41633 10103 41636
rect 10045 41627 10103 41633
rect 10594 41624 10600 41636
rect 10652 41624 10658 41676
rect 10778 41624 10784 41676
rect 10836 41664 10842 41676
rect 11241 41667 11299 41673
rect 11241 41664 11253 41667
rect 10836 41636 11253 41664
rect 10836 41624 10842 41636
rect 11241 41633 11253 41636
rect 11287 41633 11299 41667
rect 11241 41627 11299 41633
rect 12342 41624 12348 41676
rect 12400 41664 12406 41676
rect 12802 41664 12808 41676
rect 12400 41636 12808 41664
rect 12400 41624 12406 41636
rect 12802 41624 12808 41636
rect 12860 41624 12866 41676
rect 16574 41624 16580 41676
rect 16632 41664 16638 41676
rect 16776 41673 16804 41704
rect 16669 41667 16727 41673
rect 16669 41664 16681 41667
rect 16632 41636 16681 41664
rect 16632 41624 16638 41636
rect 16669 41633 16681 41636
rect 16715 41633 16727 41667
rect 16669 41627 16727 41633
rect 16761 41667 16819 41673
rect 16761 41633 16773 41667
rect 16807 41633 16819 41667
rect 16761 41627 16819 41633
rect 7314 41568 8064 41596
rect 9309 41599 9367 41605
rect 9309 41565 9321 41599
rect 9355 41596 9367 41599
rect 10502 41596 10508 41608
rect 9355 41568 10508 41596
rect 9355 41565 9367 41568
rect 9309 41559 9367 41565
rect 10502 41556 10508 41568
rect 10560 41596 10566 41608
rect 11977 41599 12035 41605
rect 11977 41596 11989 41599
rect 10560 41568 11989 41596
rect 10560 41556 10566 41568
rect 11977 41565 11989 41568
rect 12023 41596 12035 41599
rect 13173 41599 13231 41605
rect 13173 41596 13185 41599
rect 12023 41568 13185 41596
rect 12023 41565 12035 41568
rect 11977 41559 12035 41565
rect 13173 41565 13185 41568
rect 13219 41565 13231 41599
rect 13173 41559 13231 41565
rect 5077 41531 5135 41537
rect 5077 41497 5089 41531
rect 5123 41528 5135 41531
rect 6181 41531 6239 41537
rect 5123 41500 5672 41528
rect 5123 41497 5135 41500
rect 5077 41491 5135 41497
rect 5644 41469 5672 41500
rect 6181 41497 6193 41531
rect 6227 41497 6239 41531
rect 6181 41491 6239 41497
rect 11149 41531 11207 41537
rect 11149 41497 11161 41531
rect 11195 41528 11207 41531
rect 13998 41528 14004 41540
rect 11195 41500 14004 41528
rect 11195 41497 11207 41500
rect 11149 41491 11207 41497
rect 5629 41463 5687 41469
rect 5629 41429 5641 41463
rect 5675 41460 5687 41463
rect 5902 41460 5908 41472
rect 5675 41432 5908 41460
rect 5675 41429 5687 41432
rect 5629 41423 5687 41429
rect 5902 41420 5908 41432
rect 5960 41420 5966 41472
rect 6196 41460 6224 41491
rect 13998 41488 14004 41500
rect 14056 41488 14062 41540
rect 16577 41531 16635 41537
rect 16577 41497 16589 41531
rect 16623 41528 16635 41531
rect 17328 41528 17356 41763
rect 22922 41760 22928 41772
rect 22980 41760 22986 41812
rect 24210 41760 24216 41812
rect 24268 41800 24274 41812
rect 24581 41803 24639 41809
rect 24581 41800 24593 41803
rect 24268 41772 24593 41800
rect 24268 41760 24274 41772
rect 24581 41769 24593 41772
rect 24627 41769 24639 41803
rect 24581 41763 24639 41769
rect 17770 41692 17776 41744
rect 17828 41732 17834 41744
rect 17828 41704 18828 41732
rect 17828 41692 17834 41704
rect 18506 41624 18512 41676
rect 18564 41664 18570 41676
rect 18800 41673 18828 41704
rect 21174 41692 21180 41744
rect 21232 41692 21238 41744
rect 21637 41735 21695 41741
rect 21637 41701 21649 41735
rect 21683 41732 21695 41735
rect 22554 41732 22560 41744
rect 21683 41704 22560 41732
rect 21683 41701 21695 41704
rect 21637 41695 21695 41701
rect 22554 41692 22560 41704
rect 22612 41692 22618 41744
rect 22833 41735 22891 41741
rect 22833 41701 22845 41735
rect 22879 41732 22891 41735
rect 25038 41732 25044 41744
rect 22879 41704 25044 41732
rect 22879 41701 22891 41704
rect 22833 41695 22891 41701
rect 25038 41692 25044 41704
rect 25096 41692 25102 41744
rect 25133 41735 25191 41741
rect 25133 41701 25145 41735
rect 25179 41732 25191 41735
rect 25406 41732 25412 41744
rect 25179 41704 25412 41732
rect 25179 41701 25191 41704
rect 25133 41695 25191 41701
rect 25406 41692 25412 41704
rect 25464 41692 25470 41744
rect 18601 41667 18659 41673
rect 18601 41664 18613 41667
rect 18564 41636 18613 41664
rect 18564 41624 18570 41636
rect 18601 41633 18613 41636
rect 18647 41633 18659 41667
rect 18601 41627 18659 41633
rect 18785 41667 18843 41673
rect 18785 41633 18797 41667
rect 18831 41664 18843 41667
rect 18966 41664 18972 41676
rect 18831 41636 18972 41664
rect 18831 41633 18843 41636
rect 18785 41627 18843 41633
rect 18966 41624 18972 41636
rect 19024 41624 19030 41676
rect 19702 41664 19708 41676
rect 19168 41636 19708 41664
rect 19168 41596 19196 41636
rect 19702 41624 19708 41636
rect 19760 41624 19766 41676
rect 20898 41664 20904 41676
rect 20824 41636 20904 41664
rect 16623 41500 17356 41528
rect 18064 41568 19196 41596
rect 16623 41497 16635 41500
rect 16577 41491 16635 41497
rect 7742 41460 7748 41472
rect 6196 41432 7748 41460
rect 7742 41420 7748 41432
rect 7800 41420 7806 41472
rect 9674 41420 9680 41472
rect 9732 41460 9738 41472
rect 10778 41460 10784 41472
rect 9732 41432 10784 41460
rect 9732 41420 9738 41432
rect 10778 41420 10784 41432
rect 10836 41420 10842 41472
rect 11054 41420 11060 41472
rect 11112 41420 11118 41472
rect 12802 41420 12808 41472
rect 12860 41460 12866 41472
rect 13630 41460 13636 41472
rect 12860 41432 13636 41460
rect 12860 41420 12866 41432
rect 13630 41420 13636 41432
rect 13688 41420 13694 41472
rect 16206 41420 16212 41472
rect 16264 41420 16270 41472
rect 16482 41420 16488 41472
rect 16540 41460 16546 41472
rect 18064 41460 18092 41568
rect 19242 41556 19248 41608
rect 19300 41596 19306 41608
rect 19429 41599 19487 41605
rect 19429 41596 19441 41599
rect 19300 41568 19441 41596
rect 19300 41556 19306 41568
rect 19429 41565 19441 41568
rect 19475 41565 19487 41599
rect 20824 41582 20852 41636
rect 20898 41624 20904 41636
rect 20956 41624 20962 41676
rect 22281 41667 22339 41673
rect 22281 41633 22293 41667
rect 22327 41664 22339 41667
rect 22462 41664 22468 41676
rect 22327 41636 22468 41664
rect 22327 41633 22339 41636
rect 22281 41627 22339 41633
rect 22462 41624 22468 41636
rect 22520 41624 22526 41676
rect 22646 41624 22652 41676
rect 22704 41664 22710 41676
rect 23293 41667 23351 41673
rect 23293 41664 23305 41667
rect 22704 41636 23305 41664
rect 22704 41624 22710 41636
rect 23293 41633 23305 41636
rect 23339 41633 23351 41667
rect 23293 41627 23351 41633
rect 23385 41667 23443 41673
rect 23385 41633 23397 41667
rect 23431 41664 23443 41667
rect 23474 41664 23480 41676
rect 23431 41636 23480 41664
rect 23431 41633 23443 41636
rect 23385 41627 23443 41633
rect 23474 41624 23480 41636
rect 23532 41624 23538 41676
rect 24489 41599 24547 41605
rect 19429 41559 19487 41565
rect 24489 41565 24501 41599
rect 24535 41596 24547 41599
rect 25314 41596 25320 41608
rect 24535 41568 25320 41596
rect 24535 41565 24547 41568
rect 24489 41559 24547 41565
rect 25314 41556 25320 41568
rect 25372 41556 25378 41608
rect 18509 41531 18567 41537
rect 18509 41497 18521 41531
rect 18555 41528 18567 41531
rect 19150 41528 19156 41540
rect 18555 41500 19156 41528
rect 18555 41497 18567 41500
rect 18509 41491 18567 41497
rect 19150 41488 19156 41500
rect 19208 41488 19214 41540
rect 20990 41488 20996 41540
rect 21048 41528 21054 41540
rect 22097 41531 22155 41537
rect 22097 41528 22109 41531
rect 21048 41500 22109 41528
rect 21048 41488 21054 41500
rect 22097 41497 22109 41500
rect 22143 41497 22155 41531
rect 22097 41491 22155 41497
rect 22186 41488 22192 41540
rect 22244 41528 22250 41540
rect 23201 41531 23259 41537
rect 23201 41528 23213 41531
rect 22244 41500 23213 41528
rect 22244 41488 22250 41500
rect 23201 41497 23213 41500
rect 23247 41497 23259 41531
rect 23201 41491 23259 41497
rect 24213 41531 24271 41537
rect 24213 41497 24225 41531
rect 24259 41528 24271 41531
rect 24259 41500 25360 41528
rect 24259 41497 24271 41500
rect 24213 41491 24271 41497
rect 25332 41472 25360 41500
rect 16540 41432 18092 41460
rect 18141 41463 18199 41469
rect 16540 41420 16546 41432
rect 18141 41429 18153 41463
rect 18187 41460 18199 41463
rect 18414 41460 18420 41472
rect 18187 41432 18420 41460
rect 18187 41429 18199 41432
rect 18141 41423 18199 41429
rect 18414 41420 18420 41432
rect 18472 41420 18478 41472
rect 19978 41420 19984 41472
rect 20036 41460 20042 41472
rect 21634 41460 21640 41472
rect 20036 41432 21640 41460
rect 20036 41420 20042 41432
rect 21634 41420 21640 41432
rect 21692 41420 21698 41472
rect 22002 41420 22008 41472
rect 22060 41420 22066 41472
rect 24854 41420 24860 41472
rect 24912 41420 24918 41472
rect 25314 41420 25320 41472
rect 25372 41420 25378 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 1946 41216 1952 41268
rect 2004 41256 2010 41268
rect 3329 41259 3387 41265
rect 3329 41256 3341 41259
rect 2004 41228 3341 41256
rect 2004 41216 2010 41228
rect 3329 41225 3341 41228
rect 3375 41225 3387 41259
rect 3329 41219 3387 41225
rect 6178 41216 6184 41268
rect 6236 41256 6242 41268
rect 7834 41256 7840 41268
rect 6236 41228 7840 41256
rect 6236 41216 6242 41228
rect 7834 41216 7840 41228
rect 7892 41256 7898 41268
rect 8021 41259 8079 41265
rect 8021 41256 8033 41259
rect 7892 41228 8033 41256
rect 7892 41216 7898 41228
rect 8021 41225 8033 41228
rect 8067 41225 8079 41259
rect 9398 41256 9404 41268
rect 8021 41219 8079 41225
rect 8956 41228 9404 41256
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1765 41123 1823 41129
rect 1765 41120 1777 41123
rect 1360 41092 1777 41120
rect 1360 41080 1366 41092
rect 1765 41089 1777 41092
rect 1811 41120 1823 41123
rect 2041 41123 2099 41129
rect 2041 41120 2053 41123
rect 1811 41092 2053 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 2041 41089 2053 41092
rect 2087 41089 2099 41123
rect 2041 41083 2099 41089
rect 3237 41123 3295 41129
rect 3237 41089 3249 41123
rect 3283 41120 3295 41123
rect 3697 41123 3755 41129
rect 3697 41120 3709 41123
rect 3283 41092 3709 41120
rect 3283 41089 3295 41092
rect 3237 41083 3295 41089
rect 3697 41089 3709 41092
rect 3743 41120 3755 41123
rect 4614 41120 4620 41132
rect 3743 41092 4620 41120
rect 3743 41089 3755 41092
rect 3697 41083 3755 41089
rect 4614 41080 4620 41092
rect 4672 41080 4678 41132
rect 8956 41129 8984 41228
rect 9398 41216 9404 41228
rect 9456 41216 9462 41268
rect 10962 41216 10968 41268
rect 11020 41216 11026 41268
rect 11698 41216 11704 41268
rect 11756 41216 11762 41268
rect 15749 41259 15807 41265
rect 15749 41225 15761 41259
rect 15795 41256 15807 41259
rect 16114 41256 16120 41268
rect 15795 41228 16120 41256
rect 15795 41225 15807 41228
rect 15749 41219 15807 41225
rect 10980 41188 11008 41216
rect 15378 41188 15384 41200
rect 10442 41160 11008 41188
rect 15134 41160 15384 41188
rect 15378 41148 15384 41160
rect 15436 41188 15442 41200
rect 15764 41188 15792 41219
rect 16114 41216 16120 41228
rect 16172 41256 16178 41268
rect 18969 41259 19027 41265
rect 18969 41256 18981 41259
rect 16172 41228 18981 41256
rect 16172 41216 16178 41228
rect 15436 41160 15792 41188
rect 17512 41188 17540 41228
rect 18969 41225 18981 41228
rect 19015 41225 19027 41259
rect 18969 41219 19027 41225
rect 19886 41216 19892 41268
rect 19944 41216 19950 41268
rect 20162 41216 20168 41268
rect 20220 41256 20226 41268
rect 20438 41256 20444 41268
rect 20220 41228 20444 41256
rect 20220 41216 20226 41228
rect 20438 41216 20444 41228
rect 20496 41216 20502 41268
rect 20806 41216 20812 41268
rect 20864 41256 20870 41268
rect 20990 41256 20996 41268
rect 20864 41228 20996 41256
rect 20864 41216 20870 41228
rect 20990 41216 20996 41228
rect 21048 41216 21054 41268
rect 21085 41259 21143 41265
rect 21085 41225 21097 41259
rect 21131 41256 21143 41259
rect 21450 41256 21456 41268
rect 21131 41228 21456 41256
rect 21131 41225 21143 41228
rect 21085 41219 21143 41225
rect 21450 41216 21456 41228
rect 21508 41216 21514 41268
rect 22002 41216 22008 41268
rect 22060 41216 22066 41268
rect 23474 41216 23480 41268
rect 23532 41256 23538 41268
rect 24673 41259 24731 41265
rect 24673 41256 24685 41259
rect 23532 41228 24685 41256
rect 23532 41216 23538 41228
rect 24673 41225 24685 41228
rect 24719 41225 24731 41259
rect 24673 41219 24731 41225
rect 21266 41188 21272 41200
rect 17512 41160 17618 41188
rect 18984 41160 21272 41188
rect 15436 41148 15442 41160
rect 8941 41123 8999 41129
rect 8941 41089 8953 41123
rect 8987 41089 8999 41123
rect 8941 41083 8999 41089
rect 10502 41080 10508 41132
rect 10560 41120 10566 41132
rect 12069 41123 12127 41129
rect 12069 41120 12081 41123
rect 10560 41092 12081 41120
rect 10560 41080 10566 41092
rect 12069 41089 12081 41092
rect 12115 41089 12127 41123
rect 12069 41083 12127 41089
rect 12161 41123 12219 41129
rect 12161 41089 12173 41123
rect 12207 41120 12219 41123
rect 12342 41120 12348 41132
rect 12207 41092 12348 41120
rect 12207 41089 12219 41092
rect 12161 41083 12219 41089
rect 12342 41080 12348 41092
rect 12400 41080 12406 41132
rect 13630 41080 13636 41132
rect 13688 41080 13694 41132
rect 16666 41080 16672 41132
rect 16724 41120 16730 41132
rect 16853 41123 16911 41129
rect 16853 41120 16865 41123
rect 16724 41092 16865 41120
rect 16724 41080 16730 41092
rect 16853 41089 16865 41092
rect 16899 41089 16911 41123
rect 16853 41083 16911 41089
rect 9214 41012 9220 41064
rect 9272 41012 9278 41064
rect 12250 41012 12256 41064
rect 12308 41012 12314 41064
rect 13909 41055 13967 41061
rect 13909 41021 13921 41055
rect 13955 41052 13967 41055
rect 13998 41052 14004 41064
rect 13955 41024 14004 41052
rect 13955 41021 13967 41024
rect 13909 41015 13967 41021
rect 13998 41012 14004 41024
rect 14056 41052 14062 41064
rect 15286 41052 15292 41064
rect 14056 41024 15292 41052
rect 14056 41012 14062 41024
rect 15286 41012 15292 41024
rect 15344 41012 15350 41064
rect 16758 41012 16764 41064
rect 16816 41052 16822 41064
rect 17129 41055 17187 41061
rect 17129 41052 17141 41055
rect 16816 41024 17141 41052
rect 16816 41012 16822 41024
rect 17129 41021 17141 41024
rect 17175 41052 17187 41055
rect 18984 41052 19012 41160
rect 21266 41148 21272 41160
rect 21324 41148 21330 41200
rect 22278 41148 22284 41200
rect 22336 41188 22342 41200
rect 23198 41188 23204 41200
rect 22336 41160 23204 41188
rect 22336 41148 22342 41160
rect 23198 41148 23204 41160
rect 23256 41148 23262 41200
rect 24210 41148 24216 41200
rect 24268 41148 24274 41200
rect 19794 41080 19800 41132
rect 19852 41080 19858 41132
rect 19904 41092 20116 41120
rect 17175 41024 19012 41052
rect 17175 41021 17187 41024
rect 17129 41015 17187 41021
rect 19610 41012 19616 41064
rect 19668 41052 19674 41064
rect 19904 41052 19932 41092
rect 20088 41061 20116 41092
rect 25314 41080 25320 41132
rect 25372 41080 25378 41132
rect 19668 41024 19932 41052
rect 20073 41055 20131 41061
rect 19668 41012 19674 41024
rect 20073 41021 20085 41055
rect 20119 41021 20131 41055
rect 20073 41015 20131 41021
rect 20990 41012 20996 41064
rect 21048 41052 21054 41064
rect 21177 41055 21235 41061
rect 21177 41052 21189 41055
rect 21048 41024 21189 41052
rect 21048 41012 21054 41024
rect 21177 41021 21189 41024
rect 21223 41021 21235 41055
rect 21177 41015 21235 41021
rect 21266 41012 21272 41064
rect 21324 41012 21330 41064
rect 22462 41052 22468 41064
rect 22066 41024 22468 41052
rect 15381 40987 15439 40993
rect 15381 40953 15393 40987
rect 15427 40984 15439 40987
rect 15746 40984 15752 40996
rect 15427 40956 15752 40984
rect 15427 40953 15439 40956
rect 15381 40947 15439 40953
rect 15746 40944 15752 40956
rect 15804 40944 15810 40996
rect 18322 40944 18328 40996
rect 18380 40984 18386 40996
rect 18966 40984 18972 40996
rect 18380 40956 18972 40984
rect 18380 40944 18386 40956
rect 18966 40944 18972 40956
rect 19024 40984 19030 40996
rect 19978 40984 19984 40996
rect 19024 40956 19984 40984
rect 19024 40944 19030 40956
rect 19978 40944 19984 40956
rect 20036 40944 20042 40996
rect 22066 40984 22094 41024
rect 22462 41012 22468 41024
rect 22520 41012 22526 41064
rect 22830 41012 22836 41064
rect 22888 41052 22894 41064
rect 22925 41055 22983 41061
rect 22925 41052 22937 41055
rect 22888 41024 22937 41052
rect 22888 41012 22894 41024
rect 22925 41021 22937 41024
rect 22971 41021 22983 41055
rect 22925 41015 22983 41021
rect 23198 41012 23204 41064
rect 23256 41052 23262 41064
rect 24854 41052 24860 41064
rect 23256 41024 24860 41052
rect 23256 41012 23262 41024
rect 24854 41012 24860 41024
rect 24912 41012 24918 41064
rect 20088 40956 22094 40984
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 1670 40916 1676 40928
rect 1627 40888 1676 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 1670 40876 1676 40888
rect 1728 40876 1734 40928
rect 9950 40876 9956 40928
rect 10008 40916 10014 40928
rect 10686 40916 10692 40928
rect 10008 40888 10692 40916
rect 10008 40876 10014 40888
rect 10686 40876 10692 40888
rect 10744 40876 10750 40928
rect 18506 40876 18512 40928
rect 18564 40916 18570 40928
rect 18601 40919 18659 40925
rect 18601 40916 18613 40919
rect 18564 40888 18613 40916
rect 18564 40876 18570 40888
rect 18601 40885 18613 40888
rect 18647 40885 18659 40919
rect 18601 40879 18659 40885
rect 19150 40876 19156 40928
rect 19208 40876 19214 40928
rect 19426 40876 19432 40928
rect 19484 40876 19490 40928
rect 19518 40876 19524 40928
rect 19576 40916 19582 40928
rect 20088 40916 20116 40956
rect 19576 40888 20116 40916
rect 20717 40919 20775 40925
rect 19576 40876 19582 40888
rect 20717 40885 20729 40919
rect 20763 40916 20775 40919
rect 20806 40916 20812 40928
rect 20763 40888 20812 40916
rect 20763 40885 20775 40888
rect 20717 40879 20775 40885
rect 20806 40876 20812 40888
rect 20864 40876 20870 40928
rect 21450 40876 21456 40928
rect 21508 40916 21514 40928
rect 25133 40919 25191 40925
rect 25133 40916 25145 40919
rect 21508 40888 25145 40916
rect 21508 40876 21514 40888
rect 25133 40885 25145 40888
rect 25179 40885 25191 40919
rect 25133 40879 25191 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 8570 40672 8576 40724
rect 8628 40672 8634 40724
rect 8662 40672 8668 40724
rect 8720 40712 8726 40724
rect 8720 40684 10364 40712
rect 8720 40672 8726 40684
rect 9217 40647 9275 40653
rect 9217 40613 9229 40647
rect 9263 40644 9275 40647
rect 10226 40644 10232 40656
rect 9263 40616 10232 40644
rect 9263 40613 9275 40616
rect 9217 40607 9275 40613
rect 10226 40604 10232 40616
rect 10284 40604 10290 40656
rect 10336 40644 10364 40684
rect 10594 40672 10600 40724
rect 10652 40672 10658 40724
rect 11238 40672 11244 40724
rect 11296 40712 11302 40724
rect 11296 40684 12434 40712
rect 11296 40672 11302 40684
rect 11057 40647 11115 40653
rect 11057 40644 11069 40647
rect 10336 40616 11069 40644
rect 11057 40613 11069 40616
rect 11103 40644 11115 40647
rect 12406 40644 12434 40684
rect 13906 40672 13912 40724
rect 13964 40712 13970 40724
rect 14737 40715 14795 40721
rect 14737 40712 14749 40715
rect 13964 40684 14749 40712
rect 13964 40672 13970 40684
rect 14737 40681 14749 40684
rect 14783 40712 14795 40715
rect 16301 40715 16359 40721
rect 14783 40684 15884 40712
rect 14783 40681 14795 40684
rect 14737 40675 14795 40681
rect 14829 40647 14887 40653
rect 14829 40644 14841 40647
rect 11103 40616 11744 40644
rect 12406 40616 14841 40644
rect 11103 40613 11115 40616
rect 11057 40607 11115 40613
rect 6457 40579 6515 40585
rect 6457 40545 6469 40579
rect 6503 40576 6515 40579
rect 6546 40576 6552 40588
rect 6503 40548 6552 40576
rect 6503 40545 6515 40548
rect 6457 40539 6515 40545
rect 6546 40536 6552 40548
rect 6604 40576 6610 40588
rect 9861 40579 9919 40585
rect 6604 40548 8248 40576
rect 6604 40536 6610 40548
rect 6178 40468 6184 40520
rect 6236 40468 6242 40520
rect 8220 40508 8248 40548
rect 9861 40545 9873 40579
rect 9907 40576 9919 40579
rect 10318 40576 10324 40588
rect 9907 40548 10324 40576
rect 9907 40545 9919 40548
rect 9861 40539 9919 40545
rect 10318 40536 10324 40548
rect 10376 40536 10382 40588
rect 11716 40585 11744 40616
rect 14829 40613 14841 40616
rect 14875 40644 14887 40647
rect 14875 40616 15700 40644
rect 14875 40613 14887 40616
rect 14829 40607 14887 40613
rect 11517 40579 11575 40585
rect 11517 40545 11529 40579
rect 11563 40545 11575 40579
rect 11517 40539 11575 40545
rect 11701 40579 11759 40585
rect 11701 40545 11713 40579
rect 11747 40545 11759 40579
rect 11701 40539 11759 40545
rect 13265 40579 13323 40585
rect 13265 40545 13277 40579
rect 13311 40576 13323 40579
rect 13630 40576 13636 40588
rect 13311 40548 13636 40576
rect 13311 40545 13323 40548
rect 13265 40539 13323 40545
rect 11532 40508 11560 40539
rect 13630 40536 13636 40548
rect 13688 40536 13694 40588
rect 15672 40585 15700 40616
rect 15856 40588 15884 40684
rect 16301 40681 16313 40715
rect 16347 40712 16359 40715
rect 19518 40712 19524 40724
rect 16347 40684 19524 40712
rect 16347 40681 16359 40684
rect 16301 40675 16359 40681
rect 15657 40579 15715 40585
rect 15657 40545 15669 40579
rect 15703 40545 15715 40579
rect 15657 40539 15715 40545
rect 15838 40536 15844 40588
rect 15896 40536 15902 40588
rect 8220 40480 11560 40508
rect 12434 40468 12440 40520
rect 12492 40508 12498 40520
rect 12989 40511 13047 40517
rect 12989 40508 13001 40511
rect 12492 40480 13001 40508
rect 12492 40468 12498 40480
rect 12989 40477 13001 40480
rect 13035 40477 13047 40511
rect 12989 40471 13047 40477
rect 15565 40511 15623 40517
rect 15565 40477 15577 40511
rect 15611 40508 15623 40511
rect 16316 40508 16344 40675
rect 19518 40672 19524 40684
rect 19576 40672 19582 40724
rect 19610 40672 19616 40724
rect 19668 40672 19674 40724
rect 20901 40715 20959 40721
rect 20901 40681 20913 40715
rect 20947 40712 20959 40715
rect 21082 40712 21088 40724
rect 20947 40684 21088 40712
rect 20947 40681 20959 40684
rect 20901 40675 20959 40681
rect 21082 40672 21088 40684
rect 21140 40672 21146 40724
rect 21192 40684 21404 40712
rect 16942 40604 16948 40656
rect 17000 40644 17006 40656
rect 17000 40616 17264 40644
rect 17000 40604 17006 40616
rect 17034 40536 17040 40588
rect 17092 40576 17098 40588
rect 17236 40585 17264 40616
rect 17310 40604 17316 40656
rect 17368 40644 17374 40656
rect 19628 40644 19656 40672
rect 17368 40616 19656 40644
rect 17368 40604 17374 40616
rect 20162 40604 20168 40656
rect 20220 40644 20226 40656
rect 21192 40644 21220 40684
rect 20220 40616 21220 40644
rect 21376 40644 21404 40684
rect 22554 40672 22560 40724
rect 22612 40712 22618 40724
rect 23014 40712 23020 40724
rect 22612 40684 23020 40712
rect 22612 40672 22618 40684
rect 23014 40672 23020 40684
rect 23072 40672 23078 40724
rect 24029 40715 24087 40721
rect 24029 40681 24041 40715
rect 24075 40712 24087 40715
rect 24210 40712 24216 40724
rect 24075 40684 24216 40712
rect 24075 40681 24087 40684
rect 24029 40675 24087 40681
rect 24210 40672 24216 40684
rect 24268 40712 24274 40724
rect 24397 40715 24455 40721
rect 24397 40712 24409 40715
rect 24268 40684 24409 40712
rect 24268 40672 24274 40684
rect 24397 40681 24409 40684
rect 24443 40681 24455 40715
rect 24397 40675 24455 40681
rect 25133 40647 25191 40653
rect 25133 40644 25145 40647
rect 21376 40616 25145 40644
rect 20220 40604 20226 40616
rect 25133 40613 25145 40616
rect 25179 40613 25191 40647
rect 25133 40607 25191 40613
rect 17129 40579 17187 40585
rect 17129 40576 17141 40579
rect 17092 40548 17141 40576
rect 17092 40536 17098 40548
rect 17129 40545 17141 40548
rect 17175 40545 17187 40579
rect 17129 40539 17187 40545
rect 17221 40579 17279 40585
rect 17221 40545 17233 40579
rect 17267 40545 17279 40579
rect 17221 40539 17279 40545
rect 19610 40536 19616 40588
rect 19668 40576 19674 40588
rect 21453 40579 21511 40585
rect 21453 40576 21465 40579
rect 19668 40548 21465 40576
rect 19668 40536 19674 40548
rect 21453 40545 21465 40548
rect 21499 40545 21511 40579
rect 21453 40539 21511 40545
rect 15611 40480 16344 40508
rect 15611 40477 15623 40480
rect 15565 40471 15623 40477
rect 16574 40468 16580 40520
rect 16632 40508 16638 40520
rect 19150 40508 19156 40520
rect 16632 40480 19156 40508
rect 16632 40468 16638 40480
rect 19150 40468 19156 40480
rect 19208 40468 19214 40520
rect 21361 40511 21419 40517
rect 21361 40477 21373 40511
rect 21407 40477 21419 40511
rect 21468 40508 21496 40539
rect 22094 40536 22100 40588
rect 22152 40576 22158 40588
rect 22925 40579 22983 40585
rect 22925 40576 22937 40579
rect 22152 40548 22937 40576
rect 22152 40536 22158 40548
rect 22925 40545 22937 40548
rect 22971 40545 22983 40579
rect 22925 40539 22983 40545
rect 23109 40579 23167 40585
rect 23109 40545 23121 40579
rect 23155 40576 23167 40579
rect 23382 40576 23388 40588
rect 23155 40548 23388 40576
rect 23155 40545 23167 40548
rect 23109 40539 23167 40545
rect 23382 40536 23388 40548
rect 23440 40536 23446 40588
rect 22462 40508 22468 40520
rect 21468 40480 22468 40508
rect 21361 40471 21419 40477
rect 7682 40412 8340 40440
rect 8312 40384 8340 40412
rect 8570 40400 8576 40452
rect 8628 40440 8634 40452
rect 9585 40443 9643 40449
rect 9585 40440 9597 40443
rect 8628 40412 9597 40440
rect 8628 40400 8634 40412
rect 9585 40409 9597 40412
rect 9631 40440 9643 40443
rect 11238 40440 11244 40452
rect 9631 40412 11244 40440
rect 9631 40409 9643 40412
rect 9585 40403 9643 40409
rect 11238 40400 11244 40412
rect 11296 40400 11302 40452
rect 11333 40443 11391 40449
rect 11333 40409 11345 40443
rect 11379 40440 11391 40443
rect 11793 40443 11851 40449
rect 11793 40440 11805 40443
rect 11379 40412 11805 40440
rect 11379 40409 11391 40412
rect 11333 40403 11391 40409
rect 11793 40409 11805 40412
rect 11839 40440 11851 40443
rect 12250 40440 12256 40452
rect 11839 40412 12256 40440
rect 11839 40409 11851 40412
rect 11793 40403 11851 40409
rect 12250 40400 12256 40412
rect 12308 40400 12314 40452
rect 13081 40443 13139 40449
rect 13081 40409 13093 40443
rect 13127 40440 13139 40443
rect 13725 40443 13783 40449
rect 13725 40440 13737 40443
rect 13127 40412 13737 40440
rect 13127 40409 13139 40412
rect 13081 40403 13139 40409
rect 13725 40409 13737 40412
rect 13771 40440 13783 40443
rect 15930 40440 15936 40452
rect 13771 40412 15936 40440
rect 13771 40409 13783 40412
rect 13725 40403 13783 40409
rect 15930 40400 15936 40412
rect 15988 40400 15994 40452
rect 17494 40440 17500 40452
rect 16684 40412 17500 40440
rect 7282 40332 7288 40384
rect 7340 40372 7346 40384
rect 7742 40372 7748 40384
rect 7340 40344 7748 40372
rect 7340 40332 7346 40344
rect 7742 40332 7748 40344
rect 7800 40372 7806 40384
rect 7929 40375 7987 40381
rect 7929 40372 7941 40375
rect 7800 40344 7941 40372
rect 7800 40332 7806 40344
rect 7929 40341 7941 40344
rect 7975 40341 7987 40375
rect 7929 40335 7987 40341
rect 8294 40332 8300 40384
rect 8352 40332 8358 40384
rect 8757 40375 8815 40381
rect 8757 40341 8769 40375
rect 8803 40372 8815 40375
rect 9490 40372 9496 40384
rect 8803 40344 9496 40372
rect 8803 40341 8815 40344
rect 8757 40335 8815 40341
rect 9490 40332 9496 40344
rect 9548 40372 9554 40384
rect 9677 40375 9735 40381
rect 9677 40372 9689 40375
rect 9548 40344 9689 40372
rect 9548 40332 9554 40344
rect 9677 40341 9689 40344
rect 9723 40341 9735 40375
rect 9677 40335 9735 40341
rect 10318 40332 10324 40384
rect 10376 40332 10382 40384
rect 12158 40332 12164 40384
rect 12216 40332 12222 40384
rect 12618 40332 12624 40384
rect 12676 40332 12682 40384
rect 15197 40375 15255 40381
rect 15197 40341 15209 40375
rect 15243 40372 15255 40375
rect 15378 40372 15384 40384
rect 15243 40344 15384 40372
rect 15243 40341 15255 40344
rect 15197 40335 15255 40341
rect 15378 40332 15384 40344
rect 15436 40332 15442 40384
rect 16684 40381 16712 40412
rect 17494 40400 17500 40412
rect 17552 40400 17558 40452
rect 19168 40440 19196 40468
rect 21376 40440 21404 40471
rect 22462 40468 22468 40480
rect 22520 40468 22526 40520
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40508 22891 40511
rect 23014 40508 23020 40520
rect 22879 40480 23020 40508
rect 22879 40477 22891 40480
rect 22833 40471 22891 40477
rect 23014 40468 23020 40480
rect 23072 40468 23078 40520
rect 24673 40511 24731 40517
rect 24673 40477 24685 40511
rect 24719 40508 24731 40511
rect 25314 40508 25320 40520
rect 24719 40480 25320 40508
rect 24719 40477 24731 40480
rect 24673 40471 24731 40477
rect 25314 40468 25320 40480
rect 25372 40468 25378 40520
rect 21726 40440 21732 40452
rect 19168 40412 21732 40440
rect 21726 40400 21732 40412
rect 21784 40440 21790 40452
rect 21913 40443 21971 40449
rect 21913 40440 21925 40443
rect 21784 40412 21925 40440
rect 21784 40400 21790 40412
rect 21913 40409 21925 40412
rect 21959 40440 21971 40443
rect 22002 40440 22008 40452
rect 21959 40412 22008 40440
rect 21959 40409 21971 40412
rect 21913 40403 21971 40409
rect 22002 40400 22008 40412
rect 22060 40400 22066 40452
rect 22189 40443 22247 40449
rect 22189 40409 22201 40443
rect 22235 40440 22247 40443
rect 24213 40443 24271 40449
rect 22235 40412 22784 40440
rect 22235 40409 22247 40412
rect 22189 40403 22247 40409
rect 16669 40375 16727 40381
rect 16669 40341 16681 40375
rect 16715 40341 16727 40375
rect 16669 40335 16727 40341
rect 17034 40332 17040 40384
rect 17092 40332 17098 40384
rect 19794 40332 19800 40384
rect 19852 40372 19858 40384
rect 20349 40375 20407 40381
rect 20349 40372 20361 40375
rect 19852 40344 20361 40372
rect 19852 40332 19858 40344
rect 20349 40341 20361 40344
rect 20395 40372 20407 40375
rect 20438 40372 20444 40384
rect 20395 40344 20444 40372
rect 20395 40341 20407 40344
rect 20349 40335 20407 40341
rect 20438 40332 20444 40344
rect 20496 40332 20502 40384
rect 21266 40332 21272 40384
rect 21324 40372 21330 40384
rect 22204 40372 22232 40403
rect 21324 40344 22232 40372
rect 22465 40375 22523 40381
rect 21324 40332 21330 40344
rect 22465 40341 22477 40375
rect 22511 40372 22523 40375
rect 22646 40372 22652 40384
rect 22511 40344 22652 40372
rect 22511 40341 22523 40344
rect 22465 40335 22523 40341
rect 22646 40332 22652 40344
rect 22704 40332 22710 40384
rect 22756 40372 22784 40412
rect 24213 40409 24225 40443
rect 24259 40440 24271 40443
rect 24762 40440 24768 40452
rect 24259 40412 24768 40440
rect 24259 40409 24271 40412
rect 24213 40403 24271 40409
rect 24762 40400 24768 40412
rect 24820 40400 24826 40452
rect 24857 40443 24915 40449
rect 24857 40409 24869 40443
rect 24903 40440 24915 40443
rect 25222 40440 25228 40452
rect 24903 40412 25228 40440
rect 24903 40409 24915 40412
rect 24857 40403 24915 40409
rect 25222 40400 25228 40412
rect 25280 40400 25286 40452
rect 22922 40372 22928 40384
rect 22756 40344 22928 40372
rect 22922 40332 22928 40344
rect 22980 40372 22986 40384
rect 25774 40372 25780 40384
rect 22980 40344 25780 40372
rect 22980 40332 22986 40344
rect 25774 40332 25780 40344
rect 25832 40332 25838 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 7285 40171 7343 40177
rect 7285 40137 7297 40171
rect 7331 40168 7343 40171
rect 7374 40168 7380 40180
rect 7331 40140 7380 40168
rect 7331 40137 7343 40140
rect 7285 40131 7343 40137
rect 7374 40128 7380 40140
rect 7432 40128 7438 40180
rect 8754 40128 8760 40180
rect 8812 40168 8818 40180
rect 10318 40168 10324 40180
rect 8812 40140 10324 40168
rect 8812 40128 8818 40140
rect 10318 40128 10324 40140
rect 10376 40168 10382 40180
rect 10376 40140 10548 40168
rect 10376 40128 10382 40140
rect 7653 40103 7711 40109
rect 7653 40100 7665 40103
rect 7392 40072 7665 40100
rect 7392 40044 7420 40072
rect 7653 40069 7665 40072
rect 7699 40069 7711 40103
rect 7653 40063 7711 40069
rect 7834 40060 7840 40112
rect 7892 40060 7898 40112
rect 7926 40060 7932 40112
rect 7984 40100 7990 40112
rect 8294 40100 8300 40112
rect 7984 40072 8300 40100
rect 7984 40060 7990 40072
rect 8294 40060 8300 40072
rect 8352 40100 8358 40112
rect 10520 40109 10548 40140
rect 10962 40128 10968 40180
rect 11020 40168 11026 40180
rect 11517 40171 11575 40177
rect 11517 40168 11529 40171
rect 11020 40140 11529 40168
rect 11020 40128 11026 40140
rect 11517 40137 11529 40140
rect 11563 40168 11575 40171
rect 11698 40168 11704 40180
rect 11563 40140 11704 40168
rect 11563 40137 11575 40140
rect 11517 40131 11575 40137
rect 11698 40128 11704 40140
rect 11756 40128 11762 40180
rect 12250 40128 12256 40180
rect 12308 40168 12314 40180
rect 12308 40140 15516 40168
rect 12308 40128 12314 40140
rect 10505 40103 10563 40109
rect 8352 40072 9246 40100
rect 8352 40060 8358 40072
rect 10505 40069 10517 40103
rect 10551 40069 10563 40103
rect 14550 40100 14556 40112
rect 14398 40072 14556 40100
rect 10505 40063 10563 40069
rect 14550 40060 14556 40072
rect 14608 40100 14614 40112
rect 15013 40103 15071 40109
rect 15013 40100 15025 40103
rect 14608 40072 15025 40100
rect 14608 40060 14614 40072
rect 15013 40069 15025 40072
rect 15059 40100 15071 40103
rect 15286 40100 15292 40112
rect 15059 40072 15292 40100
rect 15059 40069 15071 40072
rect 15013 40063 15071 40069
rect 15286 40060 15292 40072
rect 15344 40060 15350 40112
rect 15488 40100 15516 40140
rect 15562 40128 15568 40180
rect 15620 40128 15626 40180
rect 15856 40140 18184 40168
rect 15856 40100 15884 40140
rect 15488 40072 15884 40100
rect 15933 40103 15991 40109
rect 15933 40069 15945 40103
rect 15979 40100 15991 40103
rect 16298 40100 16304 40112
rect 15979 40072 16304 40100
rect 15979 40069 15991 40072
rect 15933 40063 15991 40069
rect 16298 40060 16304 40072
rect 16356 40060 16362 40112
rect 18156 40100 18184 40140
rect 18230 40128 18236 40180
rect 18288 40128 18294 40180
rect 18414 40128 18420 40180
rect 18472 40168 18478 40180
rect 18693 40171 18751 40177
rect 18693 40168 18705 40171
rect 18472 40140 18705 40168
rect 18472 40128 18478 40140
rect 18693 40137 18705 40140
rect 18739 40137 18751 40171
rect 18693 40131 18751 40137
rect 19797 40171 19855 40177
rect 19797 40137 19809 40171
rect 19843 40168 19855 40171
rect 20622 40168 20628 40180
rect 19843 40140 20628 40168
rect 19843 40137 19855 40140
rect 19797 40131 19855 40137
rect 20622 40128 20628 40140
rect 20680 40128 20686 40180
rect 22462 40128 22468 40180
rect 22520 40168 22526 40180
rect 23290 40168 23296 40180
rect 22520 40140 23296 40168
rect 22520 40128 22526 40140
rect 23290 40128 23296 40140
rect 23348 40168 23354 40180
rect 25225 40171 25283 40177
rect 25225 40168 25237 40171
rect 23348 40140 25237 40168
rect 23348 40128 23354 40140
rect 25225 40137 25237 40140
rect 25271 40137 25283 40171
rect 25225 40131 25283 40137
rect 18322 40100 18328 40112
rect 18156 40072 18328 40100
rect 18322 40060 18328 40072
rect 18380 40060 18386 40112
rect 18601 40103 18659 40109
rect 18601 40100 18613 40103
rect 18432 40072 18613 40100
rect 7374 39992 7380 40044
rect 7432 39992 7438 40044
rect 7852 40032 7880 40060
rect 18432 40044 18460 40072
rect 18601 40069 18613 40072
rect 18647 40069 18659 40103
rect 18601 40063 18659 40069
rect 20165 40103 20223 40109
rect 20165 40069 20177 40103
rect 20211 40069 20223 40103
rect 20165 40063 20223 40069
rect 8481 40035 8539 40041
rect 8481 40032 8493 40035
rect 7852 40004 8493 40032
rect 8481 40001 8493 40004
rect 8527 40001 8539 40035
rect 8481 39995 8539 40001
rect 12802 39992 12808 40044
rect 12860 40032 12866 40044
rect 12897 40035 12955 40041
rect 12897 40032 12909 40035
rect 12860 40004 12909 40032
rect 12860 39992 12866 40004
rect 12897 40001 12909 40004
rect 12943 40001 12955 40035
rect 12897 39995 12955 40001
rect 18414 39992 18420 40044
rect 18472 39992 18478 40044
rect 19978 40032 19984 40044
rect 18892 40004 19984 40032
rect 7742 39924 7748 39976
rect 7800 39924 7806 39976
rect 7834 39924 7840 39976
rect 7892 39924 7898 39976
rect 8757 39967 8815 39973
rect 8757 39933 8769 39967
rect 8803 39964 8815 39967
rect 9950 39964 9956 39976
rect 8803 39936 9956 39964
rect 8803 39933 8815 39936
rect 8757 39927 8815 39933
rect 9950 39924 9956 39936
rect 10008 39924 10014 39976
rect 10962 39924 10968 39976
rect 11020 39924 11026 39976
rect 13173 39967 13231 39973
rect 13173 39933 13185 39967
rect 13219 39964 13231 39967
rect 15746 39964 15752 39976
rect 13219 39936 15752 39964
rect 13219 39933 13231 39936
rect 13173 39927 13231 39933
rect 15746 39924 15752 39936
rect 15804 39924 15810 39976
rect 16022 39924 16028 39976
rect 16080 39924 16086 39976
rect 16114 39924 16120 39976
rect 16172 39924 16178 39976
rect 18782 39924 18788 39976
rect 18840 39924 18846 39976
rect 10042 39856 10048 39908
rect 10100 39896 10106 39908
rect 12710 39896 12716 39908
rect 10100 39868 12716 39896
rect 10100 39856 10106 39868
rect 12710 39856 12716 39868
rect 12768 39856 12774 39908
rect 17126 39856 17132 39908
rect 17184 39896 17190 39908
rect 18892 39896 18920 40004
rect 19978 39992 19984 40004
rect 20036 40032 20042 40044
rect 20180 40032 20208 40063
rect 20438 40060 20444 40112
rect 20496 40100 20502 40112
rect 20496 40072 22416 40100
rect 20496 40060 20502 40072
rect 20809 40035 20867 40041
rect 20809 40032 20821 40035
rect 20036 40004 20208 40032
rect 20272 40004 20821 40032
rect 20036 39992 20042 40004
rect 19334 39924 19340 39976
rect 19392 39964 19398 39976
rect 19702 39964 19708 39976
rect 19392 39936 19708 39964
rect 19392 39924 19398 39936
rect 19702 39924 19708 39936
rect 19760 39964 19766 39976
rect 20272 39973 20300 40004
rect 20809 40001 20821 40004
rect 20855 40001 20867 40035
rect 20809 39995 20867 40001
rect 20257 39967 20315 39973
rect 20257 39964 20269 39967
rect 19760 39936 20269 39964
rect 19760 39924 19766 39936
rect 20257 39933 20269 39936
rect 20303 39933 20315 39967
rect 20257 39927 20315 39933
rect 20346 39924 20352 39976
rect 20404 39924 20410 39976
rect 20824 39964 20852 39995
rect 21726 39992 21732 40044
rect 21784 40032 21790 40044
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 21784 40004 22293 40032
rect 21784 39992 21790 40004
rect 22281 40001 22293 40004
rect 22327 40001 22339 40035
rect 22281 39995 22339 40001
rect 22388 39964 22416 40072
rect 22830 40060 22836 40112
rect 22888 40100 22894 40112
rect 22888 40072 23428 40100
rect 22888 40060 22894 40072
rect 22557 40035 22615 40041
rect 22557 40001 22569 40035
rect 22603 40032 22615 40035
rect 22922 40032 22928 40044
rect 22603 40004 22928 40032
rect 22603 40001 22615 40004
rect 22557 39995 22615 40001
rect 22922 39992 22928 40004
rect 22980 39992 22986 40044
rect 23400 40032 23428 40072
rect 24210 40060 24216 40112
rect 24268 40060 24274 40112
rect 23477 40035 23535 40041
rect 23477 40032 23489 40035
rect 23400 40004 23489 40032
rect 23477 40001 23489 40004
rect 23523 40001 23535 40035
rect 23477 39995 23535 40001
rect 23382 39964 23388 39976
rect 20824 39936 22094 39964
rect 22388 39936 23388 39964
rect 17184 39868 18920 39896
rect 17184 39856 17190 39868
rect 19058 39856 19064 39908
rect 19116 39896 19122 39908
rect 22066 39896 22094 39936
rect 23382 39924 23388 39936
rect 23440 39924 23446 39976
rect 23753 39967 23811 39973
rect 23753 39933 23765 39967
rect 23799 39964 23811 39967
rect 24486 39964 24492 39976
rect 23799 39936 24492 39964
rect 23799 39933 23811 39936
rect 23753 39927 23811 39933
rect 24486 39924 24492 39936
rect 24544 39924 24550 39976
rect 22830 39896 22836 39908
rect 19116 39868 21128 39896
rect 22066 39868 22836 39896
rect 19116 39856 19122 39868
rect 7098 39788 7104 39840
rect 7156 39828 7162 39840
rect 10686 39828 10692 39840
rect 7156 39800 10692 39828
rect 7156 39788 7162 39800
rect 10686 39788 10692 39800
rect 10744 39788 10750 39840
rect 14642 39788 14648 39840
rect 14700 39788 14706 39840
rect 16298 39788 16304 39840
rect 16356 39828 16362 39840
rect 16669 39831 16727 39837
rect 16669 39828 16681 39831
rect 16356 39800 16681 39828
rect 16356 39788 16362 39800
rect 16669 39797 16681 39800
rect 16715 39797 16727 39831
rect 16669 39791 16727 39797
rect 19978 39788 19984 39840
rect 20036 39828 20042 39840
rect 20622 39828 20628 39840
rect 20036 39800 20628 39828
rect 20036 39788 20042 39800
rect 20622 39788 20628 39800
rect 20680 39828 20686 39840
rect 20993 39831 21051 39837
rect 20993 39828 21005 39831
rect 20680 39800 21005 39828
rect 20680 39788 20686 39800
rect 20993 39797 21005 39800
rect 21039 39797 21051 39831
rect 21100 39828 21128 39868
rect 22830 39856 22836 39868
rect 22888 39856 22894 39908
rect 25590 39828 25596 39840
rect 21100 39800 25596 39828
rect 20993 39791 21051 39797
rect 25590 39788 25596 39800
rect 25648 39788 25654 39840
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 6546 39584 6552 39636
rect 6604 39624 6610 39636
rect 6641 39627 6699 39633
rect 6641 39624 6653 39627
rect 6604 39596 6653 39624
rect 6604 39584 6610 39596
rect 6641 39593 6653 39596
rect 6687 39593 6699 39627
rect 6641 39587 6699 39593
rect 7742 39584 7748 39636
rect 7800 39624 7806 39636
rect 9769 39627 9827 39633
rect 9769 39624 9781 39627
rect 7800 39596 9781 39624
rect 7800 39584 7806 39596
rect 9769 39593 9781 39596
rect 9815 39593 9827 39627
rect 9769 39587 9827 39593
rect 10778 39584 10784 39636
rect 10836 39624 10842 39636
rect 16114 39624 16120 39636
rect 10836 39596 16120 39624
rect 10836 39584 10842 39596
rect 16114 39584 16120 39596
rect 16172 39584 16178 39636
rect 18598 39584 18604 39636
rect 18656 39624 18662 39636
rect 18785 39627 18843 39633
rect 18785 39624 18797 39627
rect 18656 39596 18797 39624
rect 18656 39584 18662 39596
rect 18785 39593 18797 39596
rect 18831 39593 18843 39627
rect 18785 39587 18843 39593
rect 19058 39584 19064 39636
rect 19116 39584 19122 39636
rect 21269 39627 21327 39633
rect 21269 39593 21281 39627
rect 21315 39624 21327 39627
rect 22186 39624 22192 39636
rect 21315 39596 22192 39624
rect 21315 39593 21327 39596
rect 21269 39587 21327 39593
rect 22186 39584 22192 39596
rect 22244 39584 22250 39636
rect 25406 39624 25412 39636
rect 22296 39596 25412 39624
rect 12710 39516 12716 39568
rect 12768 39556 12774 39568
rect 15565 39559 15623 39565
rect 15565 39556 15577 39559
rect 12768 39528 15577 39556
rect 12768 39516 12774 39528
rect 15565 39525 15577 39528
rect 15611 39525 15623 39559
rect 15565 39519 15623 39525
rect 16022 39516 16028 39568
rect 16080 39556 16086 39568
rect 22296 39556 22324 39596
rect 25406 39584 25412 39596
rect 25464 39584 25470 39636
rect 16080 39528 22324 39556
rect 22649 39559 22707 39565
rect 16080 39516 16086 39528
rect 22649 39525 22661 39559
rect 22695 39556 22707 39559
rect 22695 39528 24992 39556
rect 22695 39525 22707 39528
rect 22649 39519 22707 39525
rect 4893 39491 4951 39497
rect 4893 39457 4905 39491
rect 4939 39488 4951 39491
rect 6178 39488 6184 39500
rect 4939 39460 6184 39488
rect 4939 39457 4951 39460
rect 4893 39451 4951 39457
rect 6178 39448 6184 39460
rect 6236 39488 6242 39500
rect 7101 39491 7159 39497
rect 7101 39488 7113 39491
rect 6236 39460 7113 39488
rect 6236 39448 6242 39460
rect 7101 39457 7113 39460
rect 7147 39457 7159 39491
rect 7101 39451 7159 39457
rect 10226 39448 10232 39500
rect 10284 39448 10290 39500
rect 10321 39491 10379 39497
rect 10321 39457 10333 39491
rect 10367 39457 10379 39491
rect 10321 39451 10379 39457
rect 10965 39491 11023 39497
rect 10965 39457 10977 39491
rect 11011 39488 11023 39491
rect 12434 39488 12440 39500
rect 11011 39460 12440 39488
rect 11011 39457 11023 39460
rect 10965 39451 11023 39457
rect 8570 39380 8576 39432
rect 8628 39420 8634 39432
rect 10336 39420 10364 39451
rect 12434 39448 12440 39460
rect 12492 39488 12498 39500
rect 12802 39488 12808 39500
rect 12492 39460 12808 39488
rect 12492 39448 12498 39460
rect 12802 39448 12808 39460
rect 12860 39448 12866 39500
rect 13814 39448 13820 39500
rect 13872 39488 13878 39500
rect 13909 39491 13967 39497
rect 13909 39488 13921 39491
rect 13872 39460 13921 39488
rect 13872 39448 13878 39460
rect 13909 39457 13921 39460
rect 13955 39488 13967 39491
rect 14829 39491 14887 39497
rect 14829 39488 14841 39491
rect 13955 39460 14841 39488
rect 13955 39457 13967 39460
rect 13909 39451 13967 39457
rect 14829 39457 14841 39460
rect 14875 39457 14887 39491
rect 14829 39451 14887 39457
rect 15013 39491 15071 39497
rect 15013 39457 15025 39491
rect 15059 39488 15071 39491
rect 15654 39488 15660 39500
rect 15059 39460 15660 39488
rect 15059 39457 15071 39460
rect 15013 39451 15071 39457
rect 15654 39448 15660 39460
rect 15712 39448 15718 39500
rect 16209 39491 16267 39497
rect 16209 39457 16221 39491
rect 16255 39488 16267 39491
rect 17678 39488 17684 39500
rect 16255 39460 17684 39488
rect 16255 39457 16267 39460
rect 16209 39451 16267 39457
rect 17678 39448 17684 39460
rect 17736 39448 17742 39500
rect 19426 39448 19432 39500
rect 19484 39488 19490 39500
rect 19889 39491 19947 39497
rect 19889 39488 19901 39491
rect 19484 39460 19901 39488
rect 19484 39448 19490 39460
rect 19889 39457 19901 39460
rect 19935 39457 19947 39491
rect 19889 39451 19947 39457
rect 20070 39448 20076 39500
rect 20128 39448 20134 39500
rect 21726 39448 21732 39500
rect 21784 39448 21790 39500
rect 21913 39491 21971 39497
rect 21913 39457 21925 39491
rect 21959 39457 21971 39491
rect 21913 39451 21971 39457
rect 23293 39491 23351 39497
rect 23293 39457 23305 39491
rect 23339 39488 23351 39491
rect 23474 39488 23480 39500
rect 23339 39460 23480 39488
rect 23339 39457 23351 39460
rect 23293 39451 23351 39457
rect 12894 39420 12900 39432
rect 8628 39392 10364 39420
rect 12374 39392 12900 39420
rect 8628 39380 8634 39392
rect 12894 39380 12900 39392
rect 12952 39420 12958 39432
rect 13081 39423 13139 39429
rect 13081 39420 13093 39423
rect 12952 39392 13093 39420
rect 12952 39380 12958 39392
rect 13081 39389 13093 39392
rect 13127 39420 13139 39423
rect 14274 39420 14280 39432
rect 13127 39392 14280 39420
rect 13127 39389 13139 39392
rect 13081 39383 13139 39389
rect 14274 39380 14280 39392
rect 14332 39420 14338 39432
rect 14550 39420 14556 39432
rect 14332 39392 14556 39420
rect 14332 39380 14338 39392
rect 14550 39380 14556 39392
rect 14608 39380 14614 39432
rect 21266 39420 21272 39432
rect 17972 39392 21272 39420
rect 5169 39355 5227 39361
rect 5169 39321 5181 39355
rect 5215 39321 5227 39355
rect 7926 39352 7932 39364
rect 6394 39324 7932 39352
rect 5169 39315 5227 39321
rect 5184 39284 5212 39315
rect 7024 39296 7052 39324
rect 7926 39312 7932 39324
rect 7984 39312 7990 39364
rect 11238 39312 11244 39364
rect 11296 39312 11302 39364
rect 14737 39355 14795 39361
rect 14737 39321 14749 39355
rect 14783 39352 14795 39355
rect 15010 39352 15016 39364
rect 14783 39324 15016 39352
rect 14783 39321 14795 39324
rect 14737 39315 14795 39321
rect 15010 39312 15016 39324
rect 15068 39312 15074 39364
rect 17034 39352 17040 39364
rect 15120 39324 17040 39352
rect 5810 39284 5816 39296
rect 5184 39256 5816 39284
rect 5810 39244 5816 39256
rect 5868 39244 5874 39296
rect 7006 39244 7012 39296
rect 7064 39244 7070 39296
rect 8294 39244 8300 39296
rect 8352 39284 8358 39296
rect 9125 39287 9183 39293
rect 9125 39284 9137 39287
rect 8352 39256 9137 39284
rect 8352 39244 8358 39256
rect 9125 39253 9137 39256
rect 9171 39253 9183 39287
rect 9125 39247 9183 39253
rect 10134 39244 10140 39296
rect 10192 39244 10198 39296
rect 12710 39244 12716 39296
rect 12768 39244 12774 39296
rect 13078 39244 13084 39296
rect 13136 39284 13142 39296
rect 13265 39287 13323 39293
rect 13265 39284 13277 39287
rect 13136 39256 13277 39284
rect 13136 39244 13142 39256
rect 13265 39253 13277 39256
rect 13311 39284 13323 39287
rect 13906 39284 13912 39296
rect 13311 39256 13912 39284
rect 13311 39253 13323 39256
rect 13265 39247 13323 39253
rect 13906 39244 13912 39256
rect 13964 39244 13970 39296
rect 14369 39287 14427 39293
rect 14369 39253 14381 39287
rect 14415 39284 14427 39287
rect 15120 39284 15148 39324
rect 17034 39312 17040 39324
rect 17092 39312 17098 39364
rect 17218 39312 17224 39364
rect 17276 39352 17282 39364
rect 17972 39352 18000 39392
rect 21266 39380 21272 39392
rect 21324 39420 21330 39432
rect 21637 39423 21695 39429
rect 21637 39420 21649 39423
rect 21324 39392 21649 39420
rect 21324 39380 21330 39392
rect 21637 39389 21649 39392
rect 21683 39389 21695 39423
rect 21637 39383 21695 39389
rect 17276 39324 18000 39352
rect 17276 39312 17282 39324
rect 18782 39312 18788 39364
rect 18840 39352 18846 39364
rect 19797 39355 19855 39361
rect 19797 39352 19809 39355
rect 18840 39324 19809 39352
rect 18840 39312 18846 39324
rect 19797 39321 19809 39324
rect 19843 39321 19855 39355
rect 19797 39315 19855 39321
rect 14415 39256 15148 39284
rect 14415 39253 14427 39256
rect 14369 39247 14427 39253
rect 15470 39244 15476 39296
rect 15528 39284 15534 39296
rect 15933 39287 15991 39293
rect 15933 39284 15945 39287
rect 15528 39256 15945 39284
rect 15528 39244 15534 39256
rect 15933 39253 15945 39256
rect 15979 39253 15991 39287
rect 15933 39247 15991 39253
rect 16022 39244 16028 39296
rect 16080 39244 16086 39296
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 18601 39287 18659 39293
rect 18601 39284 18613 39287
rect 18472 39256 18613 39284
rect 18472 39244 18478 39256
rect 18601 39253 18613 39256
rect 18647 39284 18659 39287
rect 18690 39284 18696 39296
rect 18647 39256 18696 39284
rect 18647 39253 18659 39256
rect 18601 39247 18659 39253
rect 18690 39244 18696 39256
rect 18748 39244 18754 39296
rect 19429 39287 19487 39293
rect 19429 39253 19441 39287
rect 19475 39284 19487 39287
rect 20346 39284 20352 39296
rect 19475 39256 20352 39284
rect 19475 39253 19487 39256
rect 19429 39247 19487 39253
rect 20346 39244 20352 39256
rect 20404 39244 20410 39296
rect 20438 39244 20444 39296
rect 20496 39244 20502 39296
rect 20622 39244 20628 39296
rect 20680 39284 20686 39296
rect 21082 39284 21088 39296
rect 20680 39256 21088 39284
rect 20680 39244 20686 39256
rect 21082 39244 21088 39256
rect 21140 39244 21146 39296
rect 21818 39244 21824 39296
rect 21876 39284 21882 39296
rect 21928 39284 21956 39451
rect 23474 39448 23480 39460
rect 23532 39448 23538 39500
rect 22002 39380 22008 39432
rect 22060 39420 22066 39432
rect 24964 39429 24992 39528
rect 25038 39448 25044 39500
rect 25096 39448 25102 39500
rect 25130 39448 25136 39500
rect 25188 39448 25194 39500
rect 23109 39423 23167 39429
rect 23109 39420 23121 39423
rect 22060 39392 23121 39420
rect 22060 39380 22066 39392
rect 23109 39389 23121 39392
rect 23155 39389 23167 39423
rect 23109 39383 23167 39389
rect 24949 39423 25007 39429
rect 24949 39389 24961 39423
rect 24995 39389 25007 39423
rect 24949 39383 25007 39389
rect 23017 39355 23075 39361
rect 23017 39321 23029 39355
rect 23063 39352 23075 39355
rect 23845 39355 23903 39361
rect 23845 39352 23857 39355
rect 23063 39324 23857 39352
rect 23063 39321 23075 39324
rect 23017 39315 23075 39321
rect 23845 39321 23857 39324
rect 23891 39321 23903 39355
rect 23845 39315 23903 39321
rect 22278 39284 22284 39296
rect 21876 39256 22284 39284
rect 21876 39244 21882 39256
rect 22278 39244 22284 39256
rect 22336 39244 22342 39296
rect 24302 39244 24308 39296
rect 24360 39284 24366 39296
rect 24581 39287 24639 39293
rect 24581 39284 24593 39287
rect 24360 39256 24593 39284
rect 24360 39244 24366 39256
rect 24581 39253 24593 39256
rect 24627 39253 24639 39287
rect 24581 39247 24639 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 8205 39083 8263 39089
rect 8205 39049 8217 39083
rect 8251 39080 8263 39083
rect 8662 39080 8668 39092
rect 8251 39052 8668 39080
rect 8251 39049 8263 39052
rect 8205 39043 8263 39049
rect 8662 39040 8668 39052
rect 8720 39080 8726 39092
rect 9493 39083 9551 39089
rect 9493 39080 9505 39083
rect 8720 39052 9505 39080
rect 8720 39040 8726 39052
rect 9493 39049 9505 39052
rect 9539 39049 9551 39083
rect 9493 39043 9551 39049
rect 10781 39083 10839 39089
rect 10781 39049 10793 39083
rect 10827 39080 10839 39083
rect 10962 39080 10968 39092
rect 10827 39052 10968 39080
rect 10827 39049 10839 39052
rect 10781 39043 10839 39049
rect 10962 39040 10968 39052
rect 11020 39040 11026 39092
rect 12250 39080 12256 39092
rect 11992 39052 12256 39080
rect 4062 38972 4068 39024
rect 4120 39012 4126 39024
rect 8297 39015 8355 39021
rect 8297 39012 8309 39015
rect 4120 38984 8309 39012
rect 4120 38972 4126 38984
rect 8297 38981 8309 38984
rect 8343 39012 8355 39015
rect 9585 39015 9643 39021
rect 9585 39012 9597 39015
rect 8343 38984 9597 39012
rect 8343 38981 8355 38984
rect 8297 38975 8355 38981
rect 9585 38981 9597 38984
rect 9631 39012 9643 39015
rect 11992 39012 12020 39052
rect 12250 39040 12256 39052
rect 12308 39040 12314 39092
rect 12986 39040 12992 39092
rect 13044 39080 13050 39092
rect 14277 39083 14335 39089
rect 13044 39052 13676 39080
rect 13044 39040 13050 39052
rect 12434 39012 12440 39024
rect 9631 38984 12020 39012
rect 12084 38984 12440 39012
rect 9631 38981 9643 38984
rect 9585 38975 9643 38981
rect 8386 38904 8392 38956
rect 8444 38944 8450 38956
rect 8662 38944 8668 38956
rect 8444 38916 8668 38944
rect 8444 38904 8450 38916
rect 8662 38904 8668 38916
rect 8720 38904 8726 38956
rect 8772 38916 10088 38944
rect 6730 38836 6736 38888
rect 6788 38876 6794 38888
rect 8478 38876 8484 38888
rect 6788 38848 8484 38876
rect 6788 38836 6794 38848
rect 8478 38836 8484 38848
rect 8536 38876 8542 38888
rect 8772 38876 8800 38916
rect 9582 38876 9588 38888
rect 8536 38848 8800 38876
rect 8864 38848 9588 38876
rect 8536 38836 8542 38848
rect 8665 38811 8723 38817
rect 8665 38808 8677 38811
rect 7760 38780 8677 38808
rect 7760 38752 7788 38780
rect 8665 38777 8677 38780
rect 8711 38777 8723 38811
rect 8665 38771 8723 38777
rect 7006 38700 7012 38752
rect 7064 38740 7070 38752
rect 7377 38743 7435 38749
rect 7377 38740 7389 38743
rect 7064 38712 7389 38740
rect 7064 38700 7070 38712
rect 7377 38709 7389 38712
rect 7423 38740 7435 38743
rect 7742 38740 7748 38752
rect 7423 38712 7748 38740
rect 7423 38709 7435 38712
rect 7377 38703 7435 38709
rect 7742 38700 7748 38712
rect 7800 38700 7806 38752
rect 8386 38700 8392 38752
rect 8444 38740 8450 38752
rect 8481 38743 8539 38749
rect 8481 38740 8493 38743
rect 8444 38712 8493 38740
rect 8444 38700 8450 38712
rect 8481 38709 8493 38712
rect 8527 38740 8539 38743
rect 8864 38740 8892 38848
rect 9582 38836 9588 38848
rect 9640 38876 9646 38888
rect 9677 38879 9735 38885
rect 9677 38876 9689 38879
rect 9640 38848 9689 38876
rect 9640 38836 9646 38848
rect 9677 38845 9689 38848
rect 9723 38845 9735 38879
rect 10060 38876 10088 38916
rect 10778 38904 10784 38956
rect 10836 38944 10842 38956
rect 12084 38953 12112 38984
rect 12434 38972 12440 38984
rect 12492 38972 12498 39024
rect 12894 38972 12900 39024
rect 12952 38972 12958 39024
rect 13648 39012 13676 39052
rect 14277 39049 14289 39083
rect 14323 39080 14335 39083
rect 15010 39080 15016 39092
rect 14323 39052 15016 39080
rect 14323 39049 14335 39052
rect 14277 39043 14335 39049
rect 15010 39040 15016 39052
rect 15068 39040 15074 39092
rect 15289 39083 15347 39089
rect 15289 39049 15301 39083
rect 15335 39080 15347 39083
rect 15930 39080 15936 39092
rect 15335 39052 15936 39080
rect 15335 39049 15347 39052
rect 15289 39043 15347 39049
rect 15930 39040 15936 39052
rect 15988 39040 15994 39092
rect 16022 39040 16028 39092
rect 16080 39080 16086 39092
rect 19153 39083 19211 39089
rect 19153 39080 19165 39083
rect 16080 39052 19165 39080
rect 16080 39040 16086 39052
rect 19153 39049 19165 39052
rect 19199 39049 19211 39083
rect 19153 39043 19211 39049
rect 19521 39083 19579 39089
rect 19521 39049 19533 39083
rect 19567 39080 19579 39083
rect 20622 39080 20628 39092
rect 19567 39052 20628 39080
rect 19567 39049 19579 39052
rect 19521 39043 19579 39049
rect 20622 39040 20628 39052
rect 20680 39040 20686 39092
rect 20717 39083 20775 39089
rect 20717 39049 20729 39083
rect 20763 39080 20775 39083
rect 20990 39080 20996 39092
rect 20763 39052 20996 39080
rect 20763 39049 20775 39052
rect 20717 39043 20775 39049
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 24489 39083 24547 39089
rect 24489 39080 24501 39083
rect 22066 39052 24501 39080
rect 14458 39012 14464 39024
rect 13648 38984 14464 39012
rect 14458 38972 14464 38984
rect 14516 38972 14522 39024
rect 14826 38972 14832 39024
rect 14884 39012 14890 39024
rect 17218 39012 17224 39024
rect 14884 38984 17224 39012
rect 14884 38972 14890 38984
rect 17218 38972 17224 38984
rect 17276 38972 17282 39024
rect 18325 39015 18383 39021
rect 18325 38981 18337 39015
rect 18371 39012 18383 39015
rect 18598 39012 18604 39024
rect 18371 38984 18604 39012
rect 18371 38981 18383 38984
rect 18325 38975 18383 38981
rect 18598 38972 18604 38984
rect 18656 38972 18662 39024
rect 19613 39015 19671 39021
rect 19613 38981 19625 39015
rect 19659 39012 19671 39015
rect 20806 39012 20812 39024
rect 19659 38984 20812 39012
rect 19659 38981 19671 38984
rect 19613 38975 19671 38981
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 12069 38947 12127 38953
rect 10836 38916 11008 38944
rect 10836 38904 10842 38916
rect 10980 38885 11008 38916
rect 12069 38913 12081 38947
rect 12115 38913 12127 38947
rect 12069 38907 12127 38913
rect 15381 38947 15439 38953
rect 15381 38913 15393 38947
rect 15427 38944 15439 38947
rect 15654 38944 15660 38956
rect 15427 38916 15660 38944
rect 15427 38913 15439 38916
rect 15381 38907 15439 38913
rect 15654 38904 15660 38916
rect 15712 38944 15718 38956
rect 15933 38947 15991 38953
rect 15933 38944 15945 38947
rect 15712 38916 15945 38944
rect 15712 38904 15718 38916
rect 15933 38913 15945 38916
rect 15979 38913 15991 38947
rect 15933 38907 15991 38913
rect 19886 38904 19892 38956
rect 19944 38944 19950 38956
rect 22066 38944 22094 39052
rect 24489 39049 24501 39052
rect 24535 39049 24547 39083
rect 24489 39043 24547 39049
rect 22370 38972 22376 39024
rect 22428 38972 22434 39024
rect 24210 39012 24216 39024
rect 23598 38984 24216 39012
rect 24210 38972 24216 38984
rect 24268 38972 24274 39024
rect 19944 38916 22094 38944
rect 24673 38947 24731 38953
rect 19944 38904 19950 38916
rect 24673 38913 24685 38947
rect 24719 38944 24731 38947
rect 24854 38944 24860 38956
rect 24719 38916 24860 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 24854 38904 24860 38916
rect 24912 38904 24918 38956
rect 25314 38904 25320 38956
rect 25372 38904 25378 38956
rect 10873 38879 10931 38885
rect 10873 38876 10885 38879
rect 10060 38848 10885 38876
rect 9677 38839 9735 38845
rect 8527 38712 8892 38740
rect 8527 38709 8539 38712
rect 8481 38703 8539 38709
rect 9122 38700 9128 38752
rect 9180 38700 9186 38752
rect 10336 38740 10364 38848
rect 10873 38845 10885 38848
rect 10919 38845 10931 38879
rect 10873 38839 10931 38845
rect 10965 38879 11023 38885
rect 10965 38845 10977 38879
rect 11011 38845 11023 38879
rect 10965 38839 11023 38845
rect 12345 38879 12403 38885
rect 12345 38845 12357 38879
rect 12391 38876 12403 38879
rect 14642 38876 14648 38888
rect 12391 38848 14648 38876
rect 12391 38845 12403 38848
rect 12345 38839 12403 38845
rect 14642 38836 14648 38848
rect 14700 38836 14706 38888
rect 15562 38836 15568 38888
rect 15620 38876 15626 38888
rect 16390 38876 16396 38888
rect 15620 38848 16396 38876
rect 15620 38836 15626 38848
rect 16390 38836 16396 38848
rect 16448 38836 16454 38888
rect 16853 38879 16911 38885
rect 16853 38845 16865 38879
rect 16899 38876 16911 38879
rect 17218 38876 17224 38888
rect 16899 38848 17224 38876
rect 16899 38845 16911 38848
rect 16853 38839 16911 38845
rect 17218 38836 17224 38848
rect 17276 38836 17282 38888
rect 18414 38836 18420 38888
rect 18472 38836 18478 38888
rect 18601 38879 18659 38885
rect 18601 38845 18613 38879
rect 18647 38876 18659 38879
rect 19150 38876 19156 38888
rect 18647 38848 19156 38876
rect 18647 38845 18659 38848
rect 18601 38839 18659 38845
rect 19150 38836 19156 38848
rect 19208 38836 19214 38888
rect 19705 38879 19763 38885
rect 19705 38845 19717 38879
rect 19751 38845 19763 38879
rect 19705 38839 19763 38845
rect 10413 38811 10471 38817
rect 10413 38777 10425 38811
rect 10459 38808 10471 38811
rect 11146 38808 11152 38820
rect 10459 38780 11152 38808
rect 10459 38777 10471 38780
rect 10413 38771 10471 38777
rect 11146 38768 11152 38780
rect 11204 38768 11210 38820
rect 11238 38768 11244 38820
rect 11296 38808 11302 38820
rect 13817 38811 13875 38817
rect 11296 38780 11928 38808
rect 11296 38768 11302 38780
rect 11514 38740 11520 38752
rect 10336 38712 11520 38740
rect 11514 38700 11520 38712
rect 11572 38700 11578 38752
rect 11900 38740 11928 38780
rect 13817 38777 13829 38811
rect 13863 38808 13875 38811
rect 13998 38808 14004 38820
rect 13863 38780 14004 38808
rect 13863 38777 13875 38780
rect 13817 38771 13875 38777
rect 13998 38768 14004 38780
rect 14056 38768 14062 38820
rect 18230 38768 18236 38820
rect 18288 38808 18294 38820
rect 19720 38808 19748 38839
rect 20438 38836 20444 38888
rect 20496 38876 20502 38888
rect 20809 38879 20867 38885
rect 20809 38876 20821 38879
rect 20496 38848 20821 38876
rect 20496 38836 20502 38848
rect 20809 38845 20821 38848
rect 20855 38845 20867 38879
rect 20809 38839 20867 38845
rect 20901 38879 20959 38885
rect 20901 38845 20913 38879
rect 20947 38845 20959 38879
rect 20901 38839 20959 38845
rect 18288 38780 19748 38808
rect 18288 38768 18294 38780
rect 18524 38752 18552 38780
rect 19978 38768 19984 38820
rect 20036 38808 20042 38820
rect 20916 38808 20944 38839
rect 22094 38836 22100 38888
rect 22152 38836 22158 38888
rect 22830 38836 22836 38888
rect 22888 38876 22894 38888
rect 24210 38876 24216 38888
rect 22888 38848 24216 38876
rect 22888 38836 22894 38848
rect 24210 38836 24216 38848
rect 24268 38876 24274 38888
rect 25958 38876 25964 38888
rect 24268 38848 25964 38876
rect 24268 38836 24274 38848
rect 25958 38836 25964 38848
rect 26016 38836 26022 38888
rect 20036 38780 20944 38808
rect 20036 38768 20042 38780
rect 23382 38768 23388 38820
rect 23440 38808 23446 38820
rect 25866 38808 25872 38820
rect 23440 38780 25872 38808
rect 23440 38768 23446 38780
rect 25866 38768 25872 38780
rect 25924 38768 25930 38820
rect 12066 38740 12072 38752
rect 11900 38712 12072 38740
rect 12066 38700 12072 38712
rect 12124 38740 12130 38752
rect 13078 38740 13084 38752
rect 12124 38712 13084 38740
rect 12124 38700 12130 38712
rect 13078 38700 13084 38712
rect 13136 38700 13142 38752
rect 13906 38700 13912 38752
rect 13964 38740 13970 38752
rect 14921 38743 14979 38749
rect 14921 38740 14933 38743
rect 13964 38712 14933 38740
rect 13964 38700 13970 38712
rect 14921 38709 14933 38712
rect 14967 38709 14979 38743
rect 14921 38703 14979 38709
rect 17957 38743 18015 38749
rect 17957 38709 17969 38743
rect 18003 38740 18015 38743
rect 18414 38740 18420 38752
rect 18003 38712 18420 38740
rect 18003 38709 18015 38712
rect 17957 38703 18015 38709
rect 18414 38700 18420 38712
rect 18472 38700 18478 38752
rect 18506 38700 18512 38752
rect 18564 38700 18570 38752
rect 18598 38700 18604 38752
rect 18656 38740 18662 38752
rect 18966 38740 18972 38752
rect 18656 38712 18972 38740
rect 18656 38700 18662 38712
rect 18966 38700 18972 38712
rect 19024 38700 19030 38752
rect 20349 38743 20407 38749
rect 20349 38709 20361 38743
rect 20395 38740 20407 38743
rect 21266 38740 21272 38752
rect 20395 38712 21272 38740
rect 20395 38709 20407 38712
rect 20349 38703 20407 38709
rect 21266 38700 21272 38712
rect 21324 38700 21330 38752
rect 22554 38700 22560 38752
rect 22612 38740 22618 38752
rect 23845 38743 23903 38749
rect 23845 38740 23857 38743
rect 22612 38712 23857 38740
rect 22612 38700 22618 38712
rect 23845 38709 23857 38712
rect 23891 38709 23903 38743
rect 23845 38703 23903 38709
rect 25130 38700 25136 38752
rect 25188 38700 25194 38752
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 7558 38496 7564 38548
rect 7616 38536 7622 38548
rect 7837 38539 7895 38545
rect 7837 38536 7849 38539
rect 7616 38508 7849 38536
rect 7616 38496 7622 38508
rect 7837 38505 7849 38508
rect 7883 38505 7895 38539
rect 7837 38499 7895 38505
rect 10413 38539 10471 38545
rect 10413 38505 10425 38539
rect 10459 38536 10471 38539
rect 11054 38536 11060 38548
rect 10459 38508 11060 38536
rect 10459 38505 10471 38508
rect 10413 38499 10471 38505
rect 11054 38496 11060 38508
rect 11112 38496 11118 38548
rect 11882 38496 11888 38548
rect 11940 38496 11946 38548
rect 12342 38496 12348 38548
rect 12400 38536 12406 38548
rect 12526 38536 12532 38548
rect 12400 38508 12532 38536
rect 12400 38496 12406 38508
rect 12526 38496 12532 38508
rect 12584 38496 12590 38548
rect 14182 38496 14188 38548
rect 14240 38536 14246 38548
rect 14277 38539 14335 38545
rect 14277 38536 14289 38539
rect 14240 38508 14289 38536
rect 14240 38496 14246 38508
rect 14277 38505 14289 38508
rect 14323 38505 14335 38539
rect 14277 38499 14335 38505
rect 17402 38496 17408 38548
rect 17460 38536 17466 38548
rect 19429 38539 19487 38545
rect 19429 38536 19441 38539
rect 17460 38508 19441 38536
rect 17460 38496 17466 38508
rect 19429 38505 19441 38508
rect 19475 38505 19487 38539
rect 19429 38499 19487 38505
rect 20625 38539 20683 38545
rect 20625 38505 20637 38539
rect 20671 38536 20683 38539
rect 22186 38536 22192 38548
rect 20671 38508 22192 38536
rect 20671 38505 20683 38508
rect 20625 38499 20683 38505
rect 22186 38496 22192 38508
rect 22244 38496 22250 38548
rect 22370 38496 22376 38548
rect 22428 38536 22434 38548
rect 22428 38508 23612 38536
rect 22428 38496 22434 38508
rect 8570 38468 8576 38480
rect 6840 38440 8576 38468
rect 5721 38403 5779 38409
rect 5721 38369 5733 38403
rect 5767 38400 5779 38403
rect 6840 38400 6868 38440
rect 8570 38428 8576 38440
rect 8628 38428 8634 38480
rect 9214 38428 9220 38480
rect 9272 38468 9278 38480
rect 12710 38468 12716 38480
rect 9272 38440 9904 38468
rect 9272 38428 9278 38440
rect 5767 38372 6868 38400
rect 5767 38369 5779 38372
rect 5721 38363 5779 38369
rect 6914 38360 6920 38412
rect 6972 38400 6978 38412
rect 7193 38403 7251 38409
rect 7193 38400 7205 38403
rect 6972 38372 7205 38400
rect 6972 38360 6978 38372
rect 7193 38369 7205 38372
rect 7239 38400 7251 38403
rect 7834 38400 7840 38412
rect 7239 38372 7840 38400
rect 7239 38369 7251 38372
rect 7193 38363 7251 38369
rect 7834 38360 7840 38372
rect 7892 38360 7898 38412
rect 8481 38403 8539 38409
rect 8481 38369 8493 38403
rect 8527 38369 8539 38403
rect 8481 38363 8539 38369
rect 1302 38292 1308 38344
rect 1360 38332 1366 38344
rect 1765 38335 1823 38341
rect 1765 38332 1777 38335
rect 1360 38304 1777 38332
rect 1360 38292 1366 38304
rect 1765 38301 1777 38304
rect 1811 38332 1823 38335
rect 2041 38335 2099 38341
rect 2041 38332 2053 38335
rect 1811 38304 2053 38332
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 2041 38301 2053 38304
rect 2087 38301 2099 38335
rect 2041 38295 2099 38301
rect 5445 38335 5503 38341
rect 5445 38301 5457 38335
rect 5491 38301 5503 38335
rect 5445 38295 5503 38301
rect 1578 38156 1584 38208
rect 1636 38156 1642 38208
rect 5460 38196 5488 38295
rect 7282 38292 7288 38344
rect 7340 38332 7346 38344
rect 8205 38335 8263 38341
rect 7340 38304 7880 38332
rect 7340 38292 7346 38304
rect 7742 38264 7748 38276
rect 6946 38236 7748 38264
rect 7742 38224 7748 38236
rect 7800 38224 7806 38276
rect 7852 38264 7880 38304
rect 8205 38301 8217 38335
rect 8251 38332 8263 38335
rect 8294 38332 8300 38344
rect 8251 38304 8300 38332
rect 8251 38301 8263 38304
rect 8205 38295 8263 38301
rect 8294 38292 8300 38304
rect 8352 38292 8358 38344
rect 8496 38264 8524 38363
rect 9122 38360 9128 38412
rect 9180 38400 9186 38412
rect 9677 38403 9735 38409
rect 9677 38400 9689 38403
rect 9180 38372 9689 38400
rect 9180 38360 9186 38372
rect 9677 38369 9689 38372
rect 9723 38369 9735 38403
rect 9677 38363 9735 38369
rect 9769 38403 9827 38409
rect 9769 38369 9781 38403
rect 9815 38369 9827 38403
rect 9876 38400 9904 38440
rect 10980 38440 12716 38468
rect 10980 38409 11008 38440
rect 12710 38428 12716 38440
rect 12768 38468 12774 38480
rect 12768 38440 14872 38468
rect 12768 38428 12774 38440
rect 10965 38403 11023 38409
rect 10965 38400 10977 38403
rect 9876 38372 10977 38400
rect 9769 38363 9827 38369
rect 10965 38369 10977 38372
rect 11011 38369 11023 38403
rect 10965 38363 11023 38369
rect 9214 38292 9220 38344
rect 9272 38332 9278 38344
rect 9784 38332 9812 38363
rect 12158 38360 12164 38412
rect 12216 38400 12222 38412
rect 12345 38403 12403 38409
rect 12345 38400 12357 38403
rect 12216 38372 12357 38400
rect 12216 38360 12222 38372
rect 12345 38369 12357 38372
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 12437 38403 12495 38409
rect 12437 38369 12449 38403
rect 12483 38369 12495 38403
rect 12437 38363 12495 38369
rect 13909 38403 13967 38409
rect 13909 38369 13921 38403
rect 13955 38400 13967 38403
rect 14274 38400 14280 38412
rect 13955 38372 14280 38400
rect 13955 38369 13967 38372
rect 13909 38363 13967 38369
rect 9272 38304 9812 38332
rect 9272 38292 9278 38304
rect 10594 38292 10600 38344
rect 10652 38332 10658 38344
rect 12452 38332 12480 38363
rect 14274 38360 14280 38372
rect 14332 38360 14338 38412
rect 14844 38409 14872 38440
rect 17862 38428 17868 38480
rect 17920 38468 17926 38480
rect 18141 38471 18199 38477
rect 18141 38468 18153 38471
rect 17920 38440 18153 38468
rect 17920 38428 17926 38440
rect 18141 38437 18153 38440
rect 18187 38437 18199 38471
rect 20806 38468 20812 38480
rect 18141 38431 18199 38437
rect 18524 38440 20812 38468
rect 14829 38403 14887 38409
rect 14829 38369 14841 38403
rect 14875 38369 14887 38403
rect 14829 38363 14887 38369
rect 15010 38360 15016 38412
rect 15068 38400 15074 38412
rect 16209 38403 16267 38409
rect 16209 38400 16221 38403
rect 15068 38372 16221 38400
rect 15068 38360 15074 38372
rect 16209 38369 16221 38372
rect 16255 38400 16267 38403
rect 18230 38400 18236 38412
rect 16255 38372 18236 38400
rect 16255 38369 16267 38372
rect 16209 38363 16267 38369
rect 18230 38360 18236 38372
rect 18288 38360 18294 38412
rect 10652 38304 12480 38332
rect 14737 38335 14795 38341
rect 10652 38292 10658 38304
rect 14737 38301 14749 38335
rect 14783 38332 14795 38335
rect 15378 38332 15384 38344
rect 14783 38304 15384 38332
rect 14783 38301 14795 38304
rect 14737 38295 14795 38301
rect 15378 38292 15384 38304
rect 15436 38292 15442 38344
rect 15930 38292 15936 38344
rect 15988 38292 15994 38344
rect 17586 38332 17592 38344
rect 17342 38304 17592 38332
rect 17586 38292 17592 38304
rect 17644 38292 17650 38344
rect 18524 38341 18552 38440
rect 20806 38428 20812 38440
rect 20864 38428 20870 38480
rect 22005 38471 22063 38477
rect 22005 38437 22017 38471
rect 22051 38468 22063 38471
rect 22738 38468 22744 38480
rect 22051 38440 22744 38468
rect 22051 38437 22063 38440
rect 22005 38431 22063 38437
rect 22738 38428 22744 38440
rect 22796 38428 22802 38480
rect 18690 38360 18696 38412
rect 18748 38360 18754 38412
rect 19242 38360 19248 38412
rect 19300 38400 19306 38412
rect 19981 38403 20039 38409
rect 19981 38400 19993 38403
rect 19300 38372 19993 38400
rect 19300 38360 19306 38372
rect 19981 38369 19993 38372
rect 20027 38369 20039 38403
rect 19981 38363 20039 38369
rect 20254 38360 20260 38412
rect 20312 38400 20318 38412
rect 21085 38403 21143 38409
rect 21085 38400 21097 38403
rect 20312 38372 21097 38400
rect 20312 38360 20318 38372
rect 21085 38369 21097 38372
rect 21131 38369 21143 38403
rect 21085 38363 21143 38369
rect 21174 38360 21180 38412
rect 21232 38360 21238 38412
rect 21910 38360 21916 38412
rect 21968 38400 21974 38412
rect 22465 38403 22523 38409
rect 22465 38400 22477 38403
rect 21968 38372 22477 38400
rect 21968 38360 21974 38372
rect 22465 38369 22477 38372
rect 22511 38369 22523 38403
rect 22465 38363 22523 38369
rect 22554 38360 22560 38412
rect 22612 38360 22618 38412
rect 23584 38400 23612 38508
rect 23753 38403 23811 38409
rect 23753 38400 23765 38403
rect 23584 38372 23765 38400
rect 23753 38369 23765 38372
rect 23799 38369 23811 38403
rect 23753 38363 23811 38369
rect 23842 38360 23848 38412
rect 23900 38400 23906 38412
rect 25133 38403 25191 38409
rect 25133 38400 25145 38403
rect 23900 38372 25145 38400
rect 23900 38360 23906 38372
rect 25133 38369 25145 38372
rect 25179 38369 25191 38403
rect 25133 38363 25191 38369
rect 18509 38335 18567 38341
rect 18509 38301 18521 38335
rect 18555 38301 18567 38335
rect 18509 38295 18567 38301
rect 18966 38292 18972 38344
rect 19024 38332 19030 38344
rect 20993 38335 21051 38341
rect 20993 38332 21005 38335
rect 19024 38304 21005 38332
rect 19024 38292 19030 38304
rect 20993 38301 21005 38304
rect 21039 38301 21051 38335
rect 24026 38332 24032 38344
rect 20993 38295 21051 38301
rect 21836 38304 24032 38332
rect 9585 38267 9643 38273
rect 7852 38236 9352 38264
rect 6546 38196 6552 38208
rect 5460 38168 6552 38196
rect 6546 38156 6552 38168
rect 6604 38156 6610 38208
rect 7098 38156 7104 38208
rect 7156 38196 7162 38208
rect 7561 38199 7619 38205
rect 7561 38196 7573 38199
rect 7156 38168 7573 38196
rect 7156 38156 7162 38168
rect 7561 38165 7573 38168
rect 7607 38196 7619 38199
rect 8202 38196 8208 38208
rect 7607 38168 8208 38196
rect 7607 38165 7619 38168
rect 7561 38159 7619 38165
rect 8202 38156 8208 38168
rect 8260 38196 8266 38208
rect 8297 38199 8355 38205
rect 8297 38196 8309 38199
rect 8260 38168 8309 38196
rect 8260 38156 8266 38168
rect 8297 38165 8309 38168
rect 8343 38165 8355 38199
rect 8297 38159 8355 38165
rect 8478 38156 8484 38208
rect 8536 38196 8542 38208
rect 9217 38199 9275 38205
rect 9217 38196 9229 38199
rect 8536 38168 9229 38196
rect 8536 38156 8542 38168
rect 9217 38165 9229 38168
rect 9263 38165 9275 38199
rect 9324 38196 9352 38236
rect 9585 38233 9597 38267
rect 9631 38264 9643 38267
rect 9674 38264 9680 38276
rect 9631 38236 9680 38264
rect 9631 38233 9643 38236
rect 9585 38227 9643 38233
rect 9674 38224 9680 38236
rect 9732 38224 9738 38276
rect 19518 38264 19524 38276
rect 17604 38236 19524 38264
rect 10594 38196 10600 38208
rect 9324 38168 10600 38196
rect 9217 38159 9275 38165
rect 10594 38156 10600 38168
rect 10652 38156 10658 38208
rect 10778 38156 10784 38208
rect 10836 38156 10842 38208
rect 10870 38156 10876 38208
rect 10928 38156 10934 38208
rect 12253 38199 12311 38205
rect 12253 38165 12265 38199
rect 12299 38196 12311 38199
rect 12526 38196 12532 38208
rect 12299 38168 12532 38196
rect 12299 38165 12311 38168
rect 12253 38159 12311 38165
rect 12526 38156 12532 38168
rect 12584 38196 12590 38208
rect 12897 38199 12955 38205
rect 12897 38196 12909 38199
rect 12584 38168 12909 38196
rect 12584 38156 12590 38168
rect 12897 38165 12909 38168
rect 12943 38165 12955 38199
rect 12897 38159 12955 38165
rect 13262 38156 13268 38208
rect 13320 38156 13326 38208
rect 13538 38156 13544 38208
rect 13596 38196 13602 38208
rect 13814 38196 13820 38208
rect 13596 38168 13820 38196
rect 13596 38156 13602 38168
rect 13814 38156 13820 38168
rect 13872 38156 13878 38208
rect 14645 38199 14703 38205
rect 14645 38165 14657 38199
rect 14691 38196 14703 38199
rect 17604 38196 17632 38236
rect 19518 38224 19524 38236
rect 19576 38224 19582 38276
rect 19886 38224 19892 38276
rect 19944 38224 19950 38276
rect 14691 38168 17632 38196
rect 14691 38165 14703 38168
rect 14645 38159 14703 38165
rect 17678 38156 17684 38208
rect 17736 38156 17742 38208
rect 18601 38199 18659 38205
rect 18601 38165 18613 38199
rect 18647 38196 18659 38199
rect 19058 38196 19064 38208
rect 18647 38168 19064 38196
rect 18647 38165 18659 38168
rect 18601 38159 18659 38165
rect 19058 38156 19064 38168
rect 19116 38156 19122 38208
rect 19797 38199 19855 38205
rect 19797 38165 19809 38199
rect 19843 38196 19855 38199
rect 20438 38196 20444 38208
rect 19843 38168 20444 38196
rect 19843 38165 19855 38168
rect 19797 38159 19855 38165
rect 20438 38156 20444 38168
rect 20496 38156 20502 38208
rect 21082 38156 21088 38208
rect 21140 38196 21146 38208
rect 21637 38199 21695 38205
rect 21637 38196 21649 38199
rect 21140 38168 21649 38196
rect 21140 38156 21146 38168
rect 21637 38165 21649 38168
rect 21683 38196 21695 38199
rect 21836 38196 21864 38304
rect 24026 38292 24032 38304
rect 24084 38292 24090 38344
rect 24946 38292 24952 38344
rect 25004 38332 25010 38344
rect 25041 38335 25099 38341
rect 25041 38332 25053 38335
rect 25004 38304 25053 38332
rect 25004 38292 25010 38304
rect 25041 38301 25053 38304
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 22373 38267 22431 38273
rect 22373 38233 22385 38267
rect 22419 38264 22431 38267
rect 22419 38236 23244 38264
rect 22419 38233 22431 38236
rect 22373 38227 22431 38233
rect 23216 38205 23244 38236
rect 23566 38224 23572 38276
rect 23624 38224 23630 38276
rect 23661 38267 23719 38273
rect 23661 38233 23673 38267
rect 23707 38264 23719 38267
rect 24210 38264 24216 38276
rect 23707 38236 24216 38264
rect 23707 38233 23719 38236
rect 23661 38227 23719 38233
rect 24210 38224 24216 38236
rect 24268 38224 24274 38276
rect 21683 38168 21864 38196
rect 23201 38199 23259 38205
rect 21683 38165 21695 38168
rect 21637 38159 21695 38165
rect 23201 38165 23213 38199
rect 23247 38165 23259 38199
rect 23201 38159 23259 38165
rect 23750 38156 23756 38208
rect 23808 38196 23814 38208
rect 24581 38199 24639 38205
rect 24581 38196 24593 38199
rect 23808 38168 24593 38196
rect 23808 38156 23814 38168
rect 24581 38165 24593 38168
rect 24627 38165 24639 38199
rect 24581 38159 24639 38165
rect 24670 38156 24676 38208
rect 24728 38196 24734 38208
rect 24949 38199 25007 38205
rect 24949 38196 24961 38199
rect 24728 38168 24961 38196
rect 24728 38156 24734 38168
rect 24949 38165 24961 38168
rect 24995 38165 25007 38199
rect 24949 38159 25007 38165
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 5258 37952 5264 38004
rect 5316 37952 5322 38004
rect 5721 37995 5779 38001
rect 5721 37961 5733 37995
rect 5767 37992 5779 37995
rect 8938 37992 8944 38004
rect 5767 37964 8944 37992
rect 5767 37961 5779 37964
rect 5721 37955 5779 37961
rect 8938 37952 8944 37964
rect 8996 37952 9002 38004
rect 9125 37995 9183 38001
rect 9125 37961 9137 37995
rect 9171 37992 9183 37995
rect 9306 37992 9312 38004
rect 9171 37964 9312 37992
rect 9171 37961 9183 37964
rect 9125 37955 9183 37961
rect 9306 37952 9312 37964
rect 9364 37952 9370 38004
rect 10045 37995 10103 38001
rect 10045 37961 10057 37995
rect 10091 37992 10103 37995
rect 10502 37992 10508 38004
rect 10091 37964 10508 37992
rect 10091 37961 10103 37964
rect 10045 37955 10103 37961
rect 10502 37952 10508 37964
rect 10560 37952 10566 38004
rect 10778 37952 10784 38004
rect 10836 37992 10842 38004
rect 11701 37995 11759 38001
rect 11701 37992 11713 37995
rect 10836 37964 11713 37992
rect 10836 37952 10842 37964
rect 11701 37961 11713 37964
rect 11747 37961 11759 37995
rect 11701 37955 11759 37961
rect 11790 37952 11796 38004
rect 11848 37992 11854 38004
rect 12345 37995 12403 38001
rect 12345 37992 12357 37995
rect 11848 37964 12357 37992
rect 11848 37952 11854 37964
rect 12345 37961 12357 37964
rect 12391 37961 12403 37995
rect 12345 37955 12403 37961
rect 12713 37995 12771 38001
rect 12713 37961 12725 37995
rect 12759 37992 12771 37995
rect 13262 37992 13268 38004
rect 12759 37964 13268 37992
rect 12759 37961 12771 37964
rect 12713 37955 12771 37961
rect 13262 37952 13268 37964
rect 13320 37952 13326 38004
rect 15378 37992 15384 38004
rect 13924 37964 15384 37992
rect 6825 37927 6883 37933
rect 6825 37893 6837 37927
rect 6871 37924 6883 37927
rect 6914 37924 6920 37936
rect 6871 37896 6920 37924
rect 6871 37893 6883 37896
rect 6825 37887 6883 37893
rect 6914 37884 6920 37896
rect 6972 37884 6978 37936
rect 7834 37884 7840 37936
rect 7892 37884 7898 37936
rect 9324 37924 9352 37952
rect 9324 37896 10548 37924
rect 4982 37816 4988 37868
rect 5040 37856 5046 37868
rect 5629 37859 5687 37865
rect 5629 37856 5641 37859
rect 5040 37828 5641 37856
rect 5040 37816 5046 37828
rect 5629 37825 5641 37828
rect 5675 37825 5687 37859
rect 5629 37819 5687 37825
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37856 9459 37859
rect 10413 37859 10471 37865
rect 10413 37856 10425 37859
rect 9447 37828 10425 37856
rect 9447 37825 9459 37828
rect 9401 37819 9459 37825
rect 10413 37825 10425 37828
rect 10459 37825 10471 37859
rect 10520 37856 10548 37896
rect 11330 37884 11336 37936
rect 11388 37884 11394 37936
rect 13924 37856 13952 37964
rect 15378 37952 15384 37964
rect 15436 37952 15442 38004
rect 15473 37995 15531 38001
rect 15473 37961 15485 37995
rect 15519 37992 15531 37995
rect 16298 37992 16304 38004
rect 15519 37964 16304 37992
rect 15519 37961 15531 37964
rect 15473 37955 15531 37961
rect 16298 37952 16304 37964
rect 16356 37952 16362 38004
rect 17218 37952 17224 38004
rect 17276 37952 17282 38004
rect 17586 37952 17592 38004
rect 17644 37992 17650 38004
rect 18049 37995 18107 38001
rect 18049 37992 18061 37995
rect 17644 37964 18061 37992
rect 17644 37952 17650 37964
rect 18049 37961 18061 37964
rect 18095 37961 18107 37995
rect 18049 37955 18107 37961
rect 18325 37995 18383 38001
rect 18325 37961 18337 37995
rect 18371 37992 18383 37995
rect 18690 37992 18696 38004
rect 18371 37964 18696 37992
rect 18371 37961 18383 37964
rect 18325 37955 18383 37961
rect 18690 37952 18696 37964
rect 18748 37952 18754 38004
rect 18969 37995 19027 38001
rect 18969 37961 18981 37995
rect 19015 37992 19027 37995
rect 20898 37992 20904 38004
rect 19015 37964 20904 37992
rect 19015 37961 19027 37964
rect 18969 37955 19027 37961
rect 20898 37952 20904 37964
rect 20956 37952 20962 38004
rect 21545 37995 21603 38001
rect 21545 37961 21557 37995
rect 21591 37992 21603 37995
rect 21818 37992 21824 38004
rect 21591 37964 21824 37992
rect 21591 37961 21603 37964
rect 21545 37955 21603 37961
rect 17862 37924 17868 37936
rect 10520 37828 13952 37856
rect 14108 37896 17868 37924
rect 10413 37819 10471 37825
rect 5810 37748 5816 37800
rect 5868 37748 5874 37800
rect 6546 37748 6552 37800
rect 6604 37748 6610 37800
rect 7282 37748 7288 37800
rect 7340 37788 7346 37800
rect 8386 37788 8392 37800
rect 7340 37760 8392 37788
rect 7340 37748 7346 37760
rect 8386 37748 8392 37760
rect 8444 37788 8450 37800
rect 8573 37791 8631 37797
rect 8573 37788 8585 37791
rect 8444 37760 8585 37788
rect 8444 37748 8450 37760
rect 8573 37757 8585 37760
rect 8619 37757 8631 37791
rect 8573 37751 8631 37757
rect 8941 37791 8999 37797
rect 8941 37757 8953 37791
rect 8987 37788 8999 37791
rect 10502 37788 10508 37800
rect 8987 37760 10508 37788
rect 8987 37757 8999 37760
rect 8941 37751 8999 37757
rect 6638 37612 6644 37664
rect 6696 37652 6702 37664
rect 8956 37652 8984 37751
rect 10502 37748 10508 37760
rect 10560 37748 10566 37800
rect 10612 37797 10640 37828
rect 10597 37791 10655 37797
rect 10597 37757 10609 37791
rect 10643 37757 10655 37791
rect 12805 37791 12863 37797
rect 12805 37788 12817 37791
rect 10597 37751 10655 37757
rect 12636 37760 12817 37788
rect 11330 37680 11336 37732
rect 11388 37720 11394 37732
rect 12636 37720 12664 37760
rect 12805 37757 12817 37760
rect 12851 37757 12863 37791
rect 12805 37751 12863 37757
rect 12989 37791 13047 37797
rect 12989 37757 13001 37791
rect 13035 37788 13047 37791
rect 13446 37788 13452 37800
rect 13035 37760 13452 37788
rect 13035 37757 13047 37760
rect 12989 37751 13047 37757
rect 13446 37748 13452 37760
rect 13504 37748 13510 37800
rect 13538 37748 13544 37800
rect 13596 37748 13602 37800
rect 14108 37788 14136 37896
rect 17862 37884 17868 37896
rect 17920 37884 17926 37936
rect 18230 37884 18236 37936
rect 18288 37924 18294 37936
rect 18509 37927 18567 37933
rect 18509 37924 18521 37927
rect 18288 37896 18521 37924
rect 18288 37884 18294 37896
rect 18509 37893 18521 37896
rect 18555 37924 18567 37927
rect 19242 37924 19248 37936
rect 18555 37896 19248 37924
rect 18555 37893 18567 37896
rect 18509 37887 18567 37893
rect 19242 37884 19248 37896
rect 19300 37884 19306 37936
rect 19429 37927 19487 37933
rect 19429 37893 19441 37927
rect 19475 37924 19487 37927
rect 19475 37896 20024 37924
rect 19475 37893 19487 37896
rect 19429 37887 19487 37893
rect 14369 37859 14427 37865
rect 14369 37825 14381 37859
rect 14415 37856 14427 37859
rect 15381 37859 15439 37865
rect 15381 37856 15393 37859
rect 14415 37828 15393 37856
rect 14415 37825 14427 37828
rect 14369 37819 14427 37825
rect 15381 37825 15393 37828
rect 15427 37825 15439 37859
rect 17313 37859 17371 37865
rect 17313 37856 17325 37859
rect 15381 37819 15439 37825
rect 17236 37828 17325 37856
rect 13924 37760 14136 37788
rect 11388 37692 12664 37720
rect 11388 37680 11394 37692
rect 6696 37624 8984 37652
rect 6696 37612 6702 37624
rect 9582 37612 9588 37664
rect 9640 37652 9646 37664
rect 13924 37652 13952 37760
rect 15562 37748 15568 37800
rect 15620 37788 15626 37800
rect 15657 37791 15715 37797
rect 15657 37788 15669 37791
rect 15620 37760 15669 37788
rect 15620 37748 15626 37760
rect 15657 37757 15669 37760
rect 15703 37788 15715 37791
rect 16114 37788 16120 37800
rect 15703 37760 16120 37788
rect 15703 37757 15715 37760
rect 15657 37751 15715 37757
rect 16114 37748 16120 37760
rect 16172 37748 16178 37800
rect 14274 37680 14280 37732
rect 14332 37720 14338 37732
rect 15013 37723 15071 37729
rect 15013 37720 15025 37723
rect 14332 37692 15025 37720
rect 14332 37680 14338 37692
rect 15013 37689 15025 37692
rect 15059 37689 15071 37723
rect 15013 37683 15071 37689
rect 16390 37680 16396 37732
rect 16448 37720 16454 37732
rect 17236 37720 17264 37828
rect 17313 37825 17325 37828
rect 17359 37825 17371 37859
rect 17313 37819 17371 37825
rect 18598 37816 18604 37868
rect 18656 37856 18662 37868
rect 19337 37859 19395 37865
rect 19337 37856 19349 37859
rect 18656 37828 19349 37856
rect 18656 37816 18662 37828
rect 19337 37825 19349 37828
rect 19383 37825 19395 37859
rect 19996 37856 20024 37896
rect 20070 37884 20076 37936
rect 20128 37924 20134 37936
rect 20625 37927 20683 37933
rect 20625 37924 20637 37927
rect 20128 37896 20637 37924
rect 20128 37884 20134 37896
rect 20625 37893 20637 37896
rect 20671 37924 20683 37927
rect 21269 37927 21327 37933
rect 21269 37924 21281 37927
rect 20671 37896 21281 37924
rect 20671 37893 20683 37896
rect 20625 37887 20683 37893
rect 21269 37893 21281 37896
rect 21315 37893 21327 37927
rect 21269 37887 21327 37893
rect 20717 37859 20775 37865
rect 20717 37856 20729 37859
rect 19996 37828 20729 37856
rect 19337 37819 19395 37825
rect 20717 37825 20729 37828
rect 20763 37856 20775 37859
rect 21082 37856 21088 37868
rect 20763 37828 21088 37856
rect 20763 37825 20775 37828
rect 20717 37819 20775 37825
rect 21082 37816 21088 37828
rect 21140 37816 21146 37868
rect 17497 37791 17555 37797
rect 17497 37757 17509 37791
rect 17543 37788 17555 37791
rect 17770 37788 17776 37800
rect 17543 37760 17776 37788
rect 17543 37757 17555 37760
rect 17497 37751 17555 37757
rect 17770 37748 17776 37760
rect 17828 37748 17834 37800
rect 19610 37748 19616 37800
rect 19668 37748 19674 37800
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 21560 37788 21588 37955
rect 21818 37952 21824 37964
rect 21876 37952 21882 38004
rect 22005 37995 22063 38001
rect 22005 37961 22017 37995
rect 22051 37992 22063 37995
rect 24670 37992 24676 38004
rect 22051 37964 24676 37992
rect 22051 37961 22063 37964
rect 22005 37955 22063 37961
rect 24670 37952 24676 37964
rect 24728 37952 24734 38004
rect 22465 37927 22523 37933
rect 22465 37893 22477 37927
rect 22511 37924 22523 37927
rect 23109 37927 23167 37933
rect 23109 37924 23121 37927
rect 22511 37896 23121 37924
rect 22511 37893 22523 37896
rect 22465 37887 22523 37893
rect 23109 37893 23121 37896
rect 23155 37924 23167 37927
rect 23382 37924 23388 37936
rect 23155 37896 23388 37924
rect 23155 37893 23167 37896
rect 23109 37887 23167 37893
rect 23382 37884 23388 37896
rect 23440 37884 23446 37936
rect 23842 37884 23848 37936
rect 23900 37884 23906 37936
rect 24854 37884 24860 37936
rect 24912 37884 24918 37936
rect 22373 37859 22431 37865
rect 22373 37825 22385 37859
rect 22419 37856 22431 37859
rect 23198 37856 23204 37868
rect 22419 37828 23204 37856
rect 22419 37825 22431 37828
rect 22373 37819 22431 37825
rect 23198 37816 23204 37828
rect 23256 37816 23262 37868
rect 20947 37760 21588 37788
rect 22649 37791 22707 37797
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 22649 37757 22661 37791
rect 22695 37788 22707 37791
rect 22830 37788 22836 37800
rect 22695 37760 22836 37788
rect 22695 37757 22707 37760
rect 22649 37751 22707 37757
rect 22830 37748 22836 37760
rect 22888 37748 22894 37800
rect 23569 37791 23627 37797
rect 23569 37757 23581 37791
rect 23615 37757 23627 37791
rect 23569 37751 23627 37757
rect 16448 37692 17264 37720
rect 16448 37680 16454 37692
rect 17402 37680 17408 37732
rect 17460 37720 17466 37732
rect 19794 37720 19800 37732
rect 17460 37692 19800 37720
rect 17460 37680 17466 37692
rect 19794 37680 19800 37692
rect 19852 37680 19858 37732
rect 20257 37723 20315 37729
rect 20257 37689 20269 37723
rect 20303 37720 20315 37723
rect 22002 37720 22008 37732
rect 20303 37692 22008 37720
rect 20303 37689 20315 37692
rect 20257 37683 20315 37689
rect 22002 37680 22008 37692
rect 22060 37680 22066 37732
rect 22094 37680 22100 37732
rect 22152 37720 22158 37732
rect 23584 37720 23612 37751
rect 24486 37748 24492 37800
rect 24544 37788 24550 37800
rect 25317 37791 25375 37797
rect 25317 37788 25329 37791
rect 24544 37760 25329 37788
rect 24544 37748 24550 37760
rect 25317 37757 25329 37760
rect 25363 37757 25375 37791
rect 25317 37751 25375 37757
rect 22152 37692 23612 37720
rect 22152 37680 22158 37692
rect 9640 37624 13952 37652
rect 14093 37655 14151 37661
rect 9640 37612 9646 37624
rect 14093 37621 14105 37655
rect 14139 37652 14151 37655
rect 14366 37652 14372 37664
rect 14139 37624 14372 37652
rect 14139 37621 14151 37624
rect 14093 37615 14151 37621
rect 14366 37612 14372 37624
rect 14424 37652 14430 37664
rect 15194 37652 15200 37664
rect 14424 37624 15200 37652
rect 14424 37612 14430 37624
rect 15194 37612 15200 37624
rect 15252 37612 15258 37664
rect 16117 37655 16175 37661
rect 16117 37621 16129 37655
rect 16163 37652 16175 37655
rect 16298 37652 16304 37664
rect 16163 37624 16304 37652
rect 16163 37621 16175 37624
rect 16117 37615 16175 37621
rect 16298 37612 16304 37624
rect 16356 37612 16362 37664
rect 16853 37655 16911 37661
rect 16853 37621 16865 37655
rect 16899 37652 16911 37655
rect 18322 37652 18328 37664
rect 16899 37624 18328 37652
rect 16899 37621 16911 37624
rect 16853 37615 16911 37621
rect 18322 37612 18328 37624
rect 18380 37612 18386 37664
rect 18598 37612 18604 37664
rect 18656 37612 18662 37664
rect 19288 37612 19294 37664
rect 19346 37652 19352 37664
rect 20070 37652 20076 37664
rect 19346 37624 20076 37652
rect 19346 37612 19352 37624
rect 20070 37612 20076 37624
rect 20128 37612 20134 37664
rect 23566 37612 23572 37664
rect 23624 37652 23630 37664
rect 24026 37652 24032 37664
rect 23624 37624 24032 37652
rect 23624 37612 23630 37624
rect 24026 37612 24032 37624
rect 24084 37612 24090 37664
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 8570 37408 8576 37460
rect 8628 37408 8634 37460
rect 10410 37408 10416 37460
rect 10468 37408 10474 37460
rect 10597 37451 10655 37457
rect 10597 37417 10609 37451
rect 10643 37448 10655 37451
rect 11698 37448 11704 37460
rect 10643 37420 11704 37448
rect 10643 37417 10655 37420
rect 10597 37411 10655 37417
rect 11698 37408 11704 37420
rect 11756 37408 11762 37460
rect 12250 37408 12256 37460
rect 12308 37448 12314 37460
rect 14921 37451 14979 37457
rect 14921 37448 14933 37451
rect 12308 37420 14933 37448
rect 12308 37408 12314 37420
rect 14921 37417 14933 37420
rect 14967 37417 14979 37451
rect 18690 37448 18696 37460
rect 14921 37411 14979 37417
rect 15028 37420 18696 37448
rect 12434 37340 12440 37392
rect 12492 37380 12498 37392
rect 12802 37380 12808 37392
rect 12492 37352 12808 37380
rect 12492 37340 12498 37352
rect 12802 37340 12808 37352
rect 12860 37340 12866 37392
rect 12897 37383 12955 37389
rect 12897 37349 12909 37383
rect 12943 37349 12955 37383
rect 12897 37343 12955 37349
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 8754 37312 8760 37324
rect 7147 37284 8760 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 8754 37272 8760 37284
rect 8812 37272 8818 37324
rect 10962 37272 10968 37324
rect 11020 37312 11026 37324
rect 11793 37315 11851 37321
rect 11793 37312 11805 37315
rect 11020 37284 11805 37312
rect 11020 37272 11026 37284
rect 11793 37281 11805 37284
rect 11839 37281 11851 37315
rect 11793 37275 11851 37281
rect 6546 37204 6552 37256
rect 6604 37244 6610 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6604 37216 6837 37244
rect 6604 37204 6610 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 6825 37207 6883 37213
rect 8404 37216 9873 37244
rect 6840 37108 6868 37207
rect 7742 37136 7748 37188
rect 7800 37136 7806 37188
rect 8404 37108 8432 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 10042 37204 10048 37256
rect 10100 37244 10106 37256
rect 11609 37247 11667 37253
rect 10100 37216 11284 37244
rect 10100 37204 10106 37216
rect 9125 37179 9183 37185
rect 9125 37145 9137 37179
rect 9171 37176 9183 37179
rect 10410 37176 10416 37188
rect 9171 37148 10416 37176
rect 9171 37145 9183 37148
rect 9125 37139 9183 37145
rect 10410 37136 10416 37148
rect 10468 37136 10474 37188
rect 11256 37117 11284 37216
rect 11609 37213 11621 37247
rect 11655 37244 11667 37247
rect 11882 37244 11888 37256
rect 11655 37216 11888 37244
rect 11655 37213 11667 37216
rect 11609 37207 11667 37213
rect 11882 37204 11888 37216
rect 11940 37204 11946 37256
rect 12912 37244 12940 37343
rect 12986 37340 12992 37392
rect 13044 37380 13050 37392
rect 13044 37352 13400 37380
rect 13044 37340 13050 37352
rect 13372 37321 13400 37352
rect 14458 37340 14464 37392
rect 14516 37380 14522 37392
rect 14553 37383 14611 37389
rect 14553 37380 14565 37383
rect 14516 37352 14565 37380
rect 14516 37340 14522 37352
rect 14553 37349 14565 37352
rect 14599 37349 14611 37383
rect 14553 37343 14611 37349
rect 13357 37315 13415 37321
rect 13357 37281 13369 37315
rect 13403 37281 13415 37315
rect 13357 37275 13415 37281
rect 13449 37315 13507 37321
rect 13449 37281 13461 37315
rect 13495 37312 13507 37315
rect 14090 37312 14096 37324
rect 13495 37284 14096 37312
rect 13495 37281 13507 37284
rect 13449 37275 13507 37281
rect 14090 37272 14096 37284
rect 14148 37272 14154 37324
rect 14182 37272 14188 37324
rect 14240 37312 14246 37324
rect 15028 37312 15056 37420
rect 18690 37408 18696 37420
rect 18748 37408 18754 37460
rect 21818 37408 21824 37460
rect 21876 37448 21882 37460
rect 25222 37448 25228 37460
rect 21876 37420 25228 37448
rect 21876 37408 21882 37420
rect 25222 37408 25228 37420
rect 25280 37408 25286 37460
rect 15746 37340 15752 37392
rect 15804 37380 15810 37392
rect 15804 37352 16712 37380
rect 15804 37340 15810 37352
rect 14240 37284 15056 37312
rect 14240 37272 14246 37284
rect 15378 37272 15384 37324
rect 15436 37312 15442 37324
rect 15473 37315 15531 37321
rect 15473 37312 15485 37315
rect 15436 37284 15485 37312
rect 15436 37272 15442 37284
rect 15473 37281 15485 37284
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 16206 37272 16212 37324
rect 16264 37312 16270 37324
rect 16684 37321 16712 37352
rect 17034 37340 17040 37392
rect 17092 37380 17098 37392
rect 17313 37383 17371 37389
rect 17313 37380 17325 37383
rect 17092 37352 17325 37380
rect 17092 37340 17098 37352
rect 17313 37349 17325 37352
rect 17359 37349 17371 37383
rect 17313 37343 17371 37349
rect 22462 37340 22468 37392
rect 22520 37380 22526 37392
rect 24118 37380 24124 37392
rect 22520 37352 24124 37380
rect 22520 37340 22526 37352
rect 24118 37340 24124 37352
rect 24176 37340 24182 37392
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 16264 37284 16589 37312
rect 16264 37272 16270 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 16669 37315 16727 37321
rect 16669 37281 16681 37315
rect 16715 37281 16727 37315
rect 16669 37275 16727 37281
rect 17862 37272 17868 37324
rect 17920 37272 17926 37324
rect 18506 37272 18512 37324
rect 18564 37312 18570 37324
rect 18690 37312 18696 37324
rect 18564 37284 18696 37312
rect 18564 37272 18570 37284
rect 18690 37272 18696 37284
rect 18748 37272 18754 37324
rect 19061 37315 19119 37321
rect 19061 37281 19073 37315
rect 19107 37312 19119 37315
rect 19242 37312 19248 37324
rect 19107 37284 19248 37312
rect 19107 37281 19119 37284
rect 19061 37275 19119 37281
rect 13265 37247 13323 37253
rect 12912 37216 13216 37244
rect 11701 37179 11759 37185
rect 11701 37145 11713 37179
rect 11747 37176 11759 37179
rect 13188 37176 13216 37216
rect 13265 37213 13277 37247
rect 13311 37244 13323 37247
rect 13538 37244 13544 37256
rect 13311 37216 13544 37244
rect 13311 37213 13323 37216
rect 13265 37207 13323 37213
rect 13538 37204 13544 37216
rect 13596 37204 13602 37256
rect 17773 37247 17831 37253
rect 17773 37213 17785 37247
rect 17819 37244 17831 37247
rect 19076 37244 19104 37275
rect 19242 37272 19248 37284
rect 19300 37312 19306 37324
rect 23658 37312 23664 37324
rect 19300 37284 23664 37312
rect 19300 37272 19306 37284
rect 23658 37272 23664 37284
rect 23716 37272 23722 37324
rect 24026 37272 24032 37324
rect 24084 37272 24090 37324
rect 24213 37315 24271 37321
rect 24213 37281 24225 37315
rect 24259 37312 24271 37315
rect 24394 37312 24400 37324
rect 24259 37284 24400 37312
rect 24259 37281 24271 37284
rect 24213 37275 24271 37281
rect 24394 37272 24400 37284
rect 24452 37272 24458 37324
rect 24581 37315 24639 37321
rect 24581 37281 24593 37315
rect 24627 37312 24639 37315
rect 24627 37284 25360 37312
rect 24627 37281 24639 37284
rect 24581 37275 24639 37281
rect 25332 37256 25360 37284
rect 20714 37244 20720 37256
rect 17819 37216 19104 37244
rect 19444 37216 20720 37244
rect 17819 37213 17831 37216
rect 17773 37207 17831 37213
rect 19444 37188 19472 37216
rect 20714 37204 20720 37216
rect 20772 37244 20778 37256
rect 21085 37247 21143 37253
rect 21085 37244 21097 37247
rect 20772 37216 21097 37244
rect 20772 37204 20778 37216
rect 21085 37213 21097 37216
rect 21131 37244 21143 37247
rect 21453 37247 21511 37253
rect 21453 37244 21465 37247
rect 21131 37216 21465 37244
rect 21131 37213 21143 37216
rect 21085 37207 21143 37213
rect 21453 37213 21465 37216
rect 21499 37213 21511 37247
rect 21453 37207 21511 37213
rect 22094 37204 22100 37256
rect 22152 37244 22158 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 22152 37216 22201 37244
rect 22152 37204 22158 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 25314 37204 25320 37256
rect 25372 37204 25378 37256
rect 16485 37179 16543 37185
rect 16485 37176 16497 37179
rect 11747 37148 13124 37176
rect 13188 37148 16497 37176
rect 11747 37145 11759 37148
rect 11701 37139 11759 37145
rect 6840 37080 8432 37108
rect 11241 37111 11299 37117
rect 11241 37077 11253 37111
rect 11287 37077 11299 37111
rect 11241 37071 11299 37077
rect 12621 37111 12679 37117
rect 12621 37077 12633 37111
rect 12667 37108 12679 37111
rect 12710 37108 12716 37120
rect 12667 37080 12716 37108
rect 12667 37077 12679 37080
rect 12621 37071 12679 37077
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 13096 37108 13124 37148
rect 16485 37145 16497 37148
rect 16531 37145 16543 37179
rect 17586 37176 17592 37188
rect 16485 37139 16543 37145
rect 17236 37148 17592 37176
rect 13906 37108 13912 37120
rect 13096 37080 13912 37108
rect 13906 37068 13912 37080
rect 13964 37068 13970 37120
rect 14090 37068 14096 37120
rect 14148 37108 14154 37120
rect 14185 37111 14243 37117
rect 14185 37108 14197 37111
rect 14148 37080 14197 37108
rect 14148 37068 14154 37080
rect 14185 37077 14197 37080
rect 14231 37077 14243 37111
rect 14185 37071 14243 37077
rect 14461 37111 14519 37117
rect 14461 37077 14473 37111
rect 14507 37108 14519 37111
rect 15102 37108 15108 37120
rect 14507 37080 15108 37108
rect 14507 37077 14519 37080
rect 14461 37071 14519 37077
rect 15102 37068 15108 37080
rect 15160 37068 15166 37120
rect 15194 37068 15200 37120
rect 15252 37108 15258 37120
rect 15289 37111 15347 37117
rect 15289 37108 15301 37111
rect 15252 37080 15301 37108
rect 15252 37068 15258 37080
rect 15289 37077 15301 37080
rect 15335 37077 15347 37111
rect 15289 37071 15347 37077
rect 15381 37111 15439 37117
rect 15381 37077 15393 37111
rect 15427 37108 15439 37111
rect 15562 37108 15568 37120
rect 15427 37080 15568 37108
rect 15427 37077 15439 37080
rect 15381 37071 15439 37077
rect 15562 37068 15568 37080
rect 15620 37068 15626 37120
rect 16117 37111 16175 37117
rect 16117 37077 16129 37111
rect 16163 37108 16175 37111
rect 17236 37108 17264 37148
rect 17586 37136 17592 37148
rect 17644 37136 17650 37188
rect 17681 37179 17739 37185
rect 17681 37145 17693 37179
rect 17727 37176 17739 37179
rect 17727 37148 19380 37176
rect 17727 37145 17739 37148
rect 17681 37139 17739 37145
rect 16163 37080 17264 37108
rect 16163 37077 16175 37080
rect 16117 37071 16175 37077
rect 18506 37068 18512 37120
rect 18564 37068 18570 37120
rect 19352 37108 19380 37148
rect 19426 37136 19432 37188
rect 19484 37136 19490 37188
rect 19794 37136 19800 37188
rect 19852 37176 19858 37188
rect 20165 37179 20223 37185
rect 20165 37176 20177 37179
rect 19852 37148 20177 37176
rect 19852 37136 19858 37148
rect 20165 37145 20177 37148
rect 20211 37145 20223 37179
rect 20165 37139 20223 37145
rect 20806 37136 20812 37188
rect 20864 37176 20870 37188
rect 20990 37176 20996 37188
rect 20864 37148 20996 37176
rect 20864 37136 20870 37148
rect 20990 37136 20996 37148
rect 21048 37176 21054 37188
rect 21048 37148 25176 37176
rect 21048 37136 21054 37148
rect 20070 37108 20076 37120
rect 19352 37080 20076 37108
rect 20070 37068 20076 37080
rect 20128 37068 20134 37120
rect 20714 37068 20720 37120
rect 20772 37108 20778 37120
rect 21082 37108 21088 37120
rect 20772 37080 21088 37108
rect 20772 37068 20778 37080
rect 21082 37068 21088 37080
rect 21140 37068 21146 37120
rect 23753 37111 23811 37117
rect 23753 37077 23765 37111
rect 23799 37108 23811 37111
rect 24762 37108 24768 37120
rect 23799 37080 24768 37108
rect 23799 37077 23811 37080
rect 23753 37071 23811 37077
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 25148 37117 25176 37148
rect 25133 37111 25191 37117
rect 25133 37077 25145 37111
rect 25179 37077 25191 37111
rect 25133 37071 25191 37077
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 5534 36904 5540 36916
rect 3988 36876 5540 36904
rect 3988 36777 4016 36876
rect 5534 36864 5540 36876
rect 5592 36904 5598 36916
rect 6546 36904 6552 36916
rect 5592 36876 6552 36904
rect 5592 36864 5598 36876
rect 6546 36864 6552 36876
rect 6604 36864 6610 36916
rect 7466 36864 7472 36916
rect 7524 36864 7530 36916
rect 7929 36907 7987 36913
rect 7929 36873 7941 36907
rect 7975 36904 7987 36907
rect 8478 36904 8484 36916
rect 7975 36876 8484 36904
rect 7975 36873 7987 36876
rect 7929 36867 7987 36873
rect 8478 36864 8484 36876
rect 8536 36864 8542 36916
rect 9030 36864 9036 36916
rect 9088 36864 9094 36916
rect 10778 36864 10784 36916
rect 10836 36904 10842 36916
rect 12161 36907 12219 36913
rect 12161 36904 12173 36907
rect 10836 36876 12173 36904
rect 10836 36864 10842 36876
rect 12161 36873 12173 36876
rect 12207 36873 12219 36907
rect 12161 36867 12219 36873
rect 12250 36864 12256 36916
rect 12308 36904 12314 36916
rect 12621 36907 12679 36913
rect 12621 36904 12633 36907
rect 12308 36876 12633 36904
rect 12308 36864 12314 36876
rect 12621 36873 12633 36876
rect 12667 36873 12679 36907
rect 12621 36867 12679 36873
rect 13722 36864 13728 36916
rect 13780 36904 13786 36916
rect 13817 36907 13875 36913
rect 13817 36904 13829 36907
rect 13780 36876 13829 36904
rect 13780 36864 13786 36876
rect 13817 36873 13829 36876
rect 13863 36873 13875 36907
rect 13817 36867 13875 36873
rect 14458 36864 14464 36916
rect 14516 36904 14522 36916
rect 15013 36907 15071 36913
rect 15013 36904 15025 36907
rect 14516 36876 15025 36904
rect 14516 36864 14522 36876
rect 15013 36873 15025 36876
rect 15059 36873 15071 36907
rect 15013 36867 15071 36873
rect 15378 36864 15384 36916
rect 15436 36904 15442 36916
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 15436 36876 15577 36904
rect 15436 36864 15442 36876
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 15565 36867 15623 36873
rect 15838 36864 15844 36916
rect 15896 36904 15902 36916
rect 16942 36904 16948 36916
rect 15896 36876 16948 36904
rect 15896 36864 15902 36876
rect 16942 36864 16948 36876
rect 17000 36864 17006 36916
rect 17037 36907 17095 36913
rect 17037 36873 17049 36907
rect 17083 36873 17095 36907
rect 17037 36867 17095 36873
rect 17405 36907 17463 36913
rect 17405 36873 17417 36907
rect 17451 36904 17463 36907
rect 18506 36904 18512 36916
rect 17451 36876 18512 36904
rect 17451 36873 17463 36876
rect 17405 36867 17463 36873
rect 6086 36836 6092 36848
rect 5474 36808 6092 36836
rect 6086 36796 6092 36808
rect 6144 36796 6150 36848
rect 10229 36839 10287 36845
rect 10229 36805 10241 36839
rect 10275 36836 10287 36839
rect 10410 36836 10416 36848
rect 10275 36808 10416 36836
rect 10275 36805 10287 36808
rect 10229 36799 10287 36805
rect 10410 36796 10416 36808
rect 10468 36836 10474 36848
rect 11517 36839 11575 36845
rect 11517 36836 11529 36839
rect 10468 36808 11529 36836
rect 10468 36796 10474 36808
rect 11517 36805 11529 36808
rect 11563 36805 11575 36839
rect 11517 36799 11575 36805
rect 12069 36839 12127 36845
rect 12069 36805 12081 36839
rect 12115 36836 12127 36839
rect 12529 36839 12587 36845
rect 12529 36836 12541 36839
rect 12115 36808 12541 36836
rect 12115 36805 12127 36808
rect 12069 36799 12127 36805
rect 12529 36805 12541 36808
rect 12575 36836 12587 36839
rect 12710 36836 12716 36848
rect 12575 36808 12716 36836
rect 12575 36805 12587 36808
rect 12529 36799 12587 36805
rect 3973 36771 4031 36777
rect 3973 36737 3985 36771
rect 4019 36737 4031 36771
rect 3973 36731 4031 36737
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36768 7895 36771
rect 9122 36768 9128 36780
rect 7883 36740 9128 36768
rect 7883 36737 7895 36740
rect 7837 36731 7895 36737
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 9306 36728 9312 36780
rect 9364 36768 9370 36780
rect 9401 36771 9459 36777
rect 9401 36768 9413 36771
rect 9364 36740 9413 36768
rect 9364 36728 9370 36740
rect 9401 36737 9413 36740
rect 9447 36737 9459 36771
rect 9401 36731 9459 36737
rect 9493 36771 9551 36777
rect 9493 36737 9505 36771
rect 9539 36768 9551 36771
rect 11054 36768 11060 36780
rect 9539 36740 11060 36768
rect 9539 36737 9551 36740
rect 9493 36731 9551 36737
rect 11054 36728 11060 36740
rect 11112 36728 11118 36780
rect 11532 36768 11560 36799
rect 12710 36796 12716 36808
rect 12768 36836 12774 36848
rect 13538 36836 13544 36848
rect 12768 36808 13544 36836
rect 12768 36796 12774 36808
rect 13538 36796 13544 36808
rect 13596 36796 13602 36848
rect 17052 36836 17080 36867
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 19886 36864 19892 36916
rect 19944 36904 19950 36916
rect 20349 36907 20407 36913
rect 20349 36904 20361 36907
rect 19944 36876 20361 36904
rect 19944 36864 19950 36876
rect 20349 36873 20361 36876
rect 20395 36873 20407 36907
rect 20349 36867 20407 36873
rect 20441 36907 20499 36913
rect 20441 36873 20453 36907
rect 20487 36904 20499 36907
rect 20530 36904 20536 36916
rect 20487 36876 20536 36904
rect 20487 36873 20499 36876
rect 20441 36867 20499 36873
rect 20530 36864 20536 36876
rect 20588 36904 20594 36916
rect 20993 36907 21051 36913
rect 20993 36904 21005 36907
rect 20588 36876 21005 36904
rect 20588 36864 20594 36876
rect 20993 36873 21005 36876
rect 21039 36873 21051 36907
rect 20993 36867 21051 36873
rect 22830 36864 22836 36916
rect 22888 36904 22894 36916
rect 23290 36904 23296 36916
rect 22888 36876 23296 36904
rect 22888 36864 22894 36876
rect 18782 36836 18788 36848
rect 17052 36808 18788 36836
rect 18782 36796 18788 36808
rect 18840 36796 18846 36848
rect 23124 36845 23152 36876
rect 23290 36864 23296 36876
rect 23348 36864 23354 36916
rect 23842 36864 23848 36916
rect 23900 36904 23906 36916
rect 24581 36907 24639 36913
rect 24581 36904 24593 36907
rect 23900 36876 24593 36904
rect 23900 36864 23906 36876
rect 24581 36873 24593 36876
rect 24627 36873 24639 36907
rect 24581 36867 24639 36873
rect 23109 36839 23167 36845
rect 23109 36805 23121 36839
rect 23155 36805 23167 36839
rect 24762 36836 24768 36848
rect 24334 36808 24768 36836
rect 23109 36799 23167 36805
rect 24762 36796 24768 36808
rect 24820 36796 24826 36848
rect 11532 36740 12434 36768
rect 4249 36703 4307 36709
rect 4249 36669 4261 36703
rect 4295 36700 4307 36703
rect 5442 36700 5448 36712
rect 4295 36672 5448 36700
rect 4295 36669 4307 36672
rect 4249 36663 4307 36669
rect 5442 36660 5448 36672
rect 5500 36700 5506 36712
rect 5721 36703 5779 36709
rect 5500 36672 5672 36700
rect 5500 36660 5506 36672
rect 5644 36632 5672 36672
rect 5721 36669 5733 36703
rect 5767 36700 5779 36703
rect 5810 36700 5816 36712
rect 5767 36672 5816 36700
rect 5767 36669 5779 36672
rect 5721 36663 5779 36669
rect 5810 36660 5816 36672
rect 5868 36660 5874 36712
rect 5994 36660 6000 36712
rect 6052 36700 6058 36712
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 6052 36672 8033 36700
rect 6052 36660 6058 36672
rect 8021 36669 8033 36672
rect 8067 36669 8079 36703
rect 8021 36663 8079 36669
rect 9582 36660 9588 36712
rect 9640 36660 9646 36712
rect 10962 36660 10968 36712
rect 11020 36660 11026 36712
rect 7834 36632 7840 36644
rect 5644 36604 7840 36632
rect 7834 36592 7840 36604
rect 7892 36592 7898 36644
rect 9490 36592 9496 36644
rect 9548 36632 9554 36644
rect 11793 36635 11851 36641
rect 11793 36632 11805 36635
rect 9548 36604 11805 36632
rect 9548 36592 9554 36604
rect 11793 36601 11805 36604
rect 11839 36632 11851 36635
rect 12250 36632 12256 36644
rect 11839 36604 12256 36632
rect 11839 36601 11851 36604
rect 11793 36595 11851 36601
rect 12250 36592 12256 36604
rect 12308 36592 12314 36644
rect 12406 36632 12434 36740
rect 12802 36728 12808 36780
rect 12860 36768 12866 36780
rect 13725 36771 13783 36777
rect 13725 36768 13737 36771
rect 12860 36740 13737 36768
rect 12860 36728 12866 36740
rect 13725 36737 13737 36740
rect 13771 36768 13783 36771
rect 14090 36768 14096 36780
rect 13771 36740 14096 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 14090 36728 14096 36740
rect 14148 36768 14154 36780
rect 14826 36768 14832 36780
rect 14148 36740 14832 36768
rect 14148 36728 14154 36740
rect 14826 36728 14832 36740
rect 14884 36728 14890 36780
rect 14921 36771 14979 36777
rect 14921 36737 14933 36771
rect 14967 36768 14979 36771
rect 14967 36740 15884 36768
rect 14967 36737 14979 36740
rect 14921 36731 14979 36737
rect 15856 36712 15884 36740
rect 16666 36728 16672 36780
rect 16724 36768 16730 36780
rect 17497 36771 17555 36777
rect 17497 36768 17509 36771
rect 16724 36740 17509 36768
rect 16724 36728 16730 36740
rect 17497 36737 17509 36740
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 19334 36728 19340 36780
rect 19392 36728 19398 36780
rect 22094 36728 22100 36780
rect 22152 36768 22158 36780
rect 22830 36768 22836 36780
rect 22152 36740 22836 36768
rect 22152 36728 22158 36740
rect 22830 36728 22836 36740
rect 22888 36728 22894 36780
rect 24394 36728 24400 36780
rect 24452 36768 24458 36780
rect 25314 36768 25320 36780
rect 24452 36740 25320 36768
rect 24452 36728 24458 36740
rect 25314 36728 25320 36740
rect 25372 36728 25378 36780
rect 12710 36660 12716 36712
rect 12768 36660 12774 36712
rect 13998 36660 14004 36712
rect 14056 36660 14062 36712
rect 15102 36660 15108 36712
rect 15160 36660 15166 36712
rect 15838 36660 15844 36712
rect 15896 36660 15902 36712
rect 17310 36660 17316 36712
rect 17368 36700 17374 36712
rect 17589 36703 17647 36709
rect 17589 36700 17601 36703
rect 17368 36672 17601 36700
rect 17368 36660 17374 36672
rect 17589 36669 17601 36672
rect 17635 36669 17647 36703
rect 17589 36663 17647 36669
rect 18782 36660 18788 36712
rect 18840 36700 18846 36712
rect 19242 36700 19248 36712
rect 18840 36672 19248 36700
rect 18840 36660 18846 36672
rect 19242 36660 19248 36672
rect 19300 36660 19306 36712
rect 19352 36700 19380 36728
rect 20533 36703 20591 36709
rect 20533 36700 20545 36703
rect 19352 36672 20545 36700
rect 20533 36669 20545 36672
rect 20579 36669 20591 36703
rect 20533 36663 20591 36669
rect 22370 36660 22376 36712
rect 22428 36700 22434 36712
rect 25130 36700 25136 36712
rect 22428 36672 25136 36700
rect 22428 36660 22434 36672
rect 25130 36660 25136 36672
rect 25188 36660 25194 36712
rect 16022 36632 16028 36644
rect 12406 36604 16028 36632
rect 16022 36592 16028 36604
rect 16080 36632 16086 36644
rect 19337 36635 19395 36641
rect 19337 36632 19349 36635
rect 16080 36604 19349 36632
rect 16080 36592 16086 36604
rect 19337 36601 19349 36604
rect 19383 36632 19395 36635
rect 19426 36632 19432 36644
rect 19383 36604 19432 36632
rect 19383 36601 19395 36604
rect 19337 36595 19395 36601
rect 19426 36592 19432 36604
rect 19484 36592 19490 36644
rect 6086 36524 6092 36576
rect 6144 36524 6150 36576
rect 8754 36524 8760 36576
rect 8812 36564 8818 36576
rect 9398 36564 9404 36576
rect 8812 36536 9404 36564
rect 8812 36524 8818 36536
rect 9398 36524 9404 36536
rect 9456 36524 9462 36576
rect 13357 36567 13415 36573
rect 13357 36533 13369 36567
rect 13403 36564 13415 36567
rect 14458 36564 14464 36576
rect 13403 36536 14464 36564
rect 13403 36533 13415 36536
rect 13357 36527 13415 36533
rect 14458 36524 14464 36536
rect 14516 36524 14522 36576
rect 14550 36524 14556 36576
rect 14608 36524 14614 36576
rect 17218 36524 17224 36576
rect 17276 36564 17282 36576
rect 19981 36567 20039 36573
rect 19981 36564 19993 36567
rect 17276 36536 19993 36564
rect 17276 36524 17282 36536
rect 19981 36533 19993 36536
rect 20027 36533 20039 36567
rect 19981 36527 20039 36533
rect 20070 36524 20076 36576
rect 20128 36564 20134 36576
rect 25133 36567 25191 36573
rect 25133 36564 25145 36567
rect 20128 36536 25145 36564
rect 20128 36524 20134 36536
rect 25133 36533 25145 36536
rect 25179 36533 25191 36567
rect 25133 36527 25191 36533
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 7650 36320 7656 36372
rect 7708 36320 7714 36372
rect 8938 36320 8944 36372
rect 8996 36360 9002 36372
rect 9125 36363 9183 36369
rect 9125 36360 9137 36363
rect 8996 36332 9137 36360
rect 8996 36320 9002 36332
rect 9125 36329 9137 36332
rect 9171 36329 9183 36363
rect 9125 36323 9183 36329
rect 9766 36320 9772 36372
rect 9824 36360 9830 36372
rect 12161 36363 12219 36369
rect 12161 36360 12173 36363
rect 9824 36332 12173 36360
rect 9824 36320 9830 36332
rect 12161 36329 12173 36332
rect 12207 36360 12219 36363
rect 12713 36363 12771 36369
rect 12207 36332 12664 36360
rect 12207 36329 12219 36332
rect 12161 36323 12219 36329
rect 12636 36292 12664 36332
rect 12713 36329 12725 36363
rect 12759 36360 12771 36363
rect 13354 36360 13360 36372
rect 12759 36332 13360 36360
rect 12759 36329 12771 36332
rect 12713 36323 12771 36329
rect 13354 36320 13360 36332
rect 13412 36320 13418 36372
rect 14277 36363 14335 36369
rect 14277 36329 14289 36363
rect 14323 36360 14335 36363
rect 15470 36360 15476 36372
rect 14323 36332 15476 36360
rect 14323 36329 14335 36332
rect 14277 36323 14335 36329
rect 15470 36320 15476 36332
rect 15528 36320 15534 36372
rect 19429 36363 19487 36369
rect 19429 36329 19441 36363
rect 19475 36360 19487 36363
rect 19518 36360 19524 36372
rect 19475 36332 19524 36360
rect 19475 36329 19487 36332
rect 19429 36323 19487 36329
rect 19518 36320 19524 36332
rect 19576 36320 19582 36372
rect 21726 36320 21732 36372
rect 21784 36360 21790 36372
rect 25133 36363 25191 36369
rect 25133 36360 25145 36363
rect 21784 36332 25145 36360
rect 21784 36320 21790 36332
rect 25133 36329 25145 36332
rect 25179 36329 25191 36363
rect 25133 36323 25191 36329
rect 13078 36292 13084 36304
rect 12636 36264 13084 36292
rect 13078 36252 13084 36264
rect 13136 36252 13142 36304
rect 16117 36295 16175 36301
rect 16117 36261 16129 36295
rect 16163 36292 16175 36295
rect 18966 36292 18972 36304
rect 16163 36264 18972 36292
rect 16163 36261 16175 36264
rect 16117 36255 16175 36261
rect 18966 36252 18972 36264
rect 19024 36252 19030 36304
rect 23293 36295 23351 36301
rect 23293 36261 23305 36295
rect 23339 36292 23351 36295
rect 24394 36292 24400 36304
rect 23339 36264 24400 36292
rect 23339 36261 23351 36264
rect 23293 36255 23351 36261
rect 24394 36252 24400 36264
rect 24452 36252 24458 36304
rect 7558 36184 7564 36236
rect 7616 36224 7622 36236
rect 8205 36227 8263 36233
rect 8205 36224 8217 36227
rect 7616 36196 8217 36224
rect 7616 36184 7622 36196
rect 8205 36193 8217 36196
rect 8251 36193 8263 36227
rect 9677 36227 9735 36233
rect 9677 36224 9689 36227
rect 8205 36187 8263 36193
rect 8312 36196 9689 36224
rect 1762 36116 1768 36168
rect 1820 36156 1826 36168
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 1820 36128 2053 36156
rect 1820 36116 1826 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 7834 36116 7840 36168
rect 7892 36156 7898 36168
rect 8312 36156 8340 36196
rect 9677 36193 9689 36196
rect 9723 36193 9735 36227
rect 9677 36187 9735 36193
rect 12434 36184 12440 36236
rect 12492 36224 12498 36236
rect 13173 36227 13231 36233
rect 13173 36224 13185 36227
rect 12492 36196 13185 36224
rect 12492 36184 12498 36196
rect 13173 36193 13185 36196
rect 13219 36193 13231 36227
rect 13173 36187 13231 36193
rect 13354 36184 13360 36236
rect 13412 36184 13418 36236
rect 13538 36184 13544 36236
rect 13596 36224 13602 36236
rect 14921 36227 14979 36233
rect 13596 36196 14872 36224
rect 13596 36184 13602 36196
rect 7892 36128 8340 36156
rect 9585 36159 9643 36165
rect 7892 36116 7898 36128
rect 9585 36125 9597 36159
rect 9631 36156 9643 36159
rect 11790 36156 11796 36168
rect 9631 36128 11796 36156
rect 9631 36125 9643 36128
rect 9585 36119 9643 36125
rect 11790 36116 11796 36128
rect 11848 36116 11854 36168
rect 12066 36116 12072 36168
rect 12124 36156 12130 36168
rect 13998 36156 14004 36168
rect 12124 36128 14004 36156
rect 12124 36116 12130 36128
rect 13998 36116 14004 36128
rect 14056 36116 14062 36168
rect 8113 36091 8171 36097
rect 8113 36057 8125 36091
rect 8159 36088 8171 36091
rect 10318 36088 10324 36100
rect 8159 36060 10324 36088
rect 8159 36057 8171 36060
rect 8113 36051 8171 36057
rect 10318 36048 10324 36060
rect 10376 36048 10382 36100
rect 10686 36048 10692 36100
rect 10744 36088 10750 36100
rect 12250 36088 12256 36100
rect 10744 36060 12256 36088
rect 10744 36048 10750 36060
rect 12250 36048 12256 36060
rect 12308 36088 12314 36100
rect 13817 36091 13875 36097
rect 13817 36088 13829 36091
rect 12308 36060 12434 36088
rect 12308 36048 12314 36060
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 4154 36020 4160 36032
rect 1627 35992 4160 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 4154 35980 4160 35992
rect 4212 35980 4218 36032
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 8021 36023 8079 36029
rect 8021 36020 8033 36023
rect 7524 35992 8033 36020
rect 7524 35980 7530 35992
rect 8021 35989 8033 35992
rect 8067 35989 8079 36023
rect 8021 35983 8079 35989
rect 9493 36023 9551 36029
rect 9493 35989 9505 36023
rect 9539 36020 9551 36023
rect 11238 36020 11244 36032
rect 9539 35992 11244 36020
rect 9539 35989 9551 35992
rect 9493 35983 9551 35989
rect 11238 35980 11244 35992
rect 11296 35980 11302 36032
rect 12406 36020 12434 36060
rect 12544 36060 13829 36088
rect 12544 36020 12572 36060
rect 13817 36057 13829 36060
rect 13863 36088 13875 36091
rect 14737 36091 14795 36097
rect 14737 36088 14749 36091
rect 13863 36060 14749 36088
rect 13863 36057 13875 36060
rect 13817 36051 13875 36057
rect 14737 36057 14749 36060
rect 14783 36057 14795 36091
rect 14737 36051 14795 36057
rect 12406 35992 12572 36020
rect 13078 35980 13084 36032
rect 13136 36020 13142 36032
rect 13630 36020 13636 36032
rect 13136 35992 13636 36020
rect 13136 35980 13142 35992
rect 13630 35980 13636 35992
rect 13688 35980 13694 36032
rect 14642 35980 14648 36032
rect 14700 35980 14706 36032
rect 14844 36020 14872 36196
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 15010 36224 15016 36236
rect 14967 36196 15016 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 15010 36184 15016 36196
rect 15068 36184 15074 36236
rect 15746 36184 15752 36236
rect 15804 36184 15810 36236
rect 16482 36184 16488 36236
rect 16540 36224 16546 36236
rect 16669 36227 16727 36233
rect 16669 36224 16681 36227
rect 16540 36196 16681 36224
rect 16540 36184 16546 36196
rect 16669 36193 16681 36196
rect 16715 36193 16727 36227
rect 16669 36187 16727 36193
rect 16942 36184 16948 36236
rect 17000 36224 17006 36236
rect 19061 36227 19119 36233
rect 19061 36224 19073 36227
rect 17000 36196 19073 36224
rect 17000 36184 17006 36196
rect 19061 36193 19073 36196
rect 19107 36224 19119 36227
rect 19981 36227 20039 36233
rect 19981 36224 19993 36227
rect 19107 36196 19993 36224
rect 19107 36193 19119 36196
rect 19061 36187 19119 36193
rect 19981 36193 19993 36196
rect 20027 36193 20039 36227
rect 19981 36187 20039 36193
rect 21266 36184 21272 36236
rect 21324 36184 21330 36236
rect 21453 36227 21511 36233
rect 21453 36193 21465 36227
rect 21499 36224 21511 36227
rect 21634 36224 21640 36236
rect 21499 36196 21640 36224
rect 21499 36193 21511 36196
rect 21453 36187 21511 36193
rect 21634 36184 21640 36196
rect 21692 36184 21698 36236
rect 23750 36184 23756 36236
rect 23808 36184 23814 36236
rect 23937 36227 23995 36233
rect 23937 36193 23949 36227
rect 23983 36224 23995 36227
rect 24486 36224 24492 36236
rect 23983 36196 24492 36224
rect 23983 36193 23995 36196
rect 23937 36187 23995 36193
rect 24486 36184 24492 36196
rect 24544 36184 24550 36236
rect 15764 36156 15792 36184
rect 16577 36159 16635 36165
rect 16577 36156 16589 36159
rect 15764 36128 16589 36156
rect 16577 36125 16589 36128
rect 16623 36125 16635 36159
rect 21910 36156 21916 36168
rect 16577 36119 16635 36125
rect 17420 36128 21916 36156
rect 16485 36091 16543 36097
rect 16485 36057 16497 36091
rect 16531 36088 16543 36091
rect 17313 36091 17371 36097
rect 17313 36088 17325 36091
rect 16531 36060 17325 36088
rect 16531 36057 16543 36060
rect 16485 36051 16543 36057
rect 17313 36057 17325 36060
rect 17359 36057 17371 36091
rect 17313 36051 17371 36057
rect 17420 36020 17448 36128
rect 21910 36116 21916 36128
rect 21968 36156 21974 36168
rect 24578 36156 24584 36168
rect 21968 36128 24584 36156
rect 21968 36116 21974 36128
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 19889 36091 19947 36097
rect 19889 36057 19901 36091
rect 19935 36088 19947 36091
rect 19935 36060 22094 36088
rect 19935 36057 19947 36060
rect 19889 36051 19947 36057
rect 14844 35992 17448 36020
rect 19797 36023 19855 36029
rect 19797 35989 19809 36023
rect 19843 36020 19855 36023
rect 20530 36020 20536 36032
rect 19843 35992 20536 36020
rect 19843 35989 19855 35992
rect 19797 35983 19855 35989
rect 20530 35980 20536 35992
rect 20588 35980 20594 36032
rect 20806 35980 20812 36032
rect 20864 35980 20870 36032
rect 21177 36023 21235 36029
rect 21177 35989 21189 36023
rect 21223 36020 21235 36023
rect 21450 36020 21456 36032
rect 21223 35992 21456 36020
rect 21223 35989 21235 35992
rect 21177 35983 21235 35989
rect 21450 35980 21456 35992
rect 21508 35980 21514 36032
rect 22066 36020 22094 36060
rect 22370 36020 22376 36032
rect 22066 35992 22376 36020
rect 22370 35980 22376 35992
rect 22428 35980 22434 36032
rect 23658 35980 23664 36032
rect 23716 35980 23722 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 5534 35816 5540 35828
rect 4264 35788 5540 35816
rect 4264 35689 4292 35788
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 5994 35776 6000 35828
rect 6052 35776 6058 35828
rect 13446 35816 13452 35828
rect 10244 35788 13452 35816
rect 10137 35751 10195 35757
rect 10137 35748 10149 35751
rect 9614 35720 10149 35748
rect 4249 35683 4307 35689
rect 4249 35649 4261 35683
rect 4295 35649 4307 35683
rect 6086 35680 6092 35692
rect 5658 35652 6092 35680
rect 4249 35643 4307 35649
rect 6086 35640 6092 35652
rect 6144 35680 6150 35692
rect 6144 35652 6500 35680
rect 6144 35640 6150 35652
rect 4525 35615 4583 35621
rect 4525 35581 4537 35615
rect 4571 35612 4583 35615
rect 5810 35612 5816 35624
rect 4571 35584 5816 35612
rect 4571 35581 4583 35584
rect 4525 35575 4583 35581
rect 5810 35572 5816 35584
rect 5868 35572 5874 35624
rect 6472 35485 6500 35652
rect 8113 35615 8171 35621
rect 8113 35581 8125 35615
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 8389 35615 8447 35621
rect 8389 35581 8401 35615
rect 8435 35612 8447 35615
rect 9582 35612 9588 35624
rect 8435 35584 9588 35612
rect 8435 35581 8447 35584
rect 8389 35575 8447 35581
rect 6457 35479 6515 35485
rect 6457 35445 6469 35479
rect 6503 35476 6515 35479
rect 7650 35476 7656 35488
rect 6503 35448 7656 35476
rect 6503 35445 6515 35448
rect 6457 35439 6515 35445
rect 7650 35436 7656 35448
rect 7708 35436 7714 35488
rect 8128 35476 8156 35575
rect 9582 35572 9588 35584
rect 9640 35572 9646 35624
rect 8846 35476 8852 35488
rect 8128 35448 8852 35476
rect 8846 35436 8852 35448
rect 8904 35436 8910 35488
rect 9582 35436 9588 35488
rect 9640 35476 9646 35488
rect 9692 35476 9720 35720
rect 10137 35717 10149 35720
rect 10183 35717 10195 35751
rect 10137 35711 10195 35717
rect 10244 35680 10272 35788
rect 13446 35776 13452 35788
rect 13504 35776 13510 35828
rect 14461 35819 14519 35825
rect 14461 35785 14473 35819
rect 14507 35816 14519 35819
rect 14642 35816 14648 35828
rect 14507 35788 14648 35816
rect 14507 35785 14519 35788
rect 14461 35779 14519 35785
rect 14642 35776 14648 35788
rect 14700 35776 14706 35828
rect 15010 35776 15016 35828
rect 15068 35816 15074 35828
rect 17126 35816 17132 35828
rect 15068 35788 17132 35816
rect 15068 35776 15074 35788
rect 17126 35776 17132 35788
rect 17184 35776 17190 35828
rect 17678 35776 17684 35828
rect 17736 35816 17742 35828
rect 17736 35788 17908 35816
rect 17736 35776 17742 35788
rect 11882 35708 11888 35760
rect 11940 35748 11946 35760
rect 14001 35751 14059 35757
rect 11940 35720 12466 35748
rect 11940 35708 11946 35720
rect 14001 35717 14013 35751
rect 14047 35748 14059 35751
rect 17770 35748 17776 35760
rect 14047 35720 17776 35748
rect 14047 35717 14059 35720
rect 14001 35711 14059 35717
rect 9876 35652 10272 35680
rect 9640 35448 9720 35476
rect 9640 35436 9646 35448
rect 9766 35436 9772 35488
rect 9824 35476 9830 35488
rect 9876 35485 9904 35652
rect 13354 35640 13360 35692
rect 13412 35680 13418 35692
rect 14016 35680 14044 35711
rect 17770 35708 17776 35720
rect 17828 35708 17834 35760
rect 17880 35757 17908 35788
rect 19242 35776 19248 35828
rect 19300 35776 19306 35828
rect 19337 35819 19395 35825
rect 19337 35785 19349 35819
rect 19383 35816 19395 35819
rect 21542 35816 21548 35828
rect 19383 35788 21548 35816
rect 19383 35785 19395 35788
rect 19337 35779 19395 35785
rect 21542 35776 21548 35788
rect 21600 35776 21606 35828
rect 23290 35776 23296 35828
rect 23348 35816 23354 35828
rect 24857 35819 24915 35825
rect 24857 35816 24869 35819
rect 23348 35788 24869 35816
rect 23348 35776 23354 35788
rect 24857 35785 24869 35788
rect 24903 35785 24915 35819
rect 24857 35779 24915 35785
rect 17865 35751 17923 35757
rect 17865 35717 17877 35751
rect 17911 35717 17923 35751
rect 19260 35748 19288 35776
rect 19260 35720 20392 35748
rect 17865 35711 17923 35717
rect 13412 35652 14044 35680
rect 18892 35652 18998 35680
rect 13412 35640 13418 35652
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11020 35584 11713 35612
rect 11020 35572 11026 35584
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11701 35575 11759 35581
rect 11977 35615 12035 35621
rect 11977 35581 11989 35615
rect 12023 35612 12035 35615
rect 13814 35612 13820 35624
rect 12023 35584 13820 35612
rect 12023 35581 12035 35584
rect 11977 35575 12035 35581
rect 13814 35572 13820 35584
rect 13872 35572 13878 35624
rect 17589 35615 17647 35621
rect 17589 35581 17601 35615
rect 17635 35612 17647 35615
rect 17635 35584 17724 35612
rect 17635 35581 17647 35584
rect 17589 35575 17647 35581
rect 13449 35547 13507 35553
rect 13449 35513 13461 35547
rect 13495 35544 13507 35547
rect 13538 35544 13544 35556
rect 13495 35516 13544 35544
rect 13495 35513 13507 35516
rect 13449 35507 13507 35513
rect 9861 35479 9919 35485
rect 9861 35476 9873 35479
rect 9824 35448 9873 35476
rect 9824 35436 9830 35448
rect 9861 35445 9873 35448
rect 9907 35445 9919 35479
rect 9861 35439 9919 35445
rect 12526 35436 12532 35488
rect 12584 35476 12590 35488
rect 13464 35476 13492 35507
rect 13538 35504 13544 35516
rect 13596 35504 13602 35556
rect 12584 35448 13492 35476
rect 12584 35436 12590 35448
rect 13722 35436 13728 35488
rect 13780 35436 13786 35488
rect 15930 35436 15936 35488
rect 15988 35476 15994 35488
rect 17696 35476 17724 35584
rect 18892 35544 18920 35652
rect 19242 35640 19248 35692
rect 19300 35680 19306 35692
rect 20165 35683 20223 35689
rect 20165 35680 20177 35683
rect 19300 35652 20177 35680
rect 19300 35640 19306 35652
rect 20088 35544 20116 35652
rect 20165 35649 20177 35652
rect 20211 35649 20223 35683
rect 20165 35643 20223 35649
rect 20254 35572 20260 35624
rect 20312 35572 20318 35624
rect 20364 35621 20392 35720
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 22830 35680 22836 35692
rect 22244 35652 22836 35680
rect 22244 35640 22250 35652
rect 22830 35640 22836 35652
rect 22888 35680 22894 35692
rect 23109 35683 23167 35689
rect 23109 35680 23121 35683
rect 22888 35652 23121 35680
rect 22888 35640 22894 35652
rect 23109 35649 23121 35652
rect 23155 35649 23167 35683
rect 23109 35643 23167 35649
rect 24486 35640 24492 35692
rect 24544 35640 24550 35692
rect 20349 35615 20407 35621
rect 20349 35581 20361 35615
rect 20395 35581 20407 35615
rect 20349 35575 20407 35581
rect 22462 35572 22468 35624
rect 22520 35572 22526 35624
rect 23382 35572 23388 35624
rect 23440 35572 23446 35624
rect 18892 35516 20024 35544
rect 20088 35516 22094 35544
rect 18322 35476 18328 35488
rect 15988 35448 18328 35476
rect 15988 35436 15994 35448
rect 18322 35436 18328 35448
rect 18380 35476 18386 35488
rect 19702 35476 19708 35488
rect 18380 35448 19708 35476
rect 18380 35436 18386 35448
rect 19702 35436 19708 35448
rect 19760 35436 19766 35488
rect 19794 35436 19800 35488
rect 19852 35436 19858 35488
rect 19996 35476 20024 35516
rect 20898 35476 20904 35488
rect 19996 35448 20904 35476
rect 20898 35436 20904 35448
rect 20956 35436 20962 35488
rect 22066 35476 22094 35516
rect 23934 35476 23940 35488
rect 22066 35448 23940 35476
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 24486 35436 24492 35488
rect 24544 35476 24550 35488
rect 24762 35476 24768 35488
rect 24544 35448 24768 35476
rect 24544 35436 24550 35448
rect 24762 35436 24768 35448
rect 24820 35476 24826 35488
rect 25225 35479 25283 35485
rect 25225 35476 25237 35479
rect 24820 35448 25237 35476
rect 24820 35436 24826 35448
rect 25225 35445 25237 35448
rect 25271 35445 25283 35479
rect 25225 35439 25283 35445
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 9309 35275 9367 35281
rect 9309 35272 9321 35275
rect 7432 35244 9321 35272
rect 7432 35232 7438 35244
rect 9309 35241 9321 35244
rect 9355 35241 9367 35275
rect 9309 35235 9367 35241
rect 11054 35232 11060 35284
rect 11112 35272 11118 35284
rect 12989 35275 13047 35281
rect 12989 35272 13001 35275
rect 11112 35244 13001 35272
rect 11112 35232 11118 35244
rect 12989 35241 13001 35244
rect 13035 35241 13047 35275
rect 12989 35235 13047 35241
rect 16114 35232 16120 35284
rect 16172 35272 16178 35284
rect 17129 35275 17187 35281
rect 17129 35272 17141 35275
rect 16172 35244 17141 35272
rect 16172 35232 16178 35244
rect 17129 35241 17141 35244
rect 17175 35241 17187 35275
rect 17129 35235 17187 35241
rect 19058 35232 19064 35284
rect 19116 35272 19122 35284
rect 21174 35272 21180 35284
rect 19116 35244 21180 35272
rect 19116 35232 19122 35244
rect 21174 35232 21180 35244
rect 21232 35272 21238 35284
rect 21545 35275 21603 35281
rect 21545 35272 21557 35275
rect 21232 35244 21557 35272
rect 21232 35232 21238 35244
rect 21545 35241 21557 35244
rect 21591 35241 21603 35275
rect 21545 35235 21603 35241
rect 7834 35164 7840 35216
rect 7892 35164 7898 35216
rect 8570 35164 8576 35216
rect 8628 35204 8634 35216
rect 8628 35176 9904 35204
rect 8628 35164 8634 35176
rect 5534 35096 5540 35148
rect 5592 35136 5598 35148
rect 6086 35136 6092 35148
rect 5592 35108 6092 35136
rect 5592 35096 5598 35108
rect 6086 35096 6092 35108
rect 6144 35096 6150 35148
rect 6365 35139 6423 35145
rect 6365 35105 6377 35139
rect 6411 35136 6423 35139
rect 9766 35136 9772 35148
rect 6411 35108 9772 35136
rect 6411 35105 6423 35108
rect 6365 35099 6423 35105
rect 9766 35096 9772 35108
rect 9824 35096 9830 35148
rect 9876 35145 9904 35176
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 19150 35204 19156 35216
rect 16724 35176 19156 35204
rect 16724 35164 16730 35176
rect 19150 35164 19156 35176
rect 19208 35164 19214 35216
rect 9861 35139 9919 35145
rect 9861 35105 9873 35139
rect 9907 35105 9919 35139
rect 9861 35099 9919 35105
rect 11054 35096 11060 35148
rect 11112 35136 11118 35148
rect 13541 35139 13599 35145
rect 13541 35136 13553 35139
rect 11112 35108 13553 35136
rect 11112 35096 11118 35108
rect 13541 35105 13553 35108
rect 13587 35105 13599 35139
rect 13541 35099 13599 35105
rect 15381 35139 15439 35145
rect 15381 35105 15393 35139
rect 15427 35136 15439 35139
rect 15746 35136 15752 35148
rect 15427 35108 15752 35136
rect 15427 35105 15439 35108
rect 15381 35099 15439 35105
rect 15746 35096 15752 35108
rect 15804 35096 15810 35148
rect 16114 35096 16120 35148
rect 16172 35136 16178 35148
rect 17405 35139 17463 35145
rect 17405 35136 17417 35139
rect 16172 35108 17417 35136
rect 16172 35096 16178 35108
rect 17405 35105 17417 35108
rect 17451 35105 17463 35139
rect 17405 35099 17463 35105
rect 19429 35139 19487 35145
rect 19429 35105 19441 35139
rect 19475 35136 19487 35139
rect 19702 35136 19708 35148
rect 19475 35108 19708 35136
rect 19475 35105 19487 35108
rect 19429 35099 19487 35105
rect 19702 35096 19708 35108
rect 19760 35096 19766 35148
rect 20254 35096 20260 35148
rect 20312 35136 20318 35148
rect 20714 35136 20720 35148
rect 20312 35108 20720 35136
rect 20312 35096 20318 35108
rect 20714 35096 20720 35108
rect 20772 35096 20778 35148
rect 20898 35096 20904 35148
rect 20956 35096 20962 35148
rect 21177 35139 21235 35145
rect 21177 35105 21189 35139
rect 21223 35136 21235 35139
rect 21634 35136 21640 35148
rect 21223 35108 21640 35136
rect 21223 35105 21235 35108
rect 21177 35099 21235 35105
rect 21634 35096 21640 35108
rect 21692 35096 21698 35148
rect 21821 35139 21879 35145
rect 21821 35105 21833 35139
rect 21867 35136 21879 35139
rect 21867 35108 23796 35136
rect 21867 35105 21879 35108
rect 21821 35099 21879 35105
rect 8294 35028 8300 35080
rect 8352 35068 8358 35080
rect 12710 35068 12716 35080
rect 8352 35040 12716 35068
rect 8352 35028 8358 35040
rect 12710 35028 12716 35040
rect 12768 35028 12774 35080
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35068 13507 35071
rect 14550 35068 14556 35080
rect 13495 35040 14556 35068
rect 13495 35037 13507 35040
rect 13449 35031 13507 35037
rect 14550 35028 14556 35040
rect 14608 35028 14614 35080
rect 20916 35068 20944 35096
rect 21836 35068 21864 35099
rect 20838 35040 21864 35068
rect 22186 35028 22192 35080
rect 22244 35068 22250 35080
rect 22281 35071 22339 35077
rect 22281 35068 22293 35071
rect 22244 35040 22293 35068
rect 22244 35028 22250 35040
rect 22281 35037 22293 35040
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 7650 35000 7656 35012
rect 7590 34972 7656 35000
rect 7650 34960 7656 34972
rect 7708 35000 7714 35012
rect 7708 34972 7880 35000
rect 7708 34960 7714 34972
rect 7852 34944 7880 34972
rect 8662 34960 8668 35012
rect 8720 35000 8726 35012
rect 9677 35003 9735 35009
rect 9677 35000 9689 35003
rect 8720 34972 9689 35000
rect 8720 34960 8726 34972
rect 9677 34969 9689 34972
rect 9723 34969 9735 35003
rect 9677 34963 9735 34969
rect 9769 35003 9827 35009
rect 9769 34969 9781 35003
rect 9815 35000 9827 35003
rect 14274 35000 14280 35012
rect 9815 34972 14280 35000
rect 9815 34969 9827 34972
rect 9769 34963 9827 34969
rect 14274 34960 14280 34972
rect 14332 34960 14338 35012
rect 15657 35003 15715 35009
rect 15657 34969 15669 35003
rect 15703 34969 15715 35003
rect 15657 34963 15715 34969
rect 7834 34892 7840 34944
rect 7892 34932 7898 34944
rect 8113 34935 8171 34941
rect 8113 34932 8125 34935
rect 7892 34904 8125 34932
rect 7892 34892 7898 34904
rect 8113 34901 8125 34904
rect 8159 34901 8171 34935
rect 8113 34895 8171 34901
rect 13354 34892 13360 34944
rect 13412 34892 13418 34944
rect 15672 34932 15700 34963
rect 16114 34960 16120 35012
rect 16172 34960 16178 35012
rect 19150 35000 19156 35012
rect 17052 34972 19156 35000
rect 17052 34932 17080 34972
rect 19150 34960 19156 34972
rect 19208 34960 19214 35012
rect 19702 34960 19708 35012
rect 19760 35000 19766 35012
rect 19978 35000 19984 35012
rect 19760 34972 19984 35000
rect 19760 34960 19766 34972
rect 19978 34960 19984 34972
rect 20036 34960 20042 35012
rect 22554 34960 22560 35012
rect 22612 34960 22618 35012
rect 23768 35000 23796 35108
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 23768 34986 24532 35000
rect 23782 34972 24532 34986
rect 24504 34944 24532 34972
rect 15672 34904 17080 34932
rect 23382 34892 23388 34944
rect 23440 34932 23446 34944
rect 24029 34935 24087 34941
rect 24029 34932 24041 34935
rect 23440 34904 24041 34932
rect 23440 34892 23446 34904
rect 24029 34901 24041 34904
rect 24075 34901 24087 34935
rect 24029 34895 24087 34901
rect 24486 34892 24492 34944
rect 24544 34892 24550 34944
rect 24762 34892 24768 34944
rect 24820 34932 24826 34944
rect 25133 34935 25191 34941
rect 25133 34932 25145 34935
rect 24820 34904 25145 34932
rect 24820 34892 24826 34904
rect 25133 34901 25145 34904
rect 25179 34901 25191 34935
rect 25133 34895 25191 34901
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 7098 34688 7104 34740
rect 7156 34728 7162 34740
rect 8294 34728 8300 34740
rect 7156 34700 8300 34728
rect 7156 34688 7162 34700
rect 8294 34688 8300 34700
rect 8352 34688 8358 34740
rect 9490 34688 9496 34740
rect 9548 34728 9554 34740
rect 10597 34731 10655 34737
rect 10597 34728 10609 34731
rect 9548 34700 10609 34728
rect 9548 34688 9554 34700
rect 10597 34697 10609 34700
rect 10643 34697 10655 34731
rect 13722 34728 13728 34740
rect 10597 34691 10655 34697
rect 12406 34700 13728 34728
rect 5994 34620 6000 34672
rect 6052 34660 6058 34672
rect 6825 34663 6883 34669
rect 6825 34660 6837 34663
rect 6052 34632 6837 34660
rect 6052 34620 6058 34632
rect 6825 34629 6837 34632
rect 6871 34629 6883 34663
rect 6825 34623 6883 34629
rect 9582 34620 9588 34672
rect 9640 34620 9646 34672
rect 11882 34620 11888 34672
rect 11940 34660 11946 34672
rect 12406 34660 12434 34700
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 14182 34688 14188 34740
rect 14240 34728 14246 34740
rect 15565 34731 15623 34737
rect 15565 34728 15577 34731
rect 14240 34700 15577 34728
rect 14240 34688 14246 34700
rect 15565 34697 15577 34700
rect 15611 34697 15623 34731
rect 15565 34691 15623 34697
rect 15933 34731 15991 34737
rect 15933 34697 15945 34731
rect 15979 34728 15991 34731
rect 19794 34728 19800 34740
rect 15979 34700 19800 34728
rect 15979 34697 15991 34700
rect 15933 34691 15991 34697
rect 19794 34688 19800 34700
rect 19852 34688 19858 34740
rect 20990 34688 20996 34740
rect 21048 34728 21054 34740
rect 21085 34731 21143 34737
rect 21085 34728 21097 34731
rect 21048 34700 21097 34728
rect 21048 34688 21054 34700
rect 21085 34697 21097 34700
rect 21131 34697 21143 34731
rect 21085 34691 21143 34697
rect 21174 34688 21180 34740
rect 21232 34688 21238 34740
rect 22370 34688 22376 34740
rect 22428 34688 22434 34740
rect 22462 34688 22468 34740
rect 22520 34728 22526 34740
rect 23569 34731 23627 34737
rect 23569 34728 23581 34731
rect 22520 34700 23581 34728
rect 22520 34688 22526 34700
rect 23569 34697 23581 34700
rect 23615 34697 23627 34731
rect 23569 34691 23627 34697
rect 24397 34731 24455 34737
rect 24397 34697 24409 34731
rect 24443 34728 24455 34731
rect 24670 34728 24676 34740
rect 24443 34700 24676 34728
rect 24443 34697 24455 34700
rect 24397 34691 24455 34697
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25133 34731 25191 34737
rect 25133 34697 25145 34731
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 13740 34660 13768 34688
rect 14366 34660 14372 34672
rect 11940 34632 12466 34660
rect 13740 34632 14372 34660
rect 11940 34620 11946 34632
rect 14366 34620 14372 34632
rect 14424 34620 14430 34672
rect 15194 34620 15200 34672
rect 15252 34660 15258 34672
rect 15746 34660 15752 34672
rect 15252 34632 15752 34660
rect 15252 34620 15258 34632
rect 15746 34620 15752 34632
rect 15804 34620 15810 34672
rect 16025 34663 16083 34669
rect 16025 34629 16037 34663
rect 16071 34660 16083 34663
rect 18414 34660 18420 34672
rect 16071 34632 18420 34660
rect 16071 34629 16083 34632
rect 16025 34623 16083 34629
rect 18414 34620 18420 34632
rect 18472 34620 18478 34672
rect 18782 34620 18788 34672
rect 18840 34660 18846 34672
rect 19978 34660 19984 34672
rect 18840 34632 19984 34660
rect 18840 34620 18846 34632
rect 19978 34620 19984 34632
rect 20036 34660 20042 34672
rect 20257 34663 20315 34669
rect 20257 34660 20269 34663
rect 20036 34632 20269 34660
rect 20036 34620 20042 34632
rect 20257 34629 20269 34632
rect 20303 34629 20315 34663
rect 25148 34660 25176 34691
rect 20257 34623 20315 34629
rect 20364 34632 25176 34660
rect 6086 34552 6092 34604
rect 6144 34592 6150 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 6144 34564 6561 34592
rect 6144 34552 6150 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 7926 34552 7932 34604
rect 7984 34552 7990 34604
rect 8846 34552 8852 34604
rect 8904 34552 8910 34604
rect 19610 34552 19616 34604
rect 19668 34592 19674 34604
rect 20364 34592 20392 34632
rect 19668 34564 20392 34592
rect 19668 34552 19674 34564
rect 22278 34552 22284 34604
rect 22336 34592 22342 34604
rect 22465 34595 22523 34601
rect 22465 34592 22477 34595
rect 22336 34564 22477 34592
rect 22336 34552 22342 34564
rect 22465 34561 22477 34564
rect 22511 34561 22523 34595
rect 22465 34555 22523 34561
rect 22646 34552 22652 34604
rect 22704 34592 22710 34604
rect 24581 34595 24639 34601
rect 24581 34592 24593 34595
rect 22704 34564 24593 34592
rect 22704 34552 22710 34564
rect 24581 34561 24593 34564
rect 24627 34561 24639 34595
rect 24581 34555 24639 34561
rect 25314 34552 25320 34604
rect 25372 34552 25378 34604
rect 7282 34484 7288 34536
rect 7340 34524 7346 34536
rect 8754 34524 8760 34536
rect 7340 34496 8760 34524
rect 7340 34484 7346 34496
rect 8754 34484 8760 34496
rect 8812 34484 8818 34536
rect 9582 34484 9588 34536
rect 9640 34524 9646 34536
rect 9858 34524 9864 34536
rect 9640 34496 9864 34524
rect 9640 34484 9646 34496
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 10410 34484 10416 34536
rect 10468 34524 10474 34536
rect 10962 34524 10968 34536
rect 10468 34496 10968 34524
rect 10468 34484 10474 34496
rect 10962 34484 10968 34496
rect 11020 34524 11026 34536
rect 11701 34527 11759 34533
rect 11701 34524 11713 34527
rect 11020 34496 11713 34524
rect 11020 34484 11026 34496
rect 11701 34493 11713 34496
rect 11747 34493 11759 34527
rect 11701 34487 11759 34493
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13814 34524 13820 34536
rect 13495 34496 13820 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13814 34484 13820 34496
rect 13872 34524 13878 34536
rect 14826 34524 14832 34536
rect 13872 34496 14832 34524
rect 13872 34484 13878 34496
rect 14826 34484 14832 34496
rect 14884 34484 14890 34536
rect 16117 34527 16175 34533
rect 16117 34493 16129 34527
rect 16163 34493 16175 34527
rect 16117 34487 16175 34493
rect 21269 34527 21327 34533
rect 21269 34493 21281 34527
rect 21315 34493 21327 34527
rect 21269 34487 21327 34493
rect 22557 34527 22615 34533
rect 22557 34493 22569 34527
rect 22603 34493 22615 34527
rect 23566 34524 23572 34536
rect 22557 34487 22615 34493
rect 23216 34496 23572 34524
rect 4798 34416 4804 34468
rect 4856 34456 4862 34468
rect 5626 34456 5632 34468
rect 4856 34428 5632 34456
rect 4856 34416 4862 34428
rect 5626 34416 5632 34428
rect 5684 34416 5690 34468
rect 11054 34456 11060 34468
rect 10704 34428 11060 34456
rect 9112 34391 9170 34397
rect 9112 34357 9124 34391
rect 9158 34388 9170 34391
rect 10134 34388 10140 34400
rect 9158 34360 10140 34388
rect 9158 34357 9170 34360
rect 9112 34351 9170 34357
rect 10134 34348 10140 34360
rect 10192 34388 10198 34400
rect 10704 34388 10732 34428
rect 11054 34416 11060 34428
rect 11112 34416 11118 34468
rect 15838 34416 15844 34468
rect 15896 34456 15902 34468
rect 16132 34456 16160 34487
rect 15896 34428 16160 34456
rect 15896 34416 15902 34428
rect 19886 34416 19892 34468
rect 19944 34456 19950 34468
rect 21284 34456 21312 34487
rect 19944 34428 21312 34456
rect 22572 34456 22600 34487
rect 22646 34456 22652 34468
rect 22572 34428 22652 34456
rect 19944 34416 19950 34428
rect 22646 34416 22652 34428
rect 22704 34416 22710 34468
rect 23216 34465 23244 34496
rect 23566 34484 23572 34496
rect 23624 34484 23630 34536
rect 23658 34484 23664 34536
rect 23716 34484 23722 34536
rect 23753 34527 23811 34533
rect 23753 34493 23765 34527
rect 23799 34493 23811 34527
rect 23753 34487 23811 34493
rect 23201 34459 23259 34465
rect 23201 34425 23213 34459
rect 23247 34425 23259 34459
rect 23768 34456 23796 34487
rect 23842 34456 23848 34468
rect 23768 34428 23848 34456
rect 23201 34419 23259 34425
rect 23842 34416 23848 34428
rect 23900 34416 23906 34468
rect 10192 34360 10732 34388
rect 10192 34348 10198 34360
rect 10962 34348 10968 34400
rect 11020 34388 11026 34400
rect 11790 34388 11796 34400
rect 11020 34360 11796 34388
rect 11020 34348 11026 34360
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 11964 34391 12022 34397
rect 11964 34357 11976 34391
rect 12010 34388 12022 34391
rect 12066 34388 12072 34400
rect 12010 34360 12072 34388
rect 12010 34357 12022 34360
rect 11964 34351 12022 34357
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 20714 34348 20720 34400
rect 20772 34348 20778 34400
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 5800 34187 5858 34193
rect 5800 34153 5812 34187
rect 5846 34184 5858 34187
rect 7374 34184 7380 34196
rect 5846 34156 7380 34184
rect 5846 34153 5858 34156
rect 5800 34147 5858 34153
rect 7374 34144 7380 34156
rect 7432 34144 7438 34196
rect 9122 34144 9128 34196
rect 9180 34144 9186 34196
rect 10686 34144 10692 34196
rect 10744 34184 10750 34196
rect 12161 34187 12219 34193
rect 12161 34184 12173 34187
rect 10744 34156 12173 34184
rect 10744 34144 10750 34156
rect 12161 34153 12173 34156
rect 12207 34184 12219 34187
rect 17681 34187 17739 34193
rect 12207 34156 12434 34184
rect 12207 34153 12219 34156
rect 12161 34147 12219 34153
rect 7190 34076 7196 34128
rect 7248 34116 7254 34128
rect 10226 34116 10232 34128
rect 7248 34088 10232 34116
rect 7248 34076 7254 34088
rect 10226 34076 10232 34088
rect 10284 34076 10290 34128
rect 12406 34116 12434 34156
rect 17681 34153 17693 34187
rect 17727 34184 17739 34187
rect 19702 34184 19708 34196
rect 17727 34156 19708 34184
rect 17727 34153 17739 34156
rect 17681 34147 17739 34153
rect 19702 34144 19708 34156
rect 19760 34144 19766 34196
rect 20162 34144 20168 34196
rect 20220 34184 20226 34196
rect 20533 34187 20591 34193
rect 20533 34184 20545 34187
rect 20220 34156 20545 34184
rect 20220 34144 20226 34156
rect 20533 34153 20545 34156
rect 20579 34184 20591 34187
rect 20898 34184 20904 34196
rect 20579 34156 20904 34184
rect 20579 34153 20591 34156
rect 20533 34147 20591 34153
rect 20898 34144 20904 34156
rect 20956 34144 20962 34196
rect 22278 34144 22284 34196
rect 22336 34184 22342 34196
rect 23293 34187 23351 34193
rect 23293 34184 23305 34187
rect 22336 34156 23305 34184
rect 22336 34144 22342 34156
rect 23293 34153 23305 34156
rect 23339 34153 23351 34187
rect 23293 34147 23351 34153
rect 25314 34144 25320 34196
rect 25372 34144 25378 34196
rect 12406 34088 13584 34116
rect 5534 34008 5540 34060
rect 5592 34008 5598 34060
rect 5810 34008 5816 34060
rect 5868 34048 5874 34060
rect 7285 34051 7343 34057
rect 7285 34048 7297 34051
rect 5868 34020 7297 34048
rect 5868 34008 5874 34020
rect 7285 34017 7297 34020
rect 7331 34048 7343 34051
rect 9214 34048 9220 34060
rect 7331 34020 9220 34048
rect 7331 34017 7343 34020
rect 7285 34011 7343 34017
rect 9214 34008 9220 34020
rect 9272 34048 9278 34060
rect 9677 34051 9735 34057
rect 9677 34048 9689 34051
rect 9272 34020 9689 34048
rect 9272 34008 9278 34020
rect 9677 34017 9689 34020
rect 9723 34017 9735 34051
rect 9677 34011 9735 34017
rect 10689 34051 10747 34057
rect 10689 34017 10701 34051
rect 10735 34048 10747 34051
rect 12526 34048 12532 34060
rect 10735 34020 12532 34048
rect 10735 34017 10747 34020
rect 10689 34011 10747 34017
rect 12526 34008 12532 34020
rect 12584 34008 12590 34060
rect 12618 34008 12624 34060
rect 12676 34048 12682 34060
rect 13556 34057 13584 34088
rect 13814 34076 13820 34128
rect 13872 34116 13878 34128
rect 13872 34088 16068 34116
rect 13872 34076 13878 34088
rect 13449 34051 13507 34057
rect 13449 34048 13461 34051
rect 12676 34020 13461 34048
rect 12676 34008 12682 34020
rect 13449 34017 13461 34020
rect 13495 34017 13507 34051
rect 13449 34011 13507 34017
rect 13541 34051 13599 34057
rect 13541 34017 13553 34051
rect 13587 34017 13599 34051
rect 13541 34011 13599 34017
rect 15930 34008 15936 34060
rect 15988 34008 15994 34060
rect 16040 34048 16068 34088
rect 19794 34076 19800 34128
rect 19852 34116 19858 34128
rect 21085 34119 21143 34125
rect 21085 34116 21097 34119
rect 19852 34088 21097 34116
rect 19852 34076 19858 34088
rect 21085 34085 21097 34088
rect 21131 34085 21143 34119
rect 21085 34079 21143 34085
rect 16040 34020 17448 34048
rect 7374 33940 7380 33992
rect 7432 33980 7438 33992
rect 7745 33983 7803 33989
rect 7745 33980 7757 33983
rect 7432 33952 7757 33980
rect 7432 33940 7438 33952
rect 7745 33949 7757 33952
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 8846 33940 8852 33992
rect 8904 33980 8910 33992
rect 9582 33980 9588 33992
rect 8904 33952 9588 33980
rect 8904 33940 8910 33952
rect 9582 33940 9588 33952
rect 9640 33980 9646 33992
rect 10410 33980 10416 33992
rect 9640 33952 10416 33980
rect 9640 33940 9646 33952
rect 10410 33940 10416 33952
rect 10468 33940 10474 33992
rect 11790 33940 11796 33992
rect 11848 33980 11854 33992
rect 12437 33983 12495 33989
rect 12437 33980 12449 33983
rect 11848 33952 12449 33980
rect 11848 33940 11854 33952
rect 12437 33949 12449 33952
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12802 33940 12808 33992
rect 12860 33980 12866 33992
rect 13722 33980 13728 33992
rect 12860 33952 13728 33980
rect 12860 33940 12866 33952
rect 13722 33940 13728 33952
rect 13780 33940 13786 33992
rect 17420 33980 17448 34020
rect 18414 34008 18420 34060
rect 18472 34048 18478 34060
rect 19061 34051 19119 34057
rect 19061 34048 19073 34051
rect 18472 34020 19073 34048
rect 18472 34008 18478 34020
rect 19061 34017 19073 34020
rect 19107 34048 19119 34051
rect 19981 34051 20039 34057
rect 19981 34048 19993 34051
rect 19107 34020 19993 34048
rect 19107 34017 19119 34020
rect 19061 34011 19119 34017
rect 19981 34017 19993 34020
rect 20027 34017 20039 34051
rect 19981 34011 20039 34017
rect 21634 34008 21640 34060
rect 21692 34008 21698 34060
rect 22738 34008 22744 34060
rect 22796 34008 22802 34060
rect 22925 34051 22983 34057
rect 22925 34017 22937 34051
rect 22971 34048 22983 34051
rect 23382 34048 23388 34060
rect 22971 34020 23388 34048
rect 22971 34017 22983 34020
rect 22925 34011 22983 34017
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 19610 33980 19616 33992
rect 17420 33952 19616 33980
rect 19610 33940 19616 33952
rect 19668 33940 19674 33992
rect 19797 33983 19855 33989
rect 19797 33949 19809 33983
rect 19843 33980 19855 33983
rect 20070 33980 20076 33992
rect 19843 33952 20076 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 20070 33940 20076 33952
rect 20128 33940 20134 33992
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 21545 33983 21603 33989
rect 21545 33980 21557 33983
rect 20680 33952 21557 33980
rect 20680 33940 20686 33952
rect 21545 33949 21557 33952
rect 21591 33980 21603 33983
rect 24210 33980 24216 33992
rect 21591 33952 24216 33980
rect 21591 33949 21603 33952
rect 21545 33943 21603 33949
rect 24210 33940 24216 33952
rect 24268 33940 24274 33992
rect 24302 33940 24308 33992
rect 24360 33980 24366 33992
rect 24765 33983 24823 33989
rect 24765 33980 24777 33983
rect 24360 33952 24777 33980
rect 24360 33940 24366 33952
rect 24765 33949 24777 33952
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 7038 33884 7236 33912
rect 7208 33856 7236 33884
rect 7650 33872 7656 33924
rect 7708 33912 7714 33924
rect 9493 33915 9551 33921
rect 9493 33912 9505 33915
rect 7708 33884 9505 33912
rect 7708 33872 7714 33884
rect 9493 33881 9505 33884
rect 9539 33881 9551 33915
rect 9493 33875 9551 33881
rect 9858 33872 9864 33924
rect 9916 33912 9922 33924
rect 10962 33912 10968 33924
rect 9916 33884 10968 33912
rect 9916 33872 9922 33884
rect 10962 33872 10968 33884
rect 11020 33912 11026 33924
rect 11020 33884 11178 33912
rect 11020 33872 11026 33884
rect 15562 33872 15568 33924
rect 15620 33912 15626 33924
rect 16209 33915 16267 33921
rect 16209 33912 16221 33915
rect 15620 33884 16221 33912
rect 15620 33872 15626 33884
rect 16209 33881 16221 33884
rect 16255 33881 16267 33915
rect 19889 33915 19947 33921
rect 16209 33875 16267 33881
rect 16316 33884 16698 33912
rect 17972 33884 19564 33912
rect 7190 33804 7196 33856
rect 7248 33844 7254 33856
rect 7561 33847 7619 33853
rect 7561 33844 7573 33847
rect 7248 33816 7573 33844
rect 7248 33804 7254 33816
rect 7561 33813 7573 33816
rect 7607 33844 7619 33847
rect 7926 33844 7932 33856
rect 7607 33816 7932 33844
rect 7607 33813 7619 33816
rect 7561 33807 7619 33813
rect 7926 33804 7932 33816
rect 7984 33844 7990 33856
rect 8481 33847 8539 33853
rect 8481 33844 8493 33847
rect 7984 33816 8493 33844
rect 7984 33804 7990 33816
rect 8481 33813 8493 33816
rect 8527 33813 8539 33847
rect 8481 33807 8539 33813
rect 9585 33847 9643 33853
rect 9585 33813 9597 33847
rect 9631 33844 9643 33847
rect 11974 33844 11980 33856
rect 9631 33816 11980 33844
rect 9631 33813 9643 33816
rect 9585 33807 9643 33813
rect 11974 33804 11980 33816
rect 12032 33804 12038 33856
rect 12802 33804 12808 33856
rect 12860 33844 12866 33856
rect 12989 33847 13047 33853
rect 12989 33844 13001 33847
rect 12860 33816 13001 33844
rect 12860 33804 12866 33816
rect 12989 33813 13001 33816
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 13357 33847 13415 33853
rect 13357 33813 13369 33847
rect 13403 33844 13415 33847
rect 13538 33844 13544 33856
rect 13403 33816 13544 33844
rect 13403 33813 13415 33816
rect 13357 33807 13415 33813
rect 13538 33804 13544 33816
rect 13596 33844 13602 33856
rect 14093 33847 14151 33853
rect 14093 33844 14105 33847
rect 13596 33816 14105 33844
rect 13596 33804 13602 33816
rect 14093 33813 14105 33816
rect 14139 33844 14151 33847
rect 15010 33844 15016 33856
rect 14139 33816 15016 33844
rect 14139 33813 14151 33816
rect 14093 33807 14151 33813
rect 15010 33804 15016 33816
rect 15068 33804 15074 33856
rect 16114 33804 16120 33856
rect 16172 33844 16178 33856
rect 16316 33844 16344 33884
rect 16172 33816 16344 33844
rect 16592 33844 16620 33884
rect 17972 33853 18000 33884
rect 17957 33847 18015 33853
rect 17957 33844 17969 33847
rect 16592 33816 17969 33844
rect 16172 33804 16178 33816
rect 17957 33813 17969 33816
rect 18003 33813 18015 33847
rect 17957 33807 18015 33813
rect 19058 33804 19064 33856
rect 19116 33844 19122 33856
rect 19429 33847 19487 33853
rect 19429 33844 19441 33847
rect 19116 33816 19441 33844
rect 19116 33804 19122 33816
rect 19429 33813 19441 33816
rect 19475 33813 19487 33847
rect 19536 33844 19564 33884
rect 19889 33881 19901 33915
rect 19935 33912 19947 33915
rect 19978 33912 19984 33924
rect 19935 33884 19984 33912
rect 19935 33881 19947 33884
rect 19889 33875 19947 33881
rect 19978 33872 19984 33884
rect 20036 33872 20042 33924
rect 24486 33912 24492 33924
rect 24320 33884 24492 33912
rect 24320 33856 24348 33884
rect 24486 33872 24492 33884
rect 24544 33912 24550 33924
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 24544 33884 25421 33912
rect 24544 33872 24550 33884
rect 25409 33881 25421 33884
rect 25455 33881 25467 33915
rect 25409 33875 25467 33881
rect 20162 33844 20168 33856
rect 19536 33816 20168 33844
rect 19429 33807 19487 33813
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 20622 33804 20628 33856
rect 20680 33804 20686 33856
rect 21450 33804 21456 33856
rect 21508 33804 21514 33856
rect 22278 33804 22284 33856
rect 22336 33804 22342 33856
rect 22462 33804 22468 33856
rect 22520 33844 22526 33856
rect 22649 33847 22707 33853
rect 22649 33844 22661 33847
rect 22520 33816 22661 33844
rect 22520 33804 22526 33816
rect 22649 33813 22661 33816
rect 22695 33813 22707 33847
rect 22649 33807 22707 33813
rect 24302 33804 24308 33856
rect 24360 33804 24366 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 10318 33600 10324 33652
rect 10376 33640 10382 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 10376 33612 10425 33640
rect 10376 33600 10382 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 10413 33603 10471 33609
rect 10778 33600 10784 33652
rect 10836 33640 10842 33652
rect 10873 33643 10931 33649
rect 10873 33640 10885 33643
rect 10836 33612 10885 33640
rect 10836 33600 10842 33612
rect 10873 33609 10885 33612
rect 10919 33609 10931 33643
rect 10873 33603 10931 33609
rect 11238 33600 11244 33652
rect 11296 33640 11302 33652
rect 12897 33643 12955 33649
rect 12897 33640 12909 33643
rect 11296 33612 12909 33640
rect 11296 33600 11302 33612
rect 12897 33609 12909 33612
rect 12943 33609 12955 33643
rect 12897 33603 12955 33609
rect 13357 33643 13415 33649
rect 13357 33609 13369 33643
rect 13403 33640 13415 33643
rect 13814 33640 13820 33652
rect 13403 33612 13820 33640
rect 13403 33609 13415 33612
rect 13357 33603 13415 33609
rect 1302 33464 1308 33516
rect 1360 33504 1366 33516
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 1360 33476 1777 33504
rect 1360 33464 1366 33476
rect 1765 33473 1777 33476
rect 1811 33504 1823 33507
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1811 33476 2053 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 10781 33507 10839 33513
rect 10781 33473 10793 33507
rect 10827 33504 10839 33507
rect 11606 33504 11612 33516
rect 10827 33476 11612 33504
rect 10827 33473 10839 33476
rect 10781 33467 10839 33473
rect 11606 33464 11612 33476
rect 11664 33464 11670 33516
rect 13262 33464 13268 33516
rect 13320 33464 13326 33516
rect 5350 33396 5356 33448
rect 5408 33396 5414 33448
rect 9766 33396 9772 33448
rect 9824 33396 9830 33448
rect 10965 33439 11023 33445
rect 10965 33405 10977 33439
rect 11011 33405 11023 33439
rect 10965 33399 11023 33405
rect 12805 33439 12863 33445
rect 12805 33405 12817 33439
rect 12851 33436 12863 33439
rect 13372 33436 13400 33603
rect 13814 33600 13820 33612
rect 13872 33600 13878 33652
rect 14550 33640 14556 33652
rect 14108 33612 14556 33640
rect 14108 33513 14136 33612
rect 14550 33600 14556 33612
rect 14608 33640 14614 33652
rect 15930 33640 15936 33652
rect 14608 33612 15936 33640
rect 14608 33600 14614 33612
rect 15930 33600 15936 33612
rect 15988 33600 15994 33652
rect 19150 33600 19156 33652
rect 19208 33640 19214 33652
rect 19797 33643 19855 33649
rect 19797 33640 19809 33643
rect 19208 33612 19809 33640
rect 19208 33600 19214 33612
rect 19797 33609 19809 33612
rect 19843 33640 19855 33643
rect 19978 33640 19984 33652
rect 19843 33612 19984 33640
rect 19843 33609 19855 33612
rect 19797 33603 19855 33609
rect 19978 33600 19984 33612
rect 20036 33600 20042 33652
rect 20257 33643 20315 33649
rect 20257 33609 20269 33643
rect 20303 33609 20315 33643
rect 20257 33603 20315 33609
rect 20717 33643 20775 33649
rect 20717 33609 20729 33643
rect 20763 33640 20775 33643
rect 21174 33640 21180 33652
rect 20763 33612 21180 33640
rect 20763 33609 20775 33612
rect 20717 33603 20775 33609
rect 14366 33532 14372 33584
rect 14424 33572 14430 33584
rect 14642 33572 14648 33584
rect 14424 33544 14648 33572
rect 14424 33532 14430 33544
rect 14642 33532 14648 33544
rect 14700 33572 14706 33584
rect 18322 33572 18328 33584
rect 14700 33544 14858 33572
rect 18064 33544 18328 33572
rect 14700 33532 14706 33544
rect 18064 33513 18092 33544
rect 18322 33532 18328 33544
rect 18380 33532 18386 33584
rect 20162 33572 20168 33584
rect 19550 33544 20168 33572
rect 20162 33532 20168 33544
rect 20220 33532 20226 33584
rect 20272 33572 20300 33603
rect 21174 33600 21180 33612
rect 21232 33640 21238 33652
rect 21269 33643 21327 33649
rect 21269 33640 21281 33643
rect 21232 33612 21281 33640
rect 21232 33600 21238 33612
rect 21269 33609 21281 33612
rect 21315 33609 21327 33643
rect 21269 33603 21327 33609
rect 21450 33600 21456 33652
rect 21508 33640 21514 33652
rect 22649 33643 22707 33649
rect 22649 33640 22661 33643
rect 21508 33612 22661 33640
rect 21508 33600 21514 33612
rect 22649 33609 22661 33612
rect 22695 33609 22707 33643
rect 22649 33603 22707 33609
rect 25222 33600 25228 33652
rect 25280 33600 25286 33652
rect 23658 33572 23664 33584
rect 20272 33544 23664 33572
rect 23658 33532 23664 33544
rect 23716 33532 23722 33584
rect 24302 33532 24308 33584
rect 24360 33532 24366 33584
rect 14093 33507 14151 33513
rect 14093 33473 14105 33507
rect 14139 33473 14151 33507
rect 14093 33467 14151 33473
rect 18049 33507 18107 33513
rect 18049 33473 18061 33507
rect 18095 33473 18107 33507
rect 18049 33467 18107 33473
rect 20622 33464 20628 33516
rect 20680 33464 20686 33516
rect 20916 33476 22140 33504
rect 12851 33408 13400 33436
rect 12851 33405 12863 33408
rect 12805 33399 12863 33405
rect 8294 33328 8300 33380
rect 8352 33368 8358 33380
rect 10980 33368 11008 33399
rect 13446 33396 13452 33448
rect 13504 33396 13510 33448
rect 14369 33439 14427 33445
rect 14369 33405 14381 33439
rect 14415 33436 14427 33439
rect 16666 33436 16672 33448
rect 14415 33408 16672 33436
rect 14415 33405 14427 33408
rect 14369 33399 14427 33405
rect 16666 33396 16672 33408
rect 16724 33396 16730 33448
rect 20916 33445 20944 33476
rect 18325 33439 18383 33445
rect 18325 33405 18337 33439
rect 18371 33436 18383 33439
rect 20901 33439 20959 33445
rect 18371 33408 20852 33436
rect 18371 33405 18383 33408
rect 18325 33399 18383 33405
rect 8352 33340 11008 33368
rect 20824 33368 20852 33408
rect 20901 33405 20913 33439
rect 20947 33405 20959 33439
rect 20901 33399 20959 33405
rect 20990 33396 20996 33448
rect 21048 33436 21054 33448
rect 22005 33439 22063 33445
rect 22005 33436 22017 33439
rect 21048 33408 22017 33436
rect 21048 33396 21054 33408
rect 22005 33405 22017 33408
rect 22051 33405 22063 33439
rect 22112 33436 22140 33476
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 23477 33507 23535 33513
rect 23477 33504 23489 33507
rect 22244 33476 23489 33504
rect 22244 33464 22250 33476
rect 23477 33473 23489 33476
rect 23523 33473 23535 33507
rect 23477 33467 23535 33473
rect 23290 33436 23296 33448
rect 22112 33408 23296 33436
rect 22005 33399 22063 33405
rect 23290 33396 23296 33408
rect 23348 33396 23354 33448
rect 23750 33396 23756 33448
rect 23808 33396 23814 33448
rect 21634 33368 21640 33380
rect 20824 33340 21640 33368
rect 8352 33328 8358 33340
rect 21634 33328 21640 33340
rect 21692 33328 21698 33380
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 3510 33300 3516 33312
rect 1627 33272 3516 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 3510 33260 3516 33272
rect 3568 33260 3574 33312
rect 7190 33260 7196 33312
rect 7248 33260 7254 33312
rect 12434 33260 12440 33312
rect 12492 33300 12498 33312
rect 12529 33303 12587 33309
rect 12529 33300 12541 33303
rect 12492 33272 12541 33300
rect 12492 33260 12498 33272
rect 12529 33269 12541 33272
rect 12575 33300 12587 33303
rect 13262 33300 13268 33312
rect 12575 33272 13268 33300
rect 12575 33269 12587 33272
rect 12529 33263 12587 33269
rect 13262 33260 13268 33272
rect 13320 33260 13326 33312
rect 13446 33260 13452 33312
rect 13504 33300 13510 33312
rect 15838 33300 15844 33312
rect 13504 33272 15844 33300
rect 13504 33260 13510 33272
rect 15838 33260 15844 33272
rect 15896 33260 15902 33312
rect 16114 33260 16120 33312
rect 16172 33260 16178 33312
rect 16390 33260 16396 33312
rect 16448 33300 16454 33312
rect 16850 33300 16856 33312
rect 16448 33272 16856 33300
rect 16448 33260 16454 33272
rect 16850 33260 16856 33272
rect 16908 33260 16914 33312
rect 20346 33260 20352 33312
rect 20404 33300 20410 33312
rect 22738 33300 22744 33312
rect 20404 33272 22744 33300
rect 20404 33260 20410 33272
rect 22738 33260 22744 33272
rect 22796 33260 22802 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 7466 33056 7472 33108
rect 7524 33056 7530 33108
rect 9306 33056 9312 33108
rect 9364 33096 9370 33108
rect 9401 33099 9459 33105
rect 9401 33096 9413 33099
rect 9364 33068 9413 33096
rect 9364 33056 9370 33068
rect 9401 33065 9413 33068
rect 9447 33065 9459 33099
rect 9401 33059 9459 33065
rect 10226 33056 10232 33108
rect 10284 33096 10290 33108
rect 10597 33099 10655 33105
rect 10597 33096 10609 33099
rect 10284 33068 10609 33096
rect 10284 33056 10290 33068
rect 10597 33065 10609 33068
rect 10643 33065 10655 33099
rect 10597 33059 10655 33065
rect 7009 33031 7067 33037
rect 7009 32997 7021 33031
rect 7055 33028 7067 33031
rect 7558 33028 7564 33040
rect 7055 33000 7564 33028
rect 7055 32997 7067 33000
rect 7009 32991 7067 32997
rect 7558 32988 7564 33000
rect 7616 32988 7622 33040
rect 9122 33028 9128 33040
rect 7668 33000 9128 33028
rect 5261 32963 5319 32969
rect 5261 32929 5273 32963
rect 5307 32960 5319 32963
rect 5534 32960 5540 32972
rect 5307 32932 5540 32960
rect 5307 32929 5319 32932
rect 5261 32923 5319 32929
rect 5534 32920 5540 32932
rect 5592 32920 5598 32972
rect 7190 32960 7196 32972
rect 6656 32932 7196 32960
rect 6656 32878 6684 32932
rect 7190 32920 7196 32932
rect 7248 32960 7254 32972
rect 7668 32960 7696 33000
rect 9122 32988 9128 33000
rect 9180 32988 9186 33040
rect 7248 32932 7696 32960
rect 8113 32963 8171 32969
rect 7248 32920 7254 32932
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8294 32960 8300 32972
rect 8159 32932 8300 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 8128 32892 8156 32923
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 10045 32963 10103 32969
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10134 32960 10140 32972
rect 10091 32932 10140 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 10134 32920 10140 32932
rect 10192 32920 10198 32972
rect 7668 32864 8156 32892
rect 5537 32827 5595 32833
rect 5537 32793 5549 32827
rect 5583 32793 5595 32827
rect 5537 32787 5595 32793
rect 5552 32756 5580 32787
rect 7668 32756 7696 32864
rect 9766 32852 9772 32904
rect 9824 32852 9830 32904
rect 7742 32784 7748 32836
rect 7800 32824 7806 32836
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7800 32796 7941 32824
rect 7800 32784 7806 32796
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 10612 32824 10640 33059
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 11149 33099 11207 33105
rect 11149 33096 11161 33099
rect 10928 33068 11161 33096
rect 10928 33056 10934 33068
rect 11149 33065 11161 33068
rect 11195 33065 11207 33099
rect 11149 33059 11207 33065
rect 12158 33056 12164 33108
rect 12216 33056 12222 33108
rect 14366 33096 14372 33108
rect 12406 33068 14372 33096
rect 10873 32963 10931 32969
rect 10873 32929 10885 32963
rect 10919 32960 10931 32963
rect 11514 32960 11520 32972
rect 10919 32932 11520 32960
rect 10919 32929 10931 32932
rect 10873 32923 10931 32929
rect 11514 32920 11520 32932
rect 11572 32960 11578 32972
rect 11609 32963 11667 32969
rect 11609 32960 11621 32963
rect 11572 32932 11621 32960
rect 11572 32920 11578 32932
rect 11609 32929 11621 32932
rect 11655 32929 11667 32963
rect 11609 32923 11667 32929
rect 11793 32963 11851 32969
rect 11793 32929 11805 32963
rect 11839 32960 11851 32963
rect 12176 32960 12204 33056
rect 11839 32932 12204 32960
rect 11839 32929 11851 32932
rect 11793 32923 11851 32929
rect 11624 32892 11652 32923
rect 12406 32892 12434 33068
rect 14366 33056 14372 33068
rect 14424 33056 14430 33108
rect 15010 33056 15016 33108
rect 15068 33096 15074 33108
rect 20622 33096 20628 33108
rect 15068 33068 20628 33096
rect 15068 33056 15074 33068
rect 20622 33056 20628 33068
rect 20680 33056 20686 33108
rect 20898 33056 20904 33108
rect 20956 33096 20962 33108
rect 25133 33099 25191 33105
rect 25133 33096 25145 33099
rect 20956 33068 25145 33096
rect 20956 33056 20962 33068
rect 25133 33065 25145 33068
rect 25179 33065 25191 33099
rect 25133 33059 25191 33065
rect 12618 32988 12624 33040
rect 12676 33028 12682 33040
rect 13906 33028 13912 33040
rect 12676 33000 13912 33028
rect 12676 32988 12682 33000
rect 13906 32988 13912 33000
rect 13964 32988 13970 33040
rect 14277 33031 14335 33037
rect 14277 32997 14289 33031
rect 14323 33028 14335 33031
rect 17034 33028 17040 33040
rect 14323 33000 17040 33028
rect 14323 32997 14335 33000
rect 14277 32991 14335 32997
rect 17034 32988 17040 33000
rect 17092 32988 17098 33040
rect 17126 32988 17132 33040
rect 17184 32988 17190 33040
rect 20070 33028 20076 33040
rect 17788 33000 20076 33028
rect 11624 32864 12434 32892
rect 13924 32892 13952 32988
rect 14458 32920 14464 32972
rect 14516 32960 14522 32972
rect 14737 32963 14795 32969
rect 14737 32960 14749 32963
rect 14516 32932 14749 32960
rect 14516 32920 14522 32932
rect 14737 32929 14749 32932
rect 14783 32929 14795 32963
rect 14737 32923 14795 32929
rect 14826 32920 14832 32972
rect 14884 32920 14890 32972
rect 16390 32960 16396 32972
rect 15764 32932 16396 32960
rect 15764 32901 15792 32932
rect 16390 32920 16396 32932
rect 16448 32920 16454 32972
rect 16482 32920 16488 32972
rect 16540 32960 16546 32972
rect 16669 32963 16727 32969
rect 16669 32960 16681 32963
rect 16540 32932 16681 32960
rect 16540 32920 16546 32932
rect 16669 32929 16681 32932
rect 16715 32929 16727 32963
rect 16669 32923 16727 32929
rect 16850 32920 16856 32972
rect 16908 32960 16914 32972
rect 17788 32960 17816 33000
rect 20070 32988 20076 33000
rect 20128 32988 20134 33040
rect 22554 33028 22560 33040
rect 20364 33000 20668 33028
rect 20364 32969 20392 33000
rect 20257 32963 20315 32969
rect 20257 32960 20269 32963
rect 16908 32932 17816 32960
rect 19444 32932 20269 32960
rect 16908 32920 16914 32932
rect 15749 32895 15807 32901
rect 15749 32892 15761 32895
rect 13924 32864 15761 32892
rect 15749 32861 15761 32864
rect 15795 32861 15807 32895
rect 15749 32855 15807 32861
rect 15838 32852 15844 32904
rect 15896 32892 15902 32904
rect 16577 32895 16635 32901
rect 16577 32892 16589 32895
rect 15896 32864 16589 32892
rect 15896 32852 15902 32864
rect 16577 32861 16589 32864
rect 16623 32892 16635 32895
rect 16758 32892 16764 32904
rect 16623 32864 16764 32892
rect 16623 32861 16635 32864
rect 16577 32855 16635 32861
rect 16758 32852 16764 32864
rect 16816 32892 16822 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 16816 32864 17325 32892
rect 16816 32852 16822 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17313 32855 17371 32861
rect 17494 32852 17500 32904
rect 17552 32892 17558 32904
rect 19242 32892 19248 32904
rect 17552 32864 19248 32892
rect 17552 32852 17558 32864
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 11517 32827 11575 32833
rect 11517 32824 11529 32827
rect 10612 32796 11529 32824
rect 7929 32787 7987 32793
rect 11517 32793 11529 32796
rect 11563 32824 11575 32827
rect 11882 32824 11888 32836
rect 11563 32796 11888 32824
rect 11563 32793 11575 32796
rect 11517 32787 11575 32793
rect 11882 32784 11888 32796
rect 11940 32784 11946 32836
rect 14366 32784 14372 32836
rect 14424 32824 14430 32836
rect 19444 32833 19472 32932
rect 20257 32929 20269 32932
rect 20303 32929 20315 32963
rect 20257 32923 20315 32929
rect 20349 32963 20407 32969
rect 20349 32929 20361 32963
rect 20395 32929 20407 32963
rect 20640 32960 20668 33000
rect 20824 33000 22560 33028
rect 20824 32960 20852 33000
rect 22554 32988 22560 33000
rect 22612 32988 22618 33040
rect 22925 33031 22983 33037
rect 22925 32997 22937 33031
rect 22971 33028 22983 33031
rect 24026 33028 24032 33040
rect 22971 33000 24032 33028
rect 22971 32997 22983 33000
rect 22925 32991 22983 32997
rect 20640 32932 20852 32960
rect 20349 32923 20407 32929
rect 21634 32920 21640 32972
rect 21692 32920 21698 32972
rect 22940 32960 22968 32991
rect 24026 32988 24032 33000
rect 24084 32988 24090 33040
rect 21744 32932 22968 32960
rect 20165 32895 20223 32901
rect 20165 32861 20177 32895
rect 20211 32892 20223 32895
rect 20990 32892 20996 32904
rect 20211 32864 20996 32892
rect 20211 32861 20223 32864
rect 20165 32855 20223 32861
rect 20990 32852 20996 32864
rect 21048 32852 21054 32904
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 21361 32895 21419 32901
rect 21361 32892 21373 32895
rect 21232 32864 21373 32892
rect 21232 32852 21238 32864
rect 21361 32861 21373 32864
rect 21407 32892 21419 32895
rect 21450 32892 21456 32904
rect 21407 32864 21456 32892
rect 21407 32861 21419 32864
rect 21361 32855 21419 32861
rect 21450 32852 21456 32864
rect 21508 32892 21514 32904
rect 21744 32892 21772 32932
rect 21508 32864 21772 32892
rect 21508 32852 21514 32864
rect 22370 32852 22376 32904
rect 22428 32852 22434 32904
rect 24857 32895 24915 32901
rect 24857 32861 24869 32895
rect 24903 32892 24915 32895
rect 25314 32892 25320 32904
rect 24903 32864 25320 32892
rect 24903 32861 24915 32864
rect 24857 32855 24915 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 19429 32827 19487 32833
rect 19429 32824 19441 32827
rect 14424 32796 19441 32824
rect 14424 32784 14430 32796
rect 19429 32793 19441 32796
rect 19475 32793 19487 32827
rect 22462 32824 22468 32836
rect 19429 32787 19487 32793
rect 19812 32796 22468 32824
rect 5552 32728 7696 32756
rect 7834 32716 7840 32768
rect 7892 32716 7898 32768
rect 9490 32716 9496 32768
rect 9548 32756 9554 32768
rect 9861 32759 9919 32765
rect 9861 32756 9873 32759
rect 9548 32728 9873 32756
rect 9548 32716 9554 32728
rect 9861 32725 9873 32728
rect 9907 32725 9919 32759
rect 9861 32719 9919 32725
rect 14642 32716 14648 32768
rect 14700 32716 14706 32768
rect 16114 32716 16120 32768
rect 16172 32716 16178 32768
rect 16390 32716 16396 32768
rect 16448 32756 16454 32768
rect 16485 32759 16543 32765
rect 16485 32756 16497 32759
rect 16448 32728 16497 32756
rect 16448 32716 16454 32728
rect 16485 32725 16497 32728
rect 16531 32725 16543 32759
rect 16485 32719 16543 32725
rect 17957 32759 18015 32765
rect 17957 32725 17969 32759
rect 18003 32756 18015 32759
rect 18598 32756 18604 32768
rect 18003 32728 18604 32756
rect 18003 32725 18015 32728
rect 17957 32719 18015 32725
rect 18598 32716 18604 32728
rect 18656 32716 18662 32768
rect 19812 32765 19840 32796
rect 22462 32784 22468 32796
rect 22520 32784 22526 32836
rect 19797 32759 19855 32765
rect 19797 32725 19809 32759
rect 19843 32725 19855 32759
rect 19797 32719 19855 32725
rect 20070 32716 20076 32768
rect 20128 32756 20134 32768
rect 20898 32756 20904 32768
rect 20128 32728 20904 32756
rect 20128 32716 20134 32728
rect 20898 32716 20904 32728
rect 20956 32716 20962 32768
rect 20993 32759 21051 32765
rect 20993 32725 21005 32759
rect 21039 32756 21051 32759
rect 21266 32756 21272 32768
rect 21039 32728 21272 32756
rect 21039 32725 21051 32728
rect 20993 32719 21051 32725
rect 21266 32716 21272 32728
rect 21324 32716 21330 32768
rect 21453 32759 21511 32765
rect 21453 32725 21465 32759
rect 21499 32756 21511 32759
rect 21634 32756 21640 32768
rect 21499 32728 21640 32756
rect 21499 32725 21511 32728
rect 21453 32719 21511 32725
rect 21634 32716 21640 32728
rect 21692 32716 21698 32768
rect 22189 32759 22247 32765
rect 22189 32725 22201 32759
rect 22235 32756 22247 32759
rect 22370 32756 22376 32768
rect 22235 32728 22376 32756
rect 22235 32725 22247 32728
rect 22189 32719 22247 32725
rect 22370 32716 22376 32728
rect 22428 32716 22434 32768
rect 22554 32716 22560 32768
rect 22612 32756 22618 32768
rect 22649 32759 22707 32765
rect 22649 32756 22661 32759
rect 22612 32728 22661 32756
rect 22612 32716 22618 32728
rect 22649 32725 22661 32728
rect 22695 32725 22707 32759
rect 22649 32719 22707 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 4614 32512 4620 32564
rect 4672 32512 4678 32564
rect 4982 32512 4988 32564
rect 5040 32512 5046 32564
rect 5350 32512 5356 32564
rect 5408 32512 5414 32564
rect 6917 32555 6975 32561
rect 6917 32521 6929 32555
rect 6963 32552 6975 32555
rect 7834 32552 7840 32564
rect 6963 32524 7840 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 11977 32555 12035 32561
rect 11977 32521 11989 32555
rect 12023 32552 12035 32555
rect 14642 32552 14648 32564
rect 12023 32524 14648 32552
rect 12023 32521 12035 32524
rect 11977 32515 12035 32521
rect 14642 32512 14648 32524
rect 14700 32512 14706 32564
rect 14734 32512 14740 32564
rect 14792 32552 14798 32564
rect 14792 32524 14964 32552
rect 14792 32512 14798 32524
rect 4632 32484 4660 32512
rect 4890 32484 4896 32496
rect 4632 32456 4896 32484
rect 4890 32444 4896 32456
rect 4948 32484 4954 32496
rect 5445 32487 5503 32493
rect 5445 32484 5457 32487
rect 4948 32456 5457 32484
rect 4948 32444 4954 32456
rect 5445 32453 5457 32456
rect 5491 32453 5503 32487
rect 5445 32447 5503 32453
rect 5534 32444 5540 32496
rect 5592 32484 5598 32496
rect 6178 32484 6184 32496
rect 5592 32456 6184 32484
rect 5592 32444 5598 32456
rect 6178 32444 6184 32456
rect 6236 32484 6242 32496
rect 9122 32484 9128 32496
rect 6236 32456 7604 32484
rect 9062 32456 9128 32484
rect 6236 32444 6242 32456
rect 7576 32425 7604 32456
rect 9122 32444 9128 32456
rect 9180 32484 9186 32496
rect 10226 32484 10232 32496
rect 9180 32456 10232 32484
rect 9180 32444 9186 32456
rect 10226 32444 10232 32456
rect 10284 32484 10290 32496
rect 10962 32484 10968 32496
rect 10284 32456 10968 32484
rect 10284 32444 10290 32456
rect 10962 32444 10968 32456
rect 11020 32444 11026 32496
rect 12526 32444 12532 32496
rect 12584 32484 12590 32496
rect 12584 32456 14504 32484
rect 12584 32444 12590 32456
rect 7561 32419 7619 32425
rect 7561 32385 7573 32419
rect 7607 32385 7619 32419
rect 7561 32379 7619 32385
rect 12345 32419 12403 32425
rect 12345 32385 12357 32419
rect 12391 32416 12403 32419
rect 13173 32419 13231 32425
rect 13173 32416 13185 32419
rect 12391 32388 13185 32416
rect 12391 32385 12403 32388
rect 12345 32379 12403 32385
rect 13173 32385 13185 32388
rect 13219 32385 13231 32419
rect 13173 32379 13231 32385
rect 5442 32308 5448 32360
rect 5500 32348 5506 32360
rect 5537 32351 5595 32357
rect 5537 32348 5549 32351
rect 5500 32320 5549 32348
rect 5500 32308 5506 32320
rect 5537 32317 5549 32320
rect 5583 32317 5595 32351
rect 7837 32351 7895 32357
rect 7837 32348 7849 32351
rect 5537 32311 5595 32317
rect 7576 32320 7849 32348
rect 7576 32292 7604 32320
rect 7837 32317 7849 32320
rect 7883 32317 7895 32351
rect 7837 32311 7895 32317
rect 9858 32308 9864 32360
rect 9916 32308 9922 32360
rect 11701 32351 11759 32357
rect 11701 32317 11713 32351
rect 11747 32348 11759 32351
rect 12250 32348 12256 32360
rect 11747 32320 12256 32348
rect 11747 32317 11759 32320
rect 11701 32311 11759 32317
rect 12250 32308 12256 32320
rect 12308 32348 12314 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12308 32320 12449 32348
rect 12308 32308 12314 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12437 32311 12495 32317
rect 12529 32351 12587 32357
rect 12529 32317 12541 32351
rect 12575 32317 12587 32351
rect 14476 32348 14504 32456
rect 14826 32444 14832 32496
rect 14884 32444 14890 32496
rect 14936 32484 14964 32524
rect 16114 32512 16120 32564
rect 16172 32552 16178 32564
rect 17313 32555 17371 32561
rect 17313 32552 17325 32555
rect 16172 32524 17325 32552
rect 16172 32512 16178 32524
rect 17313 32521 17325 32524
rect 17359 32521 17371 32555
rect 19245 32555 19303 32561
rect 19245 32552 19257 32555
rect 17313 32515 17371 32521
rect 18340 32524 19257 32552
rect 14936 32456 15318 32484
rect 17218 32444 17224 32496
rect 17276 32444 17282 32496
rect 14550 32376 14556 32428
rect 14608 32376 14614 32428
rect 18340 32416 18368 32524
rect 19245 32521 19257 32524
rect 19291 32552 19303 32555
rect 19291 32524 20576 32552
rect 19291 32521 19303 32524
rect 19245 32515 19303 32521
rect 18417 32419 18475 32425
rect 18417 32416 18429 32419
rect 16224 32388 18429 32416
rect 16224 32348 16252 32388
rect 18417 32385 18429 32388
rect 18463 32385 18475 32419
rect 18417 32379 18475 32385
rect 18509 32419 18567 32425
rect 18509 32385 18521 32419
rect 18555 32416 18567 32419
rect 18874 32416 18880 32428
rect 18555 32388 18880 32416
rect 18555 32385 18567 32388
rect 18509 32379 18567 32385
rect 18874 32376 18880 32388
rect 18932 32416 18938 32428
rect 19061 32419 19119 32425
rect 19061 32416 19073 32419
rect 18932 32388 19073 32416
rect 18932 32376 18938 32388
rect 19061 32385 19073 32388
rect 19107 32385 19119 32419
rect 19061 32379 19119 32385
rect 19242 32376 19248 32428
rect 19300 32416 19306 32428
rect 20257 32419 20315 32425
rect 20257 32416 20269 32419
rect 19300 32388 20269 32416
rect 19300 32376 19306 32388
rect 20257 32385 20269 32388
rect 20303 32385 20315 32419
rect 20548 32416 20576 32524
rect 20990 32512 20996 32564
rect 21048 32552 21054 32564
rect 21177 32555 21235 32561
rect 21177 32552 21189 32555
rect 21048 32524 21189 32552
rect 21048 32512 21054 32524
rect 21177 32521 21189 32524
rect 21223 32552 21235 32555
rect 21818 32552 21824 32564
rect 21223 32524 21824 32552
rect 21223 32521 21235 32524
rect 21177 32515 21235 32521
rect 21818 32512 21824 32524
rect 21876 32512 21882 32564
rect 25133 32555 25191 32561
rect 25133 32521 25145 32555
rect 25179 32521 25191 32555
rect 25133 32515 25191 32521
rect 25148 32484 25176 32515
rect 20824 32456 25176 32484
rect 20824 32416 20852 32456
rect 20548 32388 20852 32416
rect 20257 32379 20315 32385
rect 20898 32376 20904 32428
rect 20956 32416 20962 32428
rect 21085 32419 21143 32425
rect 21085 32416 21097 32419
rect 20956 32388 21097 32416
rect 20956 32376 20962 32388
rect 21085 32385 21097 32388
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22373 32419 22431 32425
rect 22373 32416 22385 32419
rect 22152 32388 22385 32416
rect 22152 32376 22158 32388
rect 22373 32385 22385 32388
rect 22419 32385 22431 32419
rect 22373 32379 22431 32385
rect 22738 32376 22744 32428
rect 22796 32416 22802 32428
rect 23017 32419 23075 32425
rect 23017 32416 23029 32419
rect 22796 32388 23029 32416
rect 22796 32376 22802 32388
rect 23017 32385 23029 32388
rect 23063 32385 23075 32419
rect 23017 32379 23075 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25317 32419 25375 32425
rect 25317 32416 25329 32419
rect 24903 32388 25329 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25317 32385 25329 32388
rect 25363 32416 25375 32419
rect 25406 32416 25412 32428
rect 25363 32388 25412 32416
rect 25363 32385 25375 32388
rect 25317 32379 25375 32385
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 14476 32320 16252 32348
rect 16301 32351 16359 32357
rect 12529 32311 12587 32317
rect 16301 32317 16313 32351
rect 16347 32348 16359 32351
rect 16666 32348 16672 32360
rect 16347 32320 16672 32348
rect 16347 32317 16359 32320
rect 16301 32311 16359 32317
rect 7558 32240 7564 32292
rect 7616 32240 7622 32292
rect 12066 32240 12072 32292
rect 12124 32280 12130 32292
rect 12544 32280 12572 32311
rect 16666 32308 16672 32320
rect 16724 32308 16730 32360
rect 17497 32351 17555 32357
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 17770 32348 17776 32360
rect 17543 32320 17776 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 17770 32308 17776 32320
rect 17828 32308 17834 32360
rect 18598 32308 18604 32360
rect 18656 32308 18662 32360
rect 20622 32348 20628 32360
rect 18708 32320 20628 32348
rect 13538 32280 13544 32292
rect 12124 32252 12572 32280
rect 12636 32252 13544 32280
rect 12124 32240 12130 32252
rect 9214 32172 9220 32224
rect 9272 32212 9278 32224
rect 9309 32215 9367 32221
rect 9309 32212 9321 32215
rect 9272 32184 9321 32212
rect 9272 32172 9278 32184
rect 9309 32181 9321 32184
rect 9355 32181 9367 32215
rect 9309 32175 9367 32181
rect 10226 32172 10232 32224
rect 10284 32212 10290 32224
rect 10321 32215 10379 32221
rect 10321 32212 10333 32215
rect 10284 32184 10333 32212
rect 10284 32172 10290 32184
rect 10321 32181 10333 32184
rect 10367 32181 10379 32215
rect 10321 32175 10379 32181
rect 12526 32172 12532 32224
rect 12584 32212 12590 32224
rect 12636 32212 12664 32252
rect 13538 32240 13544 32252
rect 13596 32240 13602 32292
rect 15930 32240 15936 32292
rect 15988 32280 15994 32292
rect 15988 32252 17080 32280
rect 15988 32240 15994 32252
rect 12584 32184 12664 32212
rect 12584 32172 12590 32184
rect 12710 32172 12716 32224
rect 12768 32212 12774 32224
rect 14458 32212 14464 32224
rect 12768 32184 14464 32212
rect 12768 32172 12774 32184
rect 14458 32172 14464 32184
rect 14516 32172 14522 32224
rect 14550 32172 14556 32224
rect 14608 32212 14614 32224
rect 15194 32212 15200 32224
rect 14608 32184 15200 32212
rect 14608 32172 14614 32184
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 16853 32215 16911 32221
rect 16853 32181 16865 32215
rect 16899 32212 16911 32215
rect 16942 32212 16948 32224
rect 16899 32184 16948 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 17052 32212 17080 32252
rect 17126 32240 17132 32292
rect 17184 32280 17190 32292
rect 18708 32280 18736 32320
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 21358 32308 21364 32360
rect 21416 32348 21422 32360
rect 21416 32320 21588 32348
rect 21416 32308 21422 32320
rect 17184 32252 18736 32280
rect 17184 32240 17190 32252
rect 17954 32212 17960 32224
rect 17052 32184 17960 32212
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 18049 32215 18107 32221
rect 18049 32181 18061 32215
rect 18095 32212 18107 32215
rect 18690 32212 18696 32224
rect 18095 32184 18696 32212
rect 18095 32181 18107 32184
rect 18049 32175 18107 32181
rect 18690 32172 18696 32184
rect 18748 32172 18754 32224
rect 20070 32172 20076 32224
rect 20128 32172 20134 32224
rect 20717 32215 20775 32221
rect 20717 32181 20729 32215
rect 20763 32212 20775 32215
rect 21358 32212 21364 32224
rect 20763 32184 21364 32212
rect 20763 32181 20775 32184
rect 20717 32175 20775 32181
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 21560 32212 21588 32320
rect 21818 32212 21824 32224
rect 21560 32184 21824 32212
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 22094 32172 22100 32224
rect 22152 32212 22158 32224
rect 22189 32215 22247 32221
rect 22189 32212 22201 32215
rect 22152 32184 22201 32212
rect 22152 32172 22158 32184
rect 22189 32181 22201 32184
rect 22235 32181 22247 32215
rect 22189 32175 22247 32181
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 22833 32215 22891 32221
rect 22833 32212 22845 32215
rect 22796 32184 22845 32212
rect 22796 32172 22802 32184
rect 22833 32181 22845 32184
rect 22879 32181 22891 32215
rect 22833 32175 22891 32181
rect 23290 32172 23296 32224
rect 23348 32172 23354 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 7929 32011 7987 32017
rect 7929 31977 7941 32011
rect 7975 32008 7987 32011
rect 8294 32008 8300 32020
rect 7975 31980 8300 32008
rect 7975 31977 7987 31980
rect 7929 31971 7987 31977
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 8573 32011 8631 32017
rect 8573 31977 8585 32011
rect 8619 32008 8631 32011
rect 9122 32008 9128 32020
rect 8619 31980 9128 32008
rect 8619 31977 8631 31980
rect 8573 31971 8631 31977
rect 6178 31832 6184 31884
rect 6236 31832 6242 31884
rect 6457 31875 6515 31881
rect 6457 31841 6469 31875
rect 6503 31872 6515 31875
rect 7098 31872 7104 31884
rect 6503 31844 7104 31872
rect 6503 31841 6515 31844
rect 6457 31835 6515 31841
rect 7098 31832 7104 31844
rect 7156 31832 7162 31884
rect 8588 31872 8616 31971
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 11149 32011 11207 32017
rect 11149 32008 11161 32011
rect 10192 31980 11161 32008
rect 10192 31968 10198 31980
rect 11149 31977 11161 31980
rect 11195 31977 11207 32011
rect 11149 31971 11207 31977
rect 11606 31968 11612 32020
rect 11664 32008 11670 32020
rect 16393 32011 16451 32017
rect 16393 32008 16405 32011
rect 11664 31980 16405 32008
rect 11664 31968 11670 31980
rect 16393 31977 16405 31980
rect 16439 31977 16451 32011
rect 16393 31971 16451 31977
rect 17954 31968 17960 32020
rect 18012 32008 18018 32020
rect 18049 32011 18107 32017
rect 18049 32008 18061 32011
rect 18012 31980 18061 32008
rect 18012 31968 18018 31980
rect 18049 31977 18061 31980
rect 18095 32008 18107 32011
rect 18414 32008 18420 32020
rect 18095 31980 18420 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18414 31968 18420 31980
rect 18472 31968 18478 32020
rect 19352 31980 20852 32008
rect 9214 31900 9220 31952
rect 9272 31940 9278 31952
rect 9272 31912 9536 31940
rect 9272 31900 9278 31912
rect 7576 31844 8616 31872
rect 9508 31872 9536 31912
rect 11238 31900 11244 31952
rect 11296 31940 11302 31952
rect 13909 31943 13967 31949
rect 13909 31940 13921 31943
rect 11296 31912 13921 31940
rect 11296 31900 11302 31912
rect 13909 31909 13921 31912
rect 13955 31940 13967 31943
rect 14090 31940 14096 31952
rect 13955 31912 14096 31940
rect 13955 31909 13967 31912
rect 13909 31903 13967 31909
rect 14090 31900 14096 31912
rect 14148 31900 14154 31952
rect 14274 31900 14280 31952
rect 14332 31900 14338 31952
rect 14642 31900 14648 31952
rect 14700 31940 14706 31952
rect 15102 31940 15108 31952
rect 14700 31912 15108 31940
rect 14700 31900 14706 31912
rect 15102 31900 15108 31912
rect 15160 31940 15166 31952
rect 15930 31940 15936 31952
rect 15160 31912 15936 31940
rect 15160 31900 15166 31912
rect 15930 31900 15936 31912
rect 15988 31900 15994 31952
rect 16114 31900 16120 31952
rect 16172 31940 16178 31952
rect 19352 31940 19380 31980
rect 16172 31912 19380 31940
rect 16172 31900 16178 31912
rect 19426 31900 19432 31952
rect 19484 31900 19490 31952
rect 19536 31912 20116 31940
rect 9677 31875 9735 31881
rect 9677 31872 9689 31875
rect 9508 31844 9689 31872
rect 7576 31790 7604 31844
rect 9677 31841 9689 31844
rect 9723 31872 9735 31875
rect 9723 31844 10916 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 8294 31764 8300 31816
rect 8352 31764 8358 31816
rect 9390 31807 9448 31813
rect 9390 31804 9402 31807
rect 9324 31776 9402 31804
rect 9324 31736 9352 31776
rect 9390 31773 9402 31776
rect 9436 31773 9448 31807
rect 10888 31804 10916 31844
rect 11422 31832 11428 31884
rect 11480 31872 11486 31884
rect 13633 31875 13691 31881
rect 13633 31872 13645 31875
rect 11480 31844 13645 31872
rect 11480 31832 11486 31844
rect 13633 31841 13645 31844
rect 13679 31872 13691 31875
rect 13814 31872 13820 31884
rect 13679 31844 13820 31872
rect 13679 31841 13691 31844
rect 13633 31835 13691 31841
rect 13814 31832 13820 31844
rect 13872 31832 13878 31884
rect 14108 31872 14136 31900
rect 14829 31875 14887 31881
rect 14829 31872 14841 31875
rect 14108 31844 14841 31872
rect 14829 31841 14841 31844
rect 14875 31841 14887 31875
rect 16945 31875 17003 31881
rect 16945 31872 16957 31875
rect 14829 31835 14887 31841
rect 14936 31844 16957 31872
rect 14642 31804 14648 31816
rect 10888 31776 14648 31804
rect 9390 31767 9448 31773
rect 14642 31764 14648 31776
rect 14700 31764 14706 31816
rect 14734 31764 14740 31816
rect 14792 31764 14798 31816
rect 14936 31804 14964 31844
rect 16945 31841 16957 31844
rect 16991 31841 17003 31875
rect 16945 31835 17003 31841
rect 18230 31832 18236 31884
rect 18288 31832 18294 31884
rect 19150 31832 19156 31884
rect 19208 31872 19214 31884
rect 19536 31872 19564 31912
rect 19208 31844 19564 31872
rect 19208 31832 19214 31844
rect 19978 31832 19984 31884
rect 20036 31832 20042 31884
rect 20088 31872 20116 31912
rect 20254 31900 20260 31952
rect 20312 31940 20318 31952
rect 20625 31943 20683 31949
rect 20625 31940 20637 31943
rect 20312 31912 20637 31940
rect 20312 31900 20318 31912
rect 20625 31909 20637 31912
rect 20671 31909 20683 31943
rect 20824 31940 20852 31980
rect 20898 31968 20904 32020
rect 20956 32008 20962 32020
rect 23290 32008 23296 32020
rect 20956 31980 23296 32008
rect 20956 31968 20962 31980
rect 23290 31968 23296 31980
rect 23348 31968 23354 32020
rect 24210 31968 24216 32020
rect 24268 32008 24274 32020
rect 25133 32011 25191 32017
rect 25133 32008 25145 32011
rect 24268 31980 25145 32008
rect 24268 31968 24274 31980
rect 25133 31977 25145 31980
rect 25179 31977 25191 32011
rect 25133 31971 25191 31977
rect 21634 31940 21640 31952
rect 20824 31912 21640 31940
rect 20625 31903 20683 31909
rect 21634 31900 21640 31912
rect 21692 31900 21698 31952
rect 21913 31943 21971 31949
rect 21913 31909 21925 31943
rect 21959 31940 21971 31943
rect 23382 31940 23388 31952
rect 21959 31912 23388 31940
rect 21959 31909 21971 31912
rect 21913 31903 21971 31909
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 20088 31844 21189 31872
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 21177 31835 21235 31841
rect 21358 31832 21364 31884
rect 21416 31872 21422 31884
rect 22373 31875 22431 31881
rect 22373 31872 22385 31875
rect 21416 31844 22385 31872
rect 21416 31832 21422 31844
rect 22373 31841 22385 31844
rect 22419 31841 22431 31875
rect 22373 31835 22431 31841
rect 22557 31875 22615 31881
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23474 31872 23480 31884
rect 22603 31844 23480 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23474 31832 23480 31844
rect 23532 31832 23538 31884
rect 14844 31776 14964 31804
rect 16853 31807 16911 31813
rect 9582 31736 9588 31748
rect 9324 31708 9588 31736
rect 9582 31696 9588 31708
rect 9640 31696 9646 31748
rect 10134 31736 10140 31748
rect 10060 31708 10140 31736
rect 7374 31628 7380 31680
rect 7432 31668 7438 31680
rect 8294 31668 8300 31680
rect 7432 31640 8300 31668
rect 7432 31628 7438 31640
rect 8294 31628 8300 31640
rect 8352 31628 8358 31680
rect 9122 31628 9128 31680
rect 9180 31628 9186 31680
rect 10060 31668 10088 31708
rect 10134 31696 10140 31708
rect 10192 31696 10198 31748
rect 14458 31696 14464 31748
rect 14516 31736 14522 31748
rect 14844 31736 14872 31776
rect 16853 31773 16865 31807
rect 16899 31804 16911 31807
rect 17126 31804 17132 31816
rect 16899 31776 17132 31804
rect 16899 31773 16911 31776
rect 16853 31767 16911 31773
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 18046 31764 18052 31816
rect 18104 31804 18110 31816
rect 18417 31807 18475 31813
rect 18417 31804 18429 31807
rect 18104 31776 18429 31804
rect 18104 31764 18110 31776
rect 18417 31773 18429 31776
rect 18463 31804 18475 31807
rect 18874 31804 18880 31816
rect 18463 31776 18880 31804
rect 18463 31773 18475 31776
rect 18417 31767 18475 31773
rect 18874 31764 18880 31776
rect 18932 31764 18938 31816
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31804 19947 31807
rect 20806 31804 20812 31816
rect 19935 31776 20812 31804
rect 19935 31773 19947 31776
rect 19889 31767 19947 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31804 21143 31807
rect 21634 31804 21640 31816
rect 21131 31776 21640 31804
rect 21131 31773 21143 31776
rect 21085 31767 21143 31773
rect 21634 31764 21640 31776
rect 21692 31804 21698 31816
rect 21910 31804 21916 31816
rect 21692 31776 21916 31804
rect 21692 31764 21698 31776
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 24121 31807 24179 31813
rect 24121 31773 24133 31807
rect 24167 31804 24179 31807
rect 24302 31804 24308 31816
rect 24167 31776 24308 31804
rect 24167 31773 24179 31776
rect 24121 31767 24179 31773
rect 24302 31764 24308 31776
rect 24360 31764 24366 31816
rect 24857 31807 24915 31813
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 14516 31708 14872 31736
rect 14516 31696 14522 31708
rect 19794 31696 19800 31748
rect 19852 31696 19858 31748
rect 20993 31739 21051 31745
rect 20993 31705 21005 31739
rect 21039 31736 21051 31739
rect 21174 31736 21180 31748
rect 21039 31708 21180 31736
rect 21039 31705 21051 31708
rect 20993 31699 21051 31705
rect 21174 31696 21180 31708
rect 21232 31696 21238 31748
rect 21266 31696 21272 31748
rect 21324 31736 21330 31748
rect 22281 31739 22339 31745
rect 22281 31736 22293 31739
rect 21324 31708 22293 31736
rect 21324 31696 21330 31708
rect 22281 31705 22293 31708
rect 22327 31705 22339 31739
rect 22281 31699 22339 31705
rect 11425 31671 11483 31677
rect 11425 31668 11437 31671
rect 10060 31640 11437 31668
rect 11425 31637 11437 31640
rect 11471 31637 11483 31671
rect 11425 31631 11483 31637
rect 13814 31628 13820 31680
rect 13872 31668 13878 31680
rect 14645 31671 14703 31677
rect 14645 31668 14657 31671
rect 13872 31640 14657 31668
rect 13872 31628 13878 31640
rect 14645 31637 14657 31640
rect 14691 31668 14703 31671
rect 15010 31668 15016 31680
rect 14691 31640 15016 31668
rect 14691 31637 14703 31640
rect 14645 31631 14703 31637
rect 15010 31628 15016 31640
rect 15068 31628 15074 31680
rect 16761 31671 16819 31677
rect 16761 31637 16773 31671
rect 16807 31668 16819 31671
rect 17678 31668 17684 31680
rect 16807 31640 17684 31668
rect 16807 31637 16819 31640
rect 16761 31631 16819 31637
rect 17678 31628 17684 31640
rect 17736 31628 17742 31680
rect 20070 31628 20076 31680
rect 20128 31668 20134 31680
rect 21450 31668 21456 31680
rect 20128 31640 21456 31668
rect 20128 31628 20134 31640
rect 21450 31628 21456 31640
rect 21508 31628 21514 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 7469 31467 7527 31473
rect 7469 31433 7481 31467
rect 7515 31464 7527 31467
rect 7650 31464 7656 31476
rect 7515 31436 7656 31464
rect 7515 31433 7527 31436
rect 7469 31427 7527 31433
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 8662 31424 8668 31476
rect 8720 31424 8726 31476
rect 9033 31467 9091 31473
rect 9033 31433 9045 31467
rect 9079 31464 9091 31467
rect 9858 31464 9864 31476
rect 9079 31436 9864 31464
rect 9079 31433 9091 31436
rect 9033 31427 9091 31433
rect 9858 31424 9864 31436
rect 9916 31424 9922 31476
rect 13354 31424 13360 31476
rect 13412 31464 13418 31476
rect 18325 31467 18383 31473
rect 18325 31464 18337 31467
rect 13412 31436 18337 31464
rect 13412 31424 13418 31436
rect 18325 31433 18337 31436
rect 18371 31433 18383 31467
rect 18325 31427 18383 31433
rect 18598 31424 18604 31476
rect 18656 31464 18662 31476
rect 18966 31464 18972 31476
rect 18656 31436 18972 31464
rect 18656 31424 18662 31436
rect 18966 31424 18972 31436
rect 19024 31424 19030 31476
rect 20070 31464 20076 31476
rect 19996 31436 20076 31464
rect 9769 31399 9827 31405
rect 9769 31365 9781 31399
rect 9815 31396 9827 31399
rect 11238 31396 11244 31408
rect 9815 31368 11244 31396
rect 9815 31365 9827 31368
rect 9769 31359 9827 31365
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 1946 31328 1952 31340
rect 1811 31300 1952 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 7834 31288 7840 31340
rect 7892 31288 7898 31340
rect 7929 31331 7987 31337
rect 7929 31297 7941 31331
rect 7975 31328 7987 31331
rect 8754 31328 8760 31340
rect 7975 31300 8760 31328
rect 7975 31297 7987 31300
rect 7929 31291 7987 31297
rect 1302 31220 1308 31272
rect 1360 31260 1366 31272
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1360 31232 2053 31260
rect 1360 31220 1366 31232
rect 2041 31229 2053 31232
rect 2087 31229 2099 31263
rect 2041 31223 2099 31229
rect 5626 31220 5632 31272
rect 5684 31260 5690 31272
rect 7193 31263 7251 31269
rect 7193 31260 7205 31263
rect 5684 31232 7205 31260
rect 5684 31220 5690 31232
rect 7193 31229 7205 31232
rect 7239 31260 7251 31263
rect 7944 31260 7972 31291
rect 8754 31288 8760 31300
rect 8812 31288 8818 31340
rect 9784 31328 9812 31359
rect 11238 31356 11244 31368
rect 11296 31356 11302 31408
rect 14921 31399 14979 31405
rect 14921 31396 14933 31399
rect 14398 31368 14933 31396
rect 14921 31365 14933 31368
rect 14967 31396 14979 31399
rect 15102 31396 15108 31408
rect 14967 31368 15108 31396
rect 14967 31365 14979 31368
rect 14921 31359 14979 31365
rect 15102 31356 15108 31368
rect 15160 31356 15166 31408
rect 18414 31356 18420 31408
rect 18472 31396 18478 31408
rect 18782 31396 18788 31408
rect 18472 31368 18788 31396
rect 18472 31356 18478 31368
rect 18782 31356 18788 31368
rect 18840 31356 18846 31408
rect 9324 31300 9812 31328
rect 17497 31331 17555 31337
rect 7239 31232 7972 31260
rect 7239 31229 7251 31232
rect 7193 31223 7251 31229
rect 8110 31220 8116 31272
rect 8168 31220 8174 31272
rect 8478 31220 8484 31272
rect 8536 31260 8542 31272
rect 9324 31269 9352 31300
rect 17497 31297 17509 31331
rect 17543 31297 17555 31331
rect 17497 31291 17555 31297
rect 17589 31331 17647 31337
rect 17589 31297 17601 31331
rect 17635 31328 17647 31331
rect 18322 31328 18328 31340
rect 17635 31300 18328 31328
rect 17635 31297 17647 31300
rect 17589 31291 17647 31297
rect 9125 31263 9183 31269
rect 9125 31260 9137 31263
rect 8536 31232 9137 31260
rect 8536 31220 8542 31232
rect 9125 31229 9137 31232
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9309 31263 9367 31269
rect 9309 31229 9321 31263
rect 9355 31229 9367 31263
rect 9309 31223 9367 31229
rect 9582 31220 9588 31272
rect 9640 31260 9646 31272
rect 12897 31263 12955 31269
rect 12897 31260 12909 31263
rect 9640 31232 12909 31260
rect 9640 31220 9646 31232
rect 12897 31229 12909 31232
rect 12943 31260 12955 31263
rect 13173 31263 13231 31269
rect 12943 31232 13032 31260
rect 12943 31229 12955 31232
rect 12897 31223 12955 31229
rect 5902 31152 5908 31204
rect 5960 31192 5966 31204
rect 8496 31192 8524 31220
rect 5960 31164 8524 31192
rect 5960 31152 5966 31164
rect 13004 31124 13032 31232
rect 13173 31229 13185 31263
rect 13219 31260 13231 31263
rect 13262 31260 13268 31272
rect 13219 31232 13268 31260
rect 13219 31229 13231 31232
rect 13173 31223 13231 31229
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 14918 31220 14924 31272
rect 14976 31260 14982 31272
rect 16761 31263 16819 31269
rect 16761 31260 16773 31263
rect 14976 31232 16773 31260
rect 14976 31220 14982 31232
rect 16761 31229 16773 31232
rect 16807 31260 16819 31263
rect 17512 31260 17540 31291
rect 18322 31288 18328 31300
rect 18380 31288 18386 31340
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31328 18751 31331
rect 18966 31328 18972 31340
rect 18739 31300 18972 31328
rect 18739 31297 18751 31300
rect 18693 31291 18751 31297
rect 18966 31288 18972 31300
rect 19024 31288 19030 31340
rect 19889 31331 19947 31337
rect 19889 31328 19901 31331
rect 19076 31300 19901 31328
rect 16807 31232 17540 31260
rect 17773 31263 17831 31269
rect 16807 31229 16819 31232
rect 16761 31223 16819 31229
rect 17773 31229 17785 31263
rect 17819 31260 17831 31263
rect 17862 31260 17868 31272
rect 17819 31232 17868 31260
rect 17819 31229 17831 31232
rect 17773 31223 17831 31229
rect 17862 31220 17868 31232
rect 17920 31220 17926 31272
rect 18782 31220 18788 31272
rect 18840 31220 18846 31272
rect 18874 31220 18880 31272
rect 18932 31220 18938 31272
rect 15470 31192 15476 31204
rect 14660 31164 15476 31192
rect 14660 31136 14688 31164
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 19076 31192 19104 31300
rect 19889 31297 19901 31300
rect 19935 31297 19947 31331
rect 19889 31291 19947 31297
rect 19334 31220 19340 31272
rect 19392 31260 19398 31272
rect 19996 31269 20024 31436
rect 20070 31424 20076 31436
rect 20128 31464 20134 31476
rect 20717 31467 20775 31473
rect 20717 31464 20729 31467
rect 20128 31436 20729 31464
rect 20128 31424 20134 31436
rect 20717 31433 20729 31436
rect 20763 31433 20775 31467
rect 20717 31427 20775 31433
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 21634 31464 21640 31476
rect 21591 31436 21640 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 21634 31424 21640 31436
rect 21692 31424 21698 31476
rect 22646 31464 22652 31476
rect 22066 31436 22652 31464
rect 22066 31396 22094 31436
rect 22646 31424 22652 31436
rect 22704 31424 22710 31476
rect 23934 31424 23940 31476
rect 23992 31464 23998 31476
rect 25133 31467 25191 31473
rect 25133 31464 25145 31467
rect 23992 31436 25145 31464
rect 23992 31424 23998 31436
rect 25133 31433 25145 31436
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 22465 31399 22523 31405
rect 22465 31396 22477 31399
rect 20640 31368 22094 31396
rect 22204 31368 22477 31396
rect 20640 31272 20668 31368
rect 21818 31288 21824 31340
rect 21876 31328 21882 31340
rect 22204 31328 22232 31368
rect 22465 31365 22477 31368
rect 22511 31365 22523 31399
rect 24302 31396 24308 31408
rect 23690 31368 24308 31396
rect 22465 31359 22523 31365
rect 24302 31356 24308 31368
rect 24360 31356 24366 31408
rect 21876 31300 22232 31328
rect 21876 31288 21882 31300
rect 24394 31288 24400 31340
rect 24452 31328 24458 31340
rect 24581 31331 24639 31337
rect 24581 31328 24593 31331
rect 24452 31300 24593 31328
rect 24452 31288 24458 31300
rect 24581 31297 24593 31300
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 25314 31288 25320 31340
rect 25372 31288 25378 31340
rect 19981 31263 20039 31269
rect 19981 31260 19993 31263
rect 19392 31232 19993 31260
rect 19392 31220 19398 31232
rect 19981 31229 19993 31232
rect 20027 31229 20039 31263
rect 19981 31223 20039 31229
rect 20165 31263 20223 31269
rect 20165 31229 20177 31263
rect 20211 31260 20223 31263
rect 20622 31260 20628 31272
rect 20211 31232 20628 31260
rect 20211 31229 20223 31232
rect 20165 31223 20223 31229
rect 20622 31220 20628 31232
rect 20680 31220 20686 31272
rect 22186 31220 22192 31272
rect 22244 31220 22250 31272
rect 17052 31164 19104 31192
rect 14458 31124 14464 31136
rect 13004 31096 14464 31124
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 14642 31084 14648 31136
rect 14700 31084 14706 31136
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 17052 31124 17080 31164
rect 15344 31096 17080 31124
rect 15344 31084 15350 31096
rect 17126 31084 17132 31136
rect 17184 31084 17190 31136
rect 19076 31124 19104 31164
rect 19521 31195 19579 31201
rect 19521 31161 19533 31195
rect 19567 31192 19579 31195
rect 21910 31192 21916 31204
rect 19567 31164 21916 31192
rect 19567 31161 19579 31164
rect 19521 31155 19579 31161
rect 21910 31152 21916 31164
rect 21968 31152 21974 31204
rect 20533 31127 20591 31133
rect 20533 31124 20545 31127
rect 19076 31096 20545 31124
rect 20533 31093 20545 31096
rect 20579 31093 20591 31127
rect 20533 31087 20591 31093
rect 23566 31084 23572 31136
rect 23624 31124 23630 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23624 31096 23949 31124
rect 23624 31084 23630 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 23937 31087 23995 31093
rect 24397 31127 24455 31133
rect 24397 31093 24409 31127
rect 24443 31124 24455 31127
rect 24486 31124 24492 31136
rect 24443 31096 24492 31124
rect 24443 31093 24455 31096
rect 24397 31087 24455 31093
rect 24486 31084 24492 31096
rect 24544 31084 24550 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 8110 30880 8116 30932
rect 8168 30920 8174 30932
rect 8168 30892 11284 30920
rect 8168 30880 8174 30892
rect 11256 30852 11284 30892
rect 11974 30880 11980 30932
rect 12032 30920 12038 30932
rect 12805 30923 12863 30929
rect 12805 30920 12817 30923
rect 12032 30892 12817 30920
rect 12032 30880 12038 30892
rect 12805 30889 12817 30892
rect 12851 30889 12863 30923
rect 18506 30920 18512 30932
rect 12805 30883 12863 30889
rect 14660 30892 18512 30920
rect 12437 30855 12495 30861
rect 12437 30852 12449 30855
rect 11256 30824 12449 30852
rect 12437 30821 12449 30824
rect 12483 30852 12495 30855
rect 12483 30824 13400 30852
rect 12483 30821 12495 30824
rect 12437 30815 12495 30821
rect 1670 30744 1676 30796
rect 1728 30784 1734 30796
rect 3973 30787 4031 30793
rect 3973 30784 3985 30787
rect 1728 30756 3985 30784
rect 1728 30744 1734 30756
rect 3973 30753 3985 30756
rect 4019 30753 4031 30787
rect 3973 30747 4031 30753
rect 7834 30744 7840 30796
rect 7892 30784 7898 30796
rect 7929 30787 7987 30793
rect 7929 30784 7941 30787
rect 7892 30756 7941 30784
rect 7892 30744 7898 30756
rect 7929 30753 7941 30756
rect 7975 30753 7987 30787
rect 7929 30747 7987 30753
rect 9582 30744 9588 30796
rect 9640 30744 9646 30796
rect 9861 30787 9919 30793
rect 9861 30753 9873 30787
rect 9907 30784 9919 30787
rect 10594 30784 10600 30796
rect 9907 30756 10600 30784
rect 9907 30753 9919 30756
rect 9861 30747 9919 30753
rect 10594 30744 10600 30756
rect 10652 30744 10658 30796
rect 13372 30793 13400 30824
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30753 13415 30787
rect 13357 30747 13415 30753
rect 11422 30676 11428 30728
rect 11480 30716 11486 30728
rect 12253 30719 12311 30725
rect 12253 30716 12265 30719
rect 11480 30688 12265 30716
rect 11480 30676 11486 30688
rect 12253 30685 12265 30688
rect 12299 30716 12311 30719
rect 13173 30719 13231 30725
rect 13173 30716 13185 30719
rect 12299 30688 13185 30716
rect 12299 30685 12311 30688
rect 12253 30679 12311 30685
rect 13173 30685 13185 30688
rect 13219 30716 13231 30719
rect 14660 30716 14688 30892
rect 18506 30880 18512 30892
rect 18564 30880 18570 30932
rect 20438 30920 20444 30932
rect 19904 30892 20444 30920
rect 15194 30744 15200 30796
rect 15252 30784 15258 30796
rect 16209 30787 16267 30793
rect 16209 30784 16221 30787
rect 15252 30756 16221 30784
rect 15252 30744 15258 30756
rect 16209 30753 16221 30756
rect 16255 30753 16267 30787
rect 16209 30747 16267 30753
rect 16482 30744 16488 30796
rect 16540 30784 16546 30796
rect 18874 30784 18880 30796
rect 16540 30756 18880 30784
rect 16540 30744 16546 30756
rect 18874 30744 18880 30756
rect 18932 30784 18938 30796
rect 19904 30793 19932 30892
rect 20438 30880 20444 30892
rect 20496 30880 20502 30932
rect 20530 30880 20536 30932
rect 20588 30920 20594 30932
rect 20588 30892 22692 30920
rect 20588 30880 20594 30892
rect 19889 30787 19947 30793
rect 18932 30756 19334 30784
rect 18932 30744 18938 30756
rect 13219 30688 14688 30716
rect 13219 30685 13231 30688
rect 13173 30679 13231 30685
rect 17494 30676 17500 30728
rect 17552 30716 17558 30728
rect 18233 30719 18291 30725
rect 18233 30716 18245 30719
rect 17552 30688 18245 30716
rect 17552 30676 17558 30688
rect 18233 30685 18245 30688
rect 18279 30685 18291 30719
rect 19306 30716 19334 30756
rect 19889 30753 19901 30787
rect 19935 30753 19947 30787
rect 19889 30747 19947 30753
rect 19978 30744 19984 30796
rect 20036 30744 20042 30796
rect 20438 30744 20444 30796
rect 20496 30784 20502 30796
rect 22557 30787 22615 30793
rect 22557 30784 22569 30787
rect 20496 30756 22569 30784
rect 20496 30744 20502 30756
rect 22557 30753 22569 30756
rect 22603 30753 22615 30787
rect 22664 30784 22692 30892
rect 22830 30880 22836 30932
rect 22888 30920 22894 30932
rect 23017 30923 23075 30929
rect 23017 30920 23029 30923
rect 22888 30892 23029 30920
rect 22888 30880 22894 30892
rect 23017 30889 23029 30892
rect 23063 30889 23075 30923
rect 23017 30883 23075 30889
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25314 30920 25320 30932
rect 24903 30892 25320 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25314 30880 25320 30892
rect 25372 30880 25378 30932
rect 25133 30855 25191 30861
rect 25133 30821 25145 30855
rect 25179 30821 25191 30855
rect 25133 30815 25191 30821
rect 25148 30784 25176 30815
rect 22664 30756 25176 30784
rect 22557 30747 22615 30753
rect 19426 30716 19432 30728
rect 19306 30688 19432 30716
rect 18233 30679 18291 30685
rect 19426 30676 19432 30688
rect 19484 30676 19490 30728
rect 19702 30676 19708 30728
rect 19760 30716 19766 30728
rect 19797 30719 19855 30725
rect 19797 30716 19809 30719
rect 19760 30688 19809 30716
rect 19760 30676 19766 30688
rect 19797 30685 19809 30688
rect 19843 30685 19855 30719
rect 19797 30679 19855 30685
rect 22278 30676 22284 30728
rect 22336 30716 22342 30728
rect 23845 30719 23903 30725
rect 23845 30716 23857 30719
rect 22336 30688 23857 30716
rect 22336 30676 22342 30688
rect 23845 30685 23857 30688
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25498 30716 25504 30728
rect 25363 30688 25504 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 25498 30676 25504 30688
rect 25556 30676 25562 30728
rect 3786 30608 3792 30660
rect 3844 30648 3850 30660
rect 4157 30651 4215 30657
rect 4157 30648 4169 30651
rect 3844 30620 4169 30648
rect 3844 30608 3850 30620
rect 4157 30617 4169 30620
rect 4203 30617 4215 30651
rect 4157 30611 4215 30617
rect 5813 30651 5871 30657
rect 5813 30617 5825 30651
rect 5859 30648 5871 30651
rect 5902 30648 5908 30660
rect 5859 30620 5908 30648
rect 5859 30617 5871 30620
rect 5813 30611 5871 30617
rect 5902 30608 5908 30620
rect 5960 30608 5966 30660
rect 11609 30651 11667 30657
rect 11609 30648 11621 30651
rect 10244 30620 10350 30648
rect 11256 30620 11621 30648
rect 10244 30592 10272 30620
rect 8478 30540 8484 30592
rect 8536 30540 8542 30592
rect 10226 30540 10232 30592
rect 10284 30580 10290 30592
rect 11256 30580 11284 30620
rect 11609 30617 11621 30620
rect 11655 30617 11667 30651
rect 11609 30611 11667 30617
rect 13265 30651 13323 30657
rect 13265 30617 13277 30651
rect 13311 30648 13323 30651
rect 13909 30651 13967 30657
rect 13909 30648 13921 30651
rect 13311 30620 13921 30648
rect 13311 30617 13323 30620
rect 13265 30611 13323 30617
rect 13909 30617 13921 30620
rect 13955 30648 13967 30651
rect 16574 30648 16580 30660
rect 13955 30620 16580 30648
rect 13955 30617 13967 30620
rect 13909 30611 13967 30617
rect 16574 30608 16580 30620
rect 16632 30608 16638 30660
rect 16684 30620 16974 30648
rect 10284 30552 11284 30580
rect 10284 30540 10290 30552
rect 11330 30540 11336 30592
rect 11388 30540 11394 30592
rect 15102 30540 15108 30592
rect 15160 30580 15166 30592
rect 15841 30583 15899 30589
rect 15841 30580 15853 30583
rect 15160 30552 15853 30580
rect 15160 30540 15166 30552
rect 15841 30549 15853 30552
rect 15887 30580 15899 30583
rect 16684 30580 16712 30620
rect 18782 30608 18788 30660
rect 18840 30648 18846 30660
rect 22373 30651 22431 30657
rect 22373 30648 22385 30651
rect 18840 30620 22385 30648
rect 18840 30608 18846 30620
rect 22373 30617 22385 30620
rect 22419 30648 22431 30651
rect 24762 30648 24768 30660
rect 22419 30620 24768 30648
rect 22419 30617 22431 30620
rect 22373 30611 22431 30617
rect 24762 30608 24768 30620
rect 24820 30608 24826 30660
rect 17402 30580 17408 30592
rect 15887 30552 17408 30580
rect 15887 30549 15899 30552
rect 15841 30543 15899 30549
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 17494 30540 17500 30592
rect 17552 30580 17558 30592
rect 17770 30580 17776 30592
rect 17552 30552 17776 30580
rect 17552 30540 17558 30552
rect 17770 30540 17776 30552
rect 17828 30580 17834 30592
rect 17957 30583 18015 30589
rect 17957 30580 17969 30583
rect 17828 30552 17969 30580
rect 17828 30540 17834 30552
rect 17957 30549 17969 30552
rect 18003 30549 18015 30583
rect 17957 30543 18015 30549
rect 18598 30540 18604 30592
rect 18656 30580 18662 30592
rect 19150 30580 19156 30592
rect 18656 30552 19156 30580
rect 18656 30540 18662 30552
rect 19150 30540 19156 30552
rect 19208 30540 19214 30592
rect 19426 30540 19432 30592
rect 19484 30540 19490 30592
rect 21818 30540 21824 30592
rect 21876 30580 21882 30592
rect 22005 30583 22063 30589
rect 22005 30580 22017 30583
rect 21876 30552 22017 30580
rect 21876 30540 21882 30552
rect 22005 30549 22017 30552
rect 22051 30549 22063 30583
rect 22005 30543 22063 30549
rect 22465 30583 22523 30589
rect 22465 30549 22477 30583
rect 22511 30580 22523 30583
rect 22830 30580 22836 30592
rect 22511 30552 22836 30580
rect 22511 30549 22523 30552
rect 22465 30543 22523 30549
rect 22830 30540 22836 30552
rect 22888 30540 22894 30592
rect 23661 30583 23719 30589
rect 23661 30549 23673 30583
rect 23707 30580 23719 30583
rect 24946 30580 24952 30592
rect 23707 30552 24952 30580
rect 23707 30549 23719 30552
rect 23661 30543 23719 30549
rect 24946 30540 24952 30552
rect 25004 30540 25010 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 15120 30348 16068 30376
rect 6362 30268 6368 30320
rect 6420 30308 6426 30320
rect 8941 30311 8999 30317
rect 8941 30308 8953 30311
rect 6420 30280 8953 30308
rect 6420 30268 6426 30280
rect 8941 30277 8953 30280
rect 8987 30308 8999 30311
rect 9582 30308 9588 30320
rect 8987 30280 9588 30308
rect 8987 30277 8999 30280
rect 8941 30271 8999 30277
rect 9582 30268 9588 30280
rect 9640 30268 9646 30320
rect 11790 30268 11796 30320
rect 11848 30308 11854 30320
rect 12529 30311 12587 30317
rect 12529 30308 12541 30311
rect 11848 30280 12541 30308
rect 11848 30268 11854 30280
rect 12529 30277 12541 30280
rect 12575 30308 12587 30311
rect 14274 30308 14280 30320
rect 12575 30280 14280 30308
rect 12575 30277 12587 30280
rect 12529 30271 12587 30277
rect 14274 30268 14280 30280
rect 14332 30268 14338 30320
rect 15120 30308 15148 30348
rect 14384 30280 15148 30308
rect 14384 30252 14412 30280
rect 15194 30268 15200 30320
rect 15252 30268 15258 30320
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 10827 30212 11713 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 14366 30240 14372 30252
rect 11701 30203 11759 30209
rect 12406 30212 14372 30240
rect 10137 30175 10195 30181
rect 10137 30141 10149 30175
rect 10183 30172 10195 30175
rect 10502 30172 10508 30184
rect 10183 30144 10508 30172
rect 10183 30141 10195 30144
rect 10137 30135 10195 30141
rect 10502 30132 10508 30144
rect 10560 30172 10566 30184
rect 10686 30172 10692 30184
rect 10560 30144 10692 30172
rect 10560 30132 10566 30144
rect 10686 30132 10692 30144
rect 10744 30172 10750 30184
rect 10873 30175 10931 30181
rect 10873 30172 10885 30175
rect 10744 30144 10885 30172
rect 10744 30132 10750 30144
rect 10873 30141 10885 30144
rect 10919 30141 10931 30175
rect 10873 30135 10931 30141
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30141 11023 30175
rect 10965 30135 11023 30141
rect 10594 30064 10600 30116
rect 10652 30104 10658 30116
rect 10980 30104 11008 30135
rect 10652 30076 11008 30104
rect 10652 30064 10658 30076
rect 10410 29996 10416 30048
rect 10468 29996 10474 30048
rect 11882 29996 11888 30048
rect 11940 30036 11946 30048
rect 12253 30039 12311 30045
rect 12253 30036 12265 30039
rect 11940 30008 12265 30036
rect 11940 29996 11946 30008
rect 12253 30005 12265 30008
rect 12299 30036 12311 30039
rect 12406 30036 12434 30212
rect 14366 30200 14372 30212
rect 14424 30200 14430 30252
rect 14458 30200 14464 30252
rect 14516 30200 14522 30252
rect 16040 30240 16068 30348
rect 18322 30336 18328 30388
rect 18380 30376 18386 30388
rect 19150 30376 19156 30388
rect 18380 30348 19156 30376
rect 18380 30336 18386 30348
rect 19150 30336 19156 30348
rect 19208 30336 19214 30388
rect 19334 30336 19340 30388
rect 19392 30376 19398 30388
rect 20898 30376 20904 30388
rect 19392 30348 20904 30376
rect 19392 30336 19398 30348
rect 20898 30336 20904 30348
rect 20956 30336 20962 30388
rect 24302 30336 24308 30388
rect 24360 30376 24366 30388
rect 24360 30348 24992 30376
rect 24360 30336 24366 30348
rect 17586 30268 17592 30320
rect 17644 30308 17650 30320
rect 17644 30280 19288 30308
rect 17644 30268 17650 30280
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 16040 30212 17969 30240
rect 17957 30209 17969 30212
rect 18003 30240 18015 30243
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 18003 30212 18613 30240
rect 18003 30209 18015 30212
rect 17957 30203 18015 30209
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 19260 30240 19288 30280
rect 23566 30268 23572 30320
rect 23624 30308 23630 30320
rect 23661 30311 23719 30317
rect 23661 30308 23673 30311
rect 23624 30280 23673 30308
rect 23624 30268 23630 30280
rect 23661 30277 23673 30280
rect 23707 30277 23719 30311
rect 24964 30308 24992 30348
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 24886 30280 25421 30308
rect 23661 30271 23719 30277
rect 25409 30277 25421 30280
rect 25455 30277 25467 30311
rect 25409 30271 25467 30277
rect 19613 30243 19671 30249
rect 19613 30240 19625 30243
rect 19260 30212 19625 30240
rect 18601 30203 18659 30209
rect 19613 30209 19625 30212
rect 19659 30209 19671 30243
rect 19613 30203 19671 30209
rect 20162 30200 20168 30252
rect 20220 30240 20226 30252
rect 20346 30240 20352 30252
rect 20220 30212 20352 30240
rect 20220 30200 20226 30212
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 22186 30200 22192 30252
rect 22244 30240 22250 30252
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22244 30212 23397 30240
rect 22244 30200 22250 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 14826 30132 14832 30184
rect 14884 30172 14890 30184
rect 16206 30172 16212 30184
rect 14884 30144 16212 30172
rect 14884 30132 14890 30144
rect 16206 30132 16212 30144
rect 16264 30132 16270 30184
rect 16945 30175 17003 30181
rect 16945 30141 16957 30175
rect 16991 30172 17003 30175
rect 17218 30172 17224 30184
rect 16991 30144 17224 30172
rect 16991 30141 17003 30144
rect 16945 30135 17003 30141
rect 17218 30132 17224 30144
rect 17276 30132 17282 30184
rect 18046 30132 18052 30184
rect 18104 30132 18110 30184
rect 18233 30175 18291 30181
rect 18233 30141 18245 30175
rect 18279 30172 18291 30175
rect 19886 30172 19892 30184
rect 18279 30144 19892 30172
rect 18279 30141 18291 30144
rect 18233 30135 18291 30141
rect 19886 30132 19892 30144
rect 19944 30132 19950 30184
rect 23750 30132 23756 30184
rect 23808 30172 23814 30184
rect 25133 30175 25191 30181
rect 25133 30172 25145 30175
rect 23808 30144 25145 30172
rect 23808 30132 23814 30144
rect 25133 30141 25145 30144
rect 25179 30141 25191 30175
rect 25133 30135 25191 30141
rect 15746 30064 15752 30116
rect 15804 30104 15810 30116
rect 21542 30104 21548 30116
rect 15804 30076 21548 30104
rect 15804 30064 15810 30076
rect 21542 30064 21548 30076
rect 21600 30064 21606 30116
rect 12299 30008 12434 30036
rect 14724 30039 14782 30045
rect 12299 30005 12311 30008
rect 12253 29999 12311 30005
rect 14724 30005 14736 30039
rect 14770 30036 14782 30039
rect 17494 30036 17500 30048
rect 14770 30008 17500 30036
rect 14770 30005 14782 30008
rect 14724 29999 14782 30005
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 17586 29996 17592 30048
rect 17644 29996 17650 30048
rect 18046 29996 18052 30048
rect 18104 30036 18110 30048
rect 18506 30036 18512 30048
rect 18104 30008 18512 30036
rect 18104 29996 18110 30008
rect 18506 29996 18512 30008
rect 18564 30036 18570 30048
rect 18785 30039 18843 30045
rect 18785 30036 18797 30039
rect 18564 30008 18797 30036
rect 18564 29996 18570 30008
rect 18785 30005 18797 30008
rect 18831 30005 18843 30039
rect 18785 29999 18843 30005
rect 18874 29996 18880 30048
rect 18932 30036 18938 30048
rect 19334 30036 19340 30048
rect 18932 30008 19340 30036
rect 18932 29996 18938 30008
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 19429 30039 19487 30045
rect 19429 30005 19441 30039
rect 19475 30036 19487 30039
rect 21726 30036 21732 30048
rect 19475 30008 21732 30036
rect 19475 30005 19487 30008
rect 19429 29999 19487 30005
rect 21726 29996 21732 30008
rect 21784 29996 21790 30048
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 4246 29792 4252 29844
rect 4304 29832 4310 29844
rect 7285 29835 7343 29841
rect 7285 29832 7297 29835
rect 4304 29804 7297 29832
rect 4304 29792 4310 29804
rect 7285 29801 7297 29804
rect 7331 29832 7343 29835
rect 7650 29832 7656 29844
rect 7331 29804 7656 29832
rect 7331 29801 7343 29804
rect 7285 29795 7343 29801
rect 7650 29792 7656 29804
rect 7708 29792 7714 29844
rect 7742 29792 7748 29844
rect 7800 29832 7806 29844
rect 7837 29835 7895 29841
rect 7837 29832 7849 29835
rect 7800 29804 7849 29832
rect 7800 29792 7806 29804
rect 7837 29801 7849 29804
rect 7883 29801 7895 29835
rect 7837 29795 7895 29801
rect 9490 29792 9496 29844
rect 9548 29792 9554 29844
rect 12894 29792 12900 29844
rect 12952 29832 12958 29844
rect 13725 29835 13783 29841
rect 13725 29832 13737 29835
rect 12952 29804 13737 29832
rect 12952 29792 12958 29804
rect 13725 29801 13737 29804
rect 13771 29832 13783 29835
rect 13771 29804 15240 29832
rect 13771 29801 13783 29804
rect 13725 29795 13783 29801
rect 11330 29724 11336 29776
rect 11388 29764 11394 29776
rect 12621 29767 12679 29773
rect 11388 29736 12434 29764
rect 11388 29724 11394 29736
rect 1578 29656 1584 29708
rect 1636 29696 1642 29708
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 1636 29668 4261 29696
rect 1636 29656 1642 29668
rect 4249 29665 4261 29668
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 8389 29699 8447 29705
rect 8389 29696 8401 29699
rect 7156 29668 8401 29696
rect 7156 29656 7162 29668
rect 8389 29665 8401 29668
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 9122 29656 9128 29708
rect 9180 29696 9186 29708
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 9180 29668 9229 29696
rect 9180 29656 9186 29668
rect 9217 29665 9229 29668
rect 9263 29696 9275 29699
rect 10045 29699 10103 29705
rect 10045 29696 10057 29699
rect 9263 29668 10057 29696
rect 9263 29665 9275 29668
rect 9217 29659 9275 29665
rect 10045 29665 10057 29668
rect 10091 29665 10103 29699
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 10045 29659 10103 29665
rect 10152 29668 11989 29696
rect 7282 29588 7288 29640
rect 7340 29588 7346 29640
rect 7834 29588 7840 29640
rect 7892 29628 7898 29640
rect 10152 29628 10180 29668
rect 11977 29665 11989 29668
rect 12023 29665 12035 29699
rect 12406 29696 12434 29736
rect 12621 29733 12633 29767
rect 12667 29764 12679 29767
rect 14734 29764 14740 29776
rect 12667 29736 14740 29764
rect 12667 29733 12679 29736
rect 12621 29727 12679 29733
rect 14734 29724 14740 29736
rect 14792 29724 14798 29776
rect 15212 29764 15240 29804
rect 16022 29792 16028 29844
rect 16080 29832 16086 29844
rect 16482 29832 16488 29844
rect 16080 29804 16488 29832
rect 16080 29792 16086 29804
rect 16482 29792 16488 29804
rect 16540 29792 16546 29844
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 17310 29832 17316 29844
rect 16632 29804 17316 29832
rect 16632 29792 16638 29804
rect 17310 29792 17316 29804
rect 17368 29832 17374 29844
rect 23934 29832 23940 29844
rect 17368 29804 23940 29832
rect 17368 29792 17374 29804
rect 23934 29792 23940 29804
rect 23992 29792 23998 29844
rect 16666 29764 16672 29776
rect 15212 29736 16672 29764
rect 16666 29724 16672 29736
rect 16724 29724 16730 29776
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 21545 29767 21603 29773
rect 17644 29736 20116 29764
rect 17644 29724 17650 29736
rect 13173 29699 13231 29705
rect 13173 29696 13185 29699
rect 12406 29668 13185 29696
rect 11977 29659 12035 29665
rect 13173 29665 13185 29668
rect 13219 29665 13231 29699
rect 13173 29659 13231 29665
rect 14458 29656 14464 29708
rect 14516 29696 14522 29708
rect 17497 29699 17555 29705
rect 17497 29696 17509 29699
rect 14516 29668 17509 29696
rect 14516 29656 14522 29668
rect 17497 29665 17509 29668
rect 17543 29665 17555 29699
rect 17497 29659 17555 29665
rect 18782 29656 18788 29708
rect 18840 29656 18846 29708
rect 20088 29705 20116 29736
rect 21545 29733 21557 29767
rect 21591 29764 21603 29767
rect 24394 29764 24400 29776
rect 21591 29736 24400 29764
rect 21591 29733 21603 29736
rect 21545 29727 21603 29733
rect 24394 29724 24400 29736
rect 24452 29724 24458 29776
rect 20073 29699 20131 29705
rect 20073 29665 20085 29699
rect 20119 29665 20131 29699
rect 20073 29659 20131 29665
rect 20257 29699 20315 29705
rect 20257 29665 20269 29699
rect 20303 29696 20315 29699
rect 21174 29696 21180 29708
rect 20303 29668 21180 29696
rect 20303 29665 20315 29668
rect 20257 29659 20315 29665
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 22189 29699 22247 29705
rect 22189 29665 22201 29699
rect 22235 29696 22247 29699
rect 22554 29696 22560 29708
rect 22235 29668 22560 29696
rect 22235 29665 22247 29668
rect 22189 29659 22247 29665
rect 22554 29656 22560 29668
rect 22612 29656 22618 29708
rect 23382 29656 23388 29708
rect 23440 29656 23446 29708
rect 23569 29699 23627 29705
rect 23569 29665 23581 29699
rect 23615 29696 23627 29699
rect 23750 29696 23756 29708
rect 23615 29668 23756 29696
rect 23615 29665 23627 29668
rect 23569 29659 23627 29665
rect 23750 29656 23756 29668
rect 23808 29656 23814 29708
rect 7892 29600 10180 29628
rect 7892 29588 7898 29600
rect 10410 29588 10416 29640
rect 10468 29628 10474 29640
rect 12989 29631 13047 29637
rect 12989 29628 13001 29631
rect 10468 29600 13001 29628
rect 10468 29588 10474 29600
rect 12989 29597 13001 29600
rect 13035 29597 13047 29631
rect 12989 29591 13047 29597
rect 16390 29588 16396 29640
rect 16448 29628 16454 29640
rect 17405 29631 17463 29637
rect 17405 29628 17417 29631
rect 16448 29600 17417 29628
rect 16448 29588 16454 29600
rect 17405 29597 17417 29600
rect 17451 29597 17463 29631
rect 17405 29591 17463 29597
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29628 20039 29631
rect 20714 29628 20720 29640
rect 20027 29600 20720 29628
rect 20027 29597 20039 29600
rect 19981 29591 20039 29597
rect 20714 29588 20720 29600
rect 20772 29588 20778 29640
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 22002 29628 22008 29640
rect 21959 29600 22008 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 3878 29520 3884 29572
rect 3936 29560 3942 29572
rect 4433 29563 4491 29569
rect 4433 29560 4445 29563
rect 3936 29532 4445 29560
rect 3936 29520 3942 29532
rect 4433 29529 4445 29532
rect 4479 29529 4491 29563
rect 4433 29523 4491 29529
rect 6089 29563 6147 29569
rect 6089 29529 6101 29563
rect 6135 29560 6147 29563
rect 6362 29560 6368 29572
rect 6135 29532 6368 29560
rect 6135 29529 6147 29532
rect 6089 29523 6147 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 7006 29520 7012 29572
rect 7064 29560 7070 29572
rect 7300 29560 7328 29588
rect 7469 29563 7527 29569
rect 7469 29560 7481 29563
rect 7064 29532 7481 29560
rect 7064 29520 7070 29532
rect 7469 29529 7481 29532
rect 7515 29560 7527 29563
rect 8297 29563 8355 29569
rect 8297 29560 8309 29563
rect 7515 29532 8309 29560
rect 7515 29529 7527 29532
rect 7469 29523 7527 29529
rect 8297 29529 8309 29532
rect 8343 29529 8355 29563
rect 8297 29523 8355 29529
rect 9306 29520 9312 29572
rect 9364 29560 9370 29572
rect 9582 29560 9588 29572
rect 9364 29532 9588 29560
rect 9364 29520 9370 29532
rect 9582 29520 9588 29532
rect 9640 29560 9646 29572
rect 9861 29563 9919 29569
rect 9861 29560 9873 29563
rect 9640 29532 9873 29560
rect 9640 29520 9646 29532
rect 9861 29529 9873 29532
rect 9907 29529 9919 29563
rect 9861 29523 9919 29529
rect 11790 29520 11796 29572
rect 11848 29520 11854 29572
rect 12802 29520 12808 29572
rect 12860 29560 12866 29572
rect 13081 29563 13139 29569
rect 13081 29560 13093 29563
rect 12860 29532 13093 29560
rect 12860 29520 12866 29532
rect 13081 29529 13093 29532
rect 13127 29529 13139 29563
rect 13081 29523 13139 29529
rect 14737 29563 14795 29569
rect 14737 29529 14749 29563
rect 14783 29560 14795 29563
rect 16758 29560 16764 29572
rect 14783 29532 16764 29560
rect 14783 29529 14795 29532
rect 14737 29523 14795 29529
rect 16758 29520 16764 29532
rect 16816 29520 16822 29572
rect 17313 29563 17371 29569
rect 17313 29529 17325 29563
rect 17359 29560 17371 29563
rect 17586 29560 17592 29572
rect 17359 29532 17592 29560
rect 17359 29529 17371 29532
rect 17313 29523 17371 29529
rect 17586 29520 17592 29532
rect 17644 29520 17650 29572
rect 18601 29563 18659 29569
rect 18601 29529 18613 29563
rect 18647 29560 18659 29563
rect 20162 29560 20168 29572
rect 18647 29532 20168 29560
rect 18647 29529 18659 29532
rect 18601 29523 18659 29529
rect 20162 29520 20168 29532
rect 20220 29560 20226 29572
rect 20220 29532 25176 29560
rect 20220 29520 20226 29532
rect 7374 29452 7380 29504
rect 7432 29492 7438 29504
rect 7650 29492 7656 29504
rect 7432 29464 7656 29492
rect 7432 29452 7438 29464
rect 7650 29452 7656 29464
rect 7708 29492 7714 29504
rect 8205 29495 8263 29501
rect 8205 29492 8217 29495
rect 7708 29464 8217 29492
rect 7708 29452 7714 29464
rect 8205 29461 8217 29464
rect 8251 29461 8263 29495
rect 8205 29455 8263 29461
rect 9033 29495 9091 29501
rect 9033 29461 9045 29495
rect 9079 29492 9091 29495
rect 9950 29492 9956 29504
rect 9079 29464 9956 29492
rect 9079 29461 9091 29464
rect 9033 29455 9091 29461
rect 9950 29452 9956 29464
rect 10008 29492 10014 29504
rect 10410 29492 10416 29504
rect 10008 29464 10416 29492
rect 10008 29452 10014 29464
rect 10410 29452 10416 29464
rect 10468 29452 10474 29504
rect 10778 29452 10784 29504
rect 10836 29492 10842 29504
rect 11425 29495 11483 29501
rect 11425 29492 11437 29495
rect 10836 29464 11437 29492
rect 10836 29452 10842 29464
rect 11425 29461 11437 29464
rect 11471 29461 11483 29495
rect 11425 29455 11483 29461
rect 11882 29452 11888 29504
rect 11940 29452 11946 29504
rect 13998 29452 14004 29504
rect 14056 29492 14062 29504
rect 14918 29492 14924 29504
rect 14056 29464 14924 29492
rect 14056 29452 14062 29464
rect 14918 29452 14924 29464
rect 14976 29452 14982 29504
rect 16574 29452 16580 29504
rect 16632 29492 16638 29504
rect 16945 29495 17003 29501
rect 16945 29492 16957 29495
rect 16632 29464 16957 29492
rect 16632 29452 16638 29464
rect 16945 29461 16957 29464
rect 16991 29461 17003 29495
rect 16945 29455 17003 29461
rect 17494 29452 17500 29504
rect 17552 29492 17558 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 17552 29464 18153 29492
rect 17552 29452 17558 29464
rect 18141 29461 18153 29464
rect 18187 29461 18199 29495
rect 18141 29455 18199 29461
rect 18322 29452 18328 29504
rect 18380 29492 18386 29504
rect 18509 29495 18567 29501
rect 18509 29492 18521 29495
rect 18380 29464 18521 29492
rect 18380 29452 18386 29464
rect 18509 29461 18521 29464
rect 18555 29461 18567 29495
rect 18509 29455 18567 29461
rect 19613 29495 19671 29501
rect 19613 29461 19625 29495
rect 19659 29492 19671 29495
rect 20346 29492 20352 29504
rect 19659 29464 20352 29492
rect 19659 29461 19671 29464
rect 19613 29455 19671 29461
rect 20346 29452 20352 29464
rect 20404 29452 20410 29504
rect 20898 29452 20904 29504
rect 20956 29452 20962 29504
rect 21910 29452 21916 29504
rect 21968 29492 21974 29504
rect 22005 29495 22063 29501
rect 22005 29492 22017 29495
rect 21968 29464 22017 29492
rect 21968 29452 21974 29464
rect 22005 29461 22017 29464
rect 22051 29461 22063 29495
rect 22005 29455 22063 29461
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22888 29464 22937 29492
rect 22888 29452 22894 29464
rect 22925 29461 22937 29464
rect 22971 29461 22983 29495
rect 22925 29455 22983 29461
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 25148 29501 25176 29532
rect 25133 29495 25191 29501
rect 25133 29461 25145 29495
rect 25179 29461 25191 29495
rect 25133 29455 25191 29461
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 7650 29248 7656 29300
rect 7708 29288 7714 29300
rect 7708 29260 12434 29288
rect 7708 29248 7714 29260
rect 9769 29223 9827 29229
rect 9769 29220 9781 29223
rect 9246 29192 9781 29220
rect 9769 29189 9781 29192
rect 9815 29220 9827 29223
rect 10226 29220 10232 29232
rect 9815 29192 10232 29220
rect 9815 29189 9827 29192
rect 9769 29183 9827 29189
rect 10226 29180 10232 29192
rect 10284 29180 10290 29232
rect 12406 29220 12434 29260
rect 12894 29248 12900 29300
rect 12952 29248 12958 29300
rect 13538 29248 13544 29300
rect 13596 29288 13602 29300
rect 13722 29288 13728 29300
rect 13596 29260 13728 29288
rect 13596 29248 13602 29260
rect 13722 29248 13728 29260
rect 13780 29248 13786 29300
rect 14182 29248 14188 29300
rect 14240 29248 14246 29300
rect 15289 29291 15347 29297
rect 15289 29257 15301 29291
rect 15335 29288 15347 29291
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15335 29260 16037 29288
rect 15335 29257 15347 29260
rect 15289 29251 15347 29257
rect 16025 29257 16037 29260
rect 16071 29288 16083 29291
rect 16114 29288 16120 29300
rect 16071 29260 16120 29288
rect 16071 29257 16083 29260
rect 16025 29251 16083 29257
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 17218 29248 17224 29300
rect 17276 29248 17282 29300
rect 17313 29291 17371 29297
rect 17313 29257 17325 29291
rect 17359 29288 17371 29291
rect 17494 29288 17500 29300
rect 17359 29260 17500 29288
rect 17359 29257 17371 29260
rect 17313 29251 17371 29257
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 17957 29291 18015 29297
rect 17957 29288 17969 29291
rect 17644 29260 17969 29288
rect 17644 29248 17650 29260
rect 17957 29257 17969 29260
rect 18003 29288 18015 29291
rect 18003 29260 19334 29288
rect 18003 29257 18015 29260
rect 17957 29251 18015 29257
rect 12406 29192 15516 29220
rect 12989 29155 13047 29161
rect 9508 29124 12756 29152
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 7745 29087 7803 29093
rect 7745 29084 7757 29087
rect 6604 29056 7757 29084
rect 6604 29044 6610 29056
rect 7745 29053 7757 29056
rect 7791 29053 7803 29087
rect 7745 29047 7803 29053
rect 9398 29044 9404 29096
rect 9456 29084 9462 29096
rect 9508 29093 9536 29124
rect 9493 29087 9551 29093
rect 9493 29084 9505 29087
rect 9456 29056 9505 29084
rect 9456 29044 9462 29056
rect 9493 29053 9505 29056
rect 9539 29053 9551 29087
rect 9493 29047 9551 29053
rect 10870 28976 10876 29028
rect 10928 29016 10934 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 10928 28988 12541 29016
rect 10928 28976 10934 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 12728 29016 12756 29124
rect 12989 29121 13001 29155
rect 13035 29152 13047 29155
rect 13035 29124 13400 29152
rect 13035 29121 13047 29124
rect 12989 29115 13047 29121
rect 13081 29087 13139 29093
rect 13081 29053 13093 29087
rect 13127 29053 13139 29087
rect 13081 29047 13139 29053
rect 13096 29016 13124 29047
rect 12728 28988 13124 29016
rect 12529 28979 12587 28985
rect 8008 28951 8066 28957
rect 8008 28917 8020 28951
rect 8054 28948 8066 28951
rect 8662 28948 8668 28960
rect 8054 28920 8668 28948
rect 8054 28917 8066 28920
rect 8008 28911 8066 28917
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 13372 28948 13400 29124
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 13780 29124 13860 29152
rect 13780 29112 13786 29124
rect 13446 28976 13452 29028
rect 13504 29016 13510 29028
rect 13725 29019 13783 29025
rect 13725 29016 13737 29019
rect 13504 28988 13737 29016
rect 13504 28976 13510 28988
rect 13725 28985 13737 28988
rect 13771 28985 13783 29019
rect 13832 29016 13860 29124
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 14274 29112 14280 29164
rect 14332 29152 14338 29164
rect 14332 29124 15056 29152
rect 14332 29112 14338 29124
rect 14369 29087 14427 29093
rect 14369 29053 14381 29087
rect 14415 29084 14427 29087
rect 14642 29084 14648 29096
rect 14415 29056 14648 29084
rect 14415 29053 14427 29056
rect 14369 29047 14427 29053
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 14921 29019 14979 29025
rect 14921 29016 14933 29019
rect 13832 28988 14933 29016
rect 13725 28979 13783 28985
rect 14921 28985 14933 28988
rect 14967 28985 14979 29019
rect 15028 29016 15056 29124
rect 15286 29044 15292 29096
rect 15344 29084 15350 29096
rect 15488 29093 15516 29192
rect 15562 29180 15568 29232
rect 15620 29220 15626 29232
rect 16209 29223 16267 29229
rect 16209 29220 16221 29223
rect 15620 29192 16221 29220
rect 15620 29180 15626 29192
rect 16132 29164 16160 29192
rect 16209 29189 16221 29192
rect 16255 29220 16267 29223
rect 18874 29220 18880 29232
rect 16255 29192 18880 29220
rect 16255 29189 16267 29192
rect 16209 29183 16267 29189
rect 18874 29180 18880 29192
rect 18932 29180 18938 29232
rect 19306 29220 19334 29260
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 22373 29291 22431 29297
rect 22373 29288 22385 29291
rect 20956 29260 22385 29288
rect 20956 29248 20962 29260
rect 22373 29257 22385 29260
rect 22419 29257 22431 29291
rect 22373 29251 22431 29257
rect 23934 29248 23940 29300
rect 23992 29248 23998 29300
rect 25314 29248 25320 29300
rect 25372 29248 25378 29300
rect 25498 29248 25504 29300
rect 25556 29248 25562 29300
rect 20070 29220 20076 29232
rect 19306 29192 20076 29220
rect 20070 29180 20076 29192
rect 20128 29220 20134 29232
rect 20128 29192 21220 29220
rect 20128 29180 20134 29192
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 16408 29124 19717 29152
rect 16408 29096 16436 29124
rect 19705 29121 19717 29124
rect 19751 29152 19763 29155
rect 20441 29155 20499 29161
rect 20441 29152 20453 29155
rect 19751 29124 20453 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 20441 29121 20453 29124
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29152 20591 29155
rect 20579 29124 21036 29152
rect 20579 29121 20591 29124
rect 20533 29115 20591 29121
rect 21008 29096 21036 29124
rect 15381 29087 15439 29093
rect 15381 29084 15393 29087
rect 15344 29056 15393 29084
rect 15344 29044 15350 29056
rect 15381 29053 15393 29056
rect 15427 29053 15439 29087
rect 15381 29047 15439 29053
rect 15473 29087 15531 29093
rect 15473 29053 15485 29087
rect 15519 29053 15531 29087
rect 15473 29047 15531 29053
rect 16390 29044 16396 29096
rect 16448 29044 16454 29096
rect 16666 29044 16672 29096
rect 16724 29084 16730 29096
rect 16724 29056 16988 29084
rect 16724 29044 16730 29056
rect 15028 28988 15976 29016
rect 14921 28979 14979 28985
rect 13998 28948 14004 28960
rect 13372 28920 14004 28948
rect 13998 28908 14004 28920
rect 14056 28908 14062 28960
rect 14182 28908 14188 28960
rect 14240 28948 14246 28960
rect 15746 28948 15752 28960
rect 14240 28920 15752 28948
rect 14240 28908 14246 28920
rect 15746 28908 15752 28920
rect 15804 28908 15810 28960
rect 15948 28948 15976 28988
rect 16022 28976 16028 29028
rect 16080 29016 16086 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 16080 28988 16865 29016
rect 16080 28976 16086 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 16960 29016 16988 29056
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 19518 29084 19524 29096
rect 17696 29056 19524 29084
rect 17586 29016 17592 29028
rect 16960 28988 17592 29016
rect 16853 28979 16911 28985
rect 17586 28976 17592 28988
rect 17644 28976 17650 29028
rect 17696 28948 17724 29056
rect 19518 29044 19524 29056
rect 19576 29044 19582 29096
rect 20625 29087 20683 29093
rect 20625 29084 20637 29087
rect 20456 29056 20637 29084
rect 20456 29028 20484 29056
rect 20625 29053 20637 29056
rect 20671 29053 20683 29087
rect 20625 29047 20683 29053
rect 20990 29044 20996 29096
rect 21048 29084 21054 29096
rect 21085 29087 21143 29093
rect 21085 29084 21097 29087
rect 21048 29056 21097 29084
rect 21048 29044 21054 29056
rect 21085 29053 21097 29056
rect 21131 29053 21143 29087
rect 21192 29084 21220 29192
rect 21542 29180 21548 29232
rect 21600 29220 21606 29232
rect 21600 29192 22094 29220
rect 21600 29180 21606 29192
rect 22066 29152 22094 29192
rect 24578 29180 24584 29232
rect 24636 29220 24642 29232
rect 24673 29223 24731 29229
rect 24673 29220 24685 29223
rect 24636 29192 24685 29220
rect 24636 29180 24642 29192
rect 24673 29189 24685 29192
rect 24719 29189 24731 29223
rect 24673 29183 24731 29189
rect 22465 29155 22523 29161
rect 22465 29152 22477 29155
rect 22066 29124 22477 29152
rect 22465 29121 22477 29124
rect 22511 29121 22523 29155
rect 23474 29152 23480 29164
rect 22465 29115 22523 29121
rect 22572 29124 23480 29152
rect 22572 29084 22600 29124
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 24118 29152 24124 29164
rect 23707 29124 24124 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 21192 29056 22600 29084
rect 22649 29087 22707 29093
rect 21085 29047 21143 29053
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23566 29084 23572 29096
rect 22695 29056 23572 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23566 29044 23572 29056
rect 23624 29044 23630 29096
rect 18046 28976 18052 29028
rect 18104 29016 18110 29028
rect 18322 29016 18328 29028
rect 18104 28988 18328 29016
rect 18104 28976 18110 28988
rect 18322 28976 18328 28988
rect 18380 28976 18386 29028
rect 20073 29019 20131 29025
rect 20073 28985 20085 29019
rect 20119 29016 20131 29019
rect 20119 28988 20392 29016
rect 20119 28985 20131 28988
rect 20073 28979 20131 28985
rect 15948 28920 17724 28948
rect 18414 28908 18420 28960
rect 18472 28948 18478 28960
rect 18874 28948 18880 28960
rect 18472 28920 18880 28948
rect 18472 28908 18478 28920
rect 18874 28908 18880 28920
rect 18932 28908 18938 28960
rect 20364 28948 20392 28988
rect 20438 28976 20444 29028
rect 20496 28976 20502 29028
rect 21634 29016 21640 29028
rect 20548 28988 21640 29016
rect 20548 28948 20576 28988
rect 21634 28976 21640 28988
rect 21692 28976 21698 29028
rect 22005 29019 22063 29025
rect 22005 28985 22017 29019
rect 22051 29016 22063 29019
rect 23290 29016 23296 29028
rect 22051 28988 23296 29016
rect 22051 28985 22063 28988
rect 22005 28979 22063 28985
rect 23290 28976 23296 28988
rect 23348 28976 23354 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 23440 28988 24869 29016
rect 23440 28976 23446 28988
rect 24857 28985 24869 28988
rect 24903 28985 24915 29019
rect 24857 28979 24915 28985
rect 20364 28920 20576 28948
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 12805 28747 12863 28753
rect 12805 28713 12817 28747
rect 12851 28744 12863 28747
rect 14090 28744 14096 28756
rect 12851 28716 14096 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 14090 28704 14096 28716
rect 14148 28704 14154 28756
rect 14826 28704 14832 28756
rect 14884 28704 14890 28756
rect 16758 28704 16764 28756
rect 16816 28744 16822 28756
rect 21266 28744 21272 28756
rect 16816 28716 21272 28744
rect 16816 28704 16822 28716
rect 21266 28704 21272 28716
rect 21324 28704 21330 28756
rect 14844 28676 14872 28704
rect 18414 28676 18420 28688
rect 14844 28648 18420 28676
rect 18414 28636 18420 28648
rect 18472 28636 18478 28688
rect 21174 28636 21180 28688
rect 21232 28636 21238 28688
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 2041 28611 2099 28617
rect 2041 28608 2053 28611
rect 1360 28580 2053 28608
rect 1360 28568 1366 28580
rect 2041 28577 2053 28580
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 4154 28568 4160 28620
rect 4212 28608 4218 28620
rect 4249 28611 4307 28617
rect 4249 28608 4261 28611
rect 4212 28580 4261 28608
rect 4212 28568 4218 28580
rect 4249 28577 4261 28580
rect 4295 28577 4307 28611
rect 4249 28571 4307 28577
rect 5626 28568 5632 28620
rect 5684 28568 5690 28620
rect 6546 28568 6552 28620
rect 6604 28568 6610 28620
rect 6825 28611 6883 28617
rect 6825 28577 6837 28611
rect 6871 28608 6883 28611
rect 8297 28611 8355 28617
rect 6871 28580 8248 28608
rect 6871 28577 6883 28580
rect 6825 28571 6883 28577
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 8110 28540 8116 28552
rect 7958 28512 8116 28540
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 8220 28540 8248 28580
rect 8297 28577 8309 28611
rect 8343 28608 8355 28611
rect 9858 28608 9864 28620
rect 8343 28580 9864 28608
rect 8343 28577 8355 28580
rect 8297 28571 8355 28577
rect 9858 28568 9864 28580
rect 9916 28568 9922 28620
rect 10873 28611 10931 28617
rect 10873 28577 10885 28611
rect 10919 28608 10931 28611
rect 11330 28608 11336 28620
rect 10919 28580 11336 28608
rect 10919 28577 10931 28580
rect 10873 28571 10931 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 12710 28608 12716 28620
rect 12406 28580 12716 28608
rect 9398 28540 9404 28552
rect 8220 28512 9404 28540
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10597 28543 10655 28549
rect 10597 28540 10609 28543
rect 10008 28512 10609 28540
rect 10008 28500 10014 28512
rect 10597 28509 10609 28512
rect 10643 28509 10655 28543
rect 12406 28540 12434 28580
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 13354 28568 13360 28620
rect 13412 28568 13418 28620
rect 14826 28568 14832 28620
rect 14884 28568 14890 28620
rect 16206 28568 16212 28620
rect 16264 28568 16270 28620
rect 17126 28568 17132 28620
rect 17184 28608 17190 28620
rect 17681 28611 17739 28617
rect 17681 28608 17693 28611
rect 17184 28580 17693 28608
rect 17184 28568 17190 28580
rect 17681 28577 17693 28580
rect 17727 28577 17739 28611
rect 17681 28571 17739 28577
rect 17770 28568 17776 28620
rect 17828 28568 17834 28620
rect 19429 28611 19487 28617
rect 19429 28577 19441 28611
rect 19475 28608 19487 28611
rect 22002 28608 22008 28620
rect 19475 28580 22008 28608
rect 19475 28577 19487 28580
rect 19429 28571 19487 28577
rect 22002 28568 22008 28580
rect 22060 28568 22066 28620
rect 22830 28568 22836 28620
rect 22888 28608 22894 28620
rect 22888 28580 24808 28608
rect 22888 28568 22894 28580
rect 12006 28512 12434 28540
rect 14645 28543 14703 28549
rect 10597 28503 10655 28509
rect 14645 28509 14657 28543
rect 14691 28540 14703 28543
rect 15562 28540 15568 28552
rect 14691 28512 15568 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15562 28500 15568 28512
rect 15620 28500 15626 28552
rect 16022 28500 16028 28552
rect 16080 28500 16086 28552
rect 16117 28543 16175 28549
rect 16117 28509 16129 28543
rect 16163 28540 16175 28543
rect 16850 28540 16856 28552
rect 16163 28512 16856 28540
rect 16163 28509 16175 28512
rect 16117 28503 16175 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 17589 28543 17647 28549
rect 17589 28509 17601 28543
rect 17635 28540 17647 28543
rect 19058 28540 19064 28552
rect 17635 28512 19064 28540
rect 17635 28509 17647 28512
rect 17589 28503 17647 28509
rect 19058 28500 19064 28512
rect 19116 28500 19122 28552
rect 24780 28549 24808 28580
rect 24029 28543 24087 28549
rect 24029 28509 24041 28543
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 24765 28543 24823 28549
rect 24765 28509 24777 28543
rect 24811 28509 24823 28543
rect 24765 28503 24823 28509
rect 3970 28432 3976 28484
rect 4028 28472 4034 28484
rect 4433 28475 4491 28481
rect 4433 28472 4445 28475
rect 4028 28444 4445 28472
rect 4028 28432 4034 28444
rect 4433 28441 4445 28444
rect 4479 28441 4491 28475
rect 18046 28472 18052 28484
rect 4433 28435 4491 28441
rect 8128 28444 11284 28472
rect 5534 28364 5540 28416
rect 5592 28404 5598 28416
rect 8128 28404 8156 28444
rect 5592 28376 8156 28404
rect 5592 28364 5598 28376
rect 8202 28364 8208 28416
rect 8260 28404 8266 28416
rect 8665 28407 8723 28413
rect 8665 28404 8677 28407
rect 8260 28376 8677 28404
rect 8260 28364 8266 28376
rect 8665 28373 8677 28376
rect 8711 28404 8723 28407
rect 10226 28404 10232 28416
rect 8711 28376 10232 28404
rect 8711 28373 8723 28376
rect 8665 28367 8723 28373
rect 10226 28364 10232 28376
rect 10284 28364 10290 28416
rect 11256 28404 11284 28444
rect 12176 28444 18052 28472
rect 12176 28404 12204 28444
rect 18046 28432 18052 28444
rect 18104 28432 18110 28484
rect 19705 28475 19763 28481
rect 19705 28441 19717 28475
rect 19751 28472 19763 28475
rect 19794 28472 19800 28484
rect 19751 28444 19800 28472
rect 19751 28441 19763 28444
rect 19705 28435 19763 28441
rect 19794 28432 19800 28444
rect 19852 28432 19858 28484
rect 21450 28472 21456 28484
rect 20930 28444 21456 28472
rect 21450 28432 21456 28444
rect 21508 28432 21514 28484
rect 24044 28472 24072 28503
rect 24210 28472 24216 28484
rect 24044 28444 24216 28472
rect 24210 28432 24216 28444
rect 24268 28472 24274 28484
rect 24854 28472 24860 28484
rect 24268 28444 24860 28472
rect 24268 28432 24274 28444
rect 24854 28432 24860 28444
rect 24912 28432 24918 28484
rect 11256 28376 12204 28404
rect 12345 28407 12403 28413
rect 12345 28373 12357 28407
rect 12391 28404 12403 28407
rect 12802 28404 12808 28416
rect 12391 28376 12808 28404
rect 12391 28373 12403 28376
rect 12345 28367 12403 28373
rect 12802 28364 12808 28376
rect 12860 28364 12866 28416
rect 13170 28364 13176 28416
rect 13228 28364 13234 28416
rect 13262 28364 13268 28416
rect 13320 28364 13326 28416
rect 13909 28407 13967 28413
rect 13909 28373 13921 28407
rect 13955 28404 13967 28407
rect 13998 28404 14004 28416
rect 13955 28376 14004 28404
rect 13955 28373 13967 28376
rect 13909 28367 13967 28373
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 14274 28364 14280 28416
rect 14332 28364 14338 28416
rect 14550 28364 14556 28416
rect 14608 28404 14614 28416
rect 14737 28407 14795 28413
rect 14737 28404 14749 28407
rect 14608 28376 14749 28404
rect 14608 28364 14614 28376
rect 14737 28373 14749 28376
rect 14783 28373 14795 28407
rect 14737 28367 14795 28373
rect 15286 28364 15292 28416
rect 15344 28364 15350 28416
rect 15657 28407 15715 28413
rect 15657 28373 15669 28407
rect 15703 28404 15715 28407
rect 15746 28404 15752 28416
rect 15703 28376 15752 28404
rect 15703 28373 15715 28376
rect 15657 28367 15715 28373
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16942 28364 16948 28416
rect 17000 28404 17006 28416
rect 17221 28407 17279 28413
rect 17221 28404 17233 28407
rect 17000 28376 17233 28404
rect 17000 28364 17006 28376
rect 17221 28373 17233 28376
rect 17267 28373 17279 28407
rect 17221 28367 17279 28373
rect 18414 28364 18420 28416
rect 18472 28404 18478 28416
rect 23845 28407 23903 28413
rect 23845 28404 23857 28407
rect 18472 28376 23857 28404
rect 18472 28364 18478 28376
rect 23845 28373 23857 28376
rect 23891 28373 23903 28407
rect 23845 28367 23903 28373
rect 24578 28364 24584 28416
rect 24636 28364 24642 28416
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 1946 28160 1952 28212
rect 2004 28200 2010 28212
rect 3786 28209 3792 28212
rect 2041 28203 2099 28209
rect 2041 28200 2053 28203
rect 2004 28172 2053 28200
rect 2004 28160 2010 28172
rect 2041 28169 2053 28172
rect 2087 28169 2099 28203
rect 2041 28163 2099 28169
rect 3743 28203 3792 28209
rect 3743 28169 3755 28203
rect 3789 28169 3792 28203
rect 3743 28163 3792 28169
rect 3786 28160 3792 28163
rect 3844 28160 3850 28212
rect 10226 28160 10232 28212
rect 10284 28200 10290 28212
rect 10321 28203 10379 28209
rect 10321 28200 10333 28203
rect 10284 28172 10333 28200
rect 10284 28160 10290 28172
rect 10321 28169 10333 28172
rect 10367 28169 10379 28203
rect 10321 28163 10379 28169
rect 12621 28203 12679 28209
rect 12621 28169 12633 28203
rect 12667 28200 12679 28203
rect 13170 28200 13176 28212
rect 12667 28172 13176 28200
rect 12667 28169 12679 28172
rect 12621 28163 12679 28169
rect 13170 28160 13176 28172
rect 13228 28160 13234 28212
rect 15838 28160 15844 28212
rect 15896 28200 15902 28212
rect 15933 28203 15991 28209
rect 15933 28200 15945 28203
rect 15896 28172 15945 28200
rect 15896 28160 15902 28172
rect 15933 28169 15945 28172
rect 15979 28200 15991 28203
rect 16853 28203 16911 28209
rect 16853 28200 16865 28203
rect 15979 28172 16865 28200
rect 15979 28169 15991 28172
rect 15933 28163 15991 28169
rect 16853 28169 16865 28172
rect 16899 28169 16911 28203
rect 16853 28163 16911 28169
rect 18322 28160 18328 28212
rect 18380 28160 18386 28212
rect 19521 28203 19579 28209
rect 19521 28169 19533 28203
rect 19567 28200 19579 28203
rect 20162 28200 20168 28212
rect 19567 28172 20168 28200
rect 19567 28169 19579 28172
rect 19521 28163 19579 28169
rect 20162 28160 20168 28172
rect 20220 28160 20226 28212
rect 22646 28160 22652 28212
rect 22704 28200 22710 28212
rect 24121 28203 24179 28209
rect 24121 28200 24133 28203
rect 22704 28172 24133 28200
rect 22704 28160 22710 28172
rect 24121 28169 24133 28172
rect 24167 28169 24179 28203
rect 24121 28163 24179 28169
rect 10244 28132 10272 28160
rect 16761 28135 16819 28141
rect 9798 28104 12434 28132
rect 2225 28067 2283 28073
rect 2225 28033 2237 28067
rect 2271 28064 2283 28067
rect 3418 28064 3424 28076
rect 2271 28036 3424 28064
rect 2271 28033 2283 28036
rect 2225 28027 2283 28033
rect 3418 28024 3424 28036
rect 3476 28024 3482 28076
rect 3602 28024 3608 28076
rect 3660 28073 3666 28076
rect 3660 28067 3698 28073
rect 3686 28033 3698 28067
rect 3660 28027 3698 28033
rect 3660 28024 3666 28027
rect 8297 27999 8355 28005
rect 8297 27965 8309 27999
rect 8343 27996 8355 27999
rect 8343 27968 8432 27996
rect 8343 27965 8355 27968
rect 8297 27959 8355 27965
rect 8404 27860 8432 27968
rect 8570 27956 8576 28008
rect 8628 27956 8634 28008
rect 8662 27956 8668 28008
rect 8720 27996 8726 28008
rect 8720 27968 10088 27996
rect 8720 27956 8726 27968
rect 10060 27937 10088 27968
rect 10045 27931 10103 27937
rect 10045 27897 10057 27931
rect 10091 27928 10103 27931
rect 11238 27928 11244 27940
rect 10091 27900 11244 27928
rect 10091 27897 10103 27900
rect 10045 27891 10103 27897
rect 11238 27888 11244 27900
rect 11296 27888 11302 27940
rect 9950 27860 9956 27872
rect 8404 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27820 10014 27872
rect 12406 27860 12434 28104
rect 16761 28101 16773 28135
rect 16807 28132 16819 28135
rect 18874 28132 18880 28144
rect 16807 28104 18880 28132
rect 16807 28101 16819 28104
rect 16761 28095 16819 28101
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28064 13231 28067
rect 13262 28064 13268 28076
rect 13219 28036 13268 28064
rect 13219 28033 13231 28036
rect 13173 28027 13231 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 16022 27956 16028 28008
rect 16080 27956 16086 28008
rect 16206 27956 16212 28008
rect 16264 27996 16270 28008
rect 16776 27996 16804 28095
rect 18874 28092 18880 28104
rect 18932 28092 18938 28144
rect 20806 28132 20812 28144
rect 18984 28104 20812 28132
rect 17494 28024 17500 28076
rect 17552 28064 17558 28076
rect 18233 28067 18291 28073
rect 18233 28064 18245 28067
rect 17552 28036 18245 28064
rect 17552 28024 17558 28036
rect 18233 28033 18245 28036
rect 18279 28033 18291 28067
rect 18984 28064 19012 28104
rect 20806 28092 20812 28104
rect 20864 28092 20870 28144
rect 21450 28092 21456 28144
rect 21508 28132 21514 28144
rect 22664 28132 22692 28160
rect 21508 28104 22770 28132
rect 21508 28092 21514 28104
rect 24670 28092 24676 28144
rect 24728 28092 24734 28144
rect 18233 28027 18291 28033
rect 18708 28036 19012 28064
rect 16264 27968 16804 27996
rect 18509 27999 18567 28005
rect 16264 27956 16270 27968
rect 18509 27965 18521 27999
rect 18555 27996 18567 27999
rect 18598 27996 18604 28008
rect 18555 27968 18604 27996
rect 18555 27965 18567 27968
rect 18509 27959 18567 27965
rect 18598 27956 18604 27968
rect 18656 27956 18662 28008
rect 16040 27928 16068 27956
rect 17037 27931 17095 27937
rect 17037 27928 17049 27931
rect 15396 27900 15700 27928
rect 16040 27900 17049 27928
rect 15396 27872 15424 27900
rect 12710 27860 12716 27872
rect 12406 27832 12716 27860
rect 12710 27820 12716 27832
rect 12768 27860 12774 27872
rect 13265 27863 13323 27869
rect 13265 27860 13277 27863
rect 12768 27832 13277 27860
rect 12768 27820 12774 27832
rect 13265 27829 13277 27832
rect 13311 27829 13323 27863
rect 13265 27823 13323 27829
rect 14550 27820 14556 27872
rect 14608 27860 14614 27872
rect 15105 27863 15163 27869
rect 15105 27860 15117 27863
rect 14608 27832 15117 27860
rect 14608 27820 14614 27832
rect 15105 27829 15117 27832
rect 15151 27860 15163 27863
rect 15378 27860 15384 27872
rect 15151 27832 15384 27860
rect 15151 27829 15163 27832
rect 15105 27823 15163 27829
rect 15378 27820 15384 27832
rect 15436 27820 15442 27872
rect 15562 27820 15568 27872
rect 15620 27820 15626 27872
rect 15672 27860 15700 27900
rect 17037 27897 17049 27900
rect 17083 27928 17095 27931
rect 18708 27928 18736 28036
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19429 28067 19487 28073
rect 19429 28064 19441 28067
rect 19392 28036 19441 28064
rect 19392 28024 19398 28036
rect 19429 28033 19441 28036
rect 19475 28033 19487 28067
rect 19429 28027 19487 28033
rect 22002 28024 22008 28076
rect 22060 28024 22066 28076
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27996 19763 27999
rect 19978 27996 19984 28008
rect 19751 27968 19984 27996
rect 19751 27965 19763 27968
rect 19705 27959 19763 27965
rect 19978 27956 19984 27968
rect 20036 27956 20042 28008
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 24670 27996 24676 28008
rect 22327 27968 24676 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 17083 27900 18736 27928
rect 17083 27897 17095 27900
rect 17037 27891 17095 27897
rect 18782 27888 18788 27940
rect 18840 27928 18846 27940
rect 24857 27931 24915 27937
rect 18840 27900 22094 27928
rect 18840 27888 18846 27900
rect 17494 27860 17500 27872
rect 15672 27832 17500 27860
rect 17494 27820 17500 27832
rect 17552 27820 17558 27872
rect 17865 27863 17923 27869
rect 17865 27829 17877 27863
rect 17911 27860 17923 27863
rect 18966 27860 18972 27872
rect 17911 27832 18972 27860
rect 17911 27829 17923 27832
rect 17865 27823 17923 27829
rect 18966 27820 18972 27832
rect 19024 27820 19030 27872
rect 19058 27820 19064 27872
rect 19116 27820 19122 27872
rect 22066 27860 22094 27900
rect 24857 27897 24869 27931
rect 24903 27928 24915 27931
rect 25130 27928 25136 27940
rect 24903 27900 25136 27928
rect 24903 27897 24915 27900
rect 24857 27891 24915 27897
rect 25130 27888 25136 27900
rect 25188 27888 25194 27940
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 22066 27832 23765 27860
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 6444 27659 6502 27665
rect 6444 27625 6456 27659
rect 6490 27656 6502 27659
rect 9858 27656 9864 27668
rect 6490 27628 9864 27656
rect 6490 27625 6502 27628
rect 6444 27619 6502 27625
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 18322 27616 18328 27668
rect 18380 27656 18386 27668
rect 18693 27659 18751 27665
rect 18693 27656 18705 27659
rect 18380 27628 18705 27656
rect 18380 27616 18386 27628
rect 18693 27625 18705 27628
rect 18739 27625 18751 27659
rect 18693 27619 18751 27625
rect 18782 27616 18788 27668
rect 18840 27656 18846 27668
rect 19334 27656 19340 27668
rect 18840 27628 19340 27656
rect 18840 27616 18846 27628
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 24210 27616 24216 27668
rect 24268 27616 24274 27668
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 7929 27591 7987 27597
rect 7929 27588 7941 27591
rect 7892 27560 7941 27588
rect 7892 27548 7898 27560
rect 7929 27557 7941 27560
rect 7975 27557 7987 27591
rect 7929 27551 7987 27557
rect 8294 27548 8300 27600
rect 8352 27588 8358 27600
rect 8389 27591 8447 27597
rect 8389 27588 8401 27591
rect 8352 27560 8401 27588
rect 8352 27548 8358 27560
rect 8389 27557 8401 27560
rect 8435 27557 8447 27591
rect 8389 27551 8447 27557
rect 20073 27591 20131 27597
rect 20073 27557 20085 27591
rect 20119 27588 20131 27591
rect 21082 27588 21088 27600
rect 20119 27560 21088 27588
rect 20119 27557 20131 27560
rect 20073 27551 20131 27557
rect 21082 27548 21088 27560
rect 21140 27548 21146 27600
rect 6181 27523 6239 27529
rect 6181 27489 6193 27523
rect 6227 27520 6239 27523
rect 6546 27520 6552 27532
rect 6227 27492 6552 27520
rect 6227 27489 6239 27492
rect 6181 27483 6239 27489
rect 6546 27480 6552 27492
rect 6604 27480 6610 27532
rect 7558 27412 7564 27464
rect 7616 27452 7622 27464
rect 8312 27452 8340 27548
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 12860 27492 15669 27520
rect 12860 27480 12866 27492
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 17126 27480 17132 27532
rect 17184 27520 17190 27532
rect 17184 27492 18736 27520
rect 17184 27480 17190 27492
rect 7616 27424 8340 27452
rect 7616 27412 7622 27424
rect 9950 27412 9956 27464
rect 10008 27452 10014 27464
rect 10962 27452 10968 27464
rect 10008 27424 10968 27452
rect 10008 27412 10014 27424
rect 10962 27412 10968 27424
rect 11020 27452 11026 27464
rect 11149 27455 11207 27461
rect 11149 27452 11161 27455
rect 11020 27424 11161 27452
rect 11020 27412 11026 27424
rect 11149 27421 11161 27424
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 15470 27412 15476 27464
rect 15528 27452 15534 27464
rect 15565 27455 15623 27461
rect 15565 27452 15577 27455
rect 15528 27424 15577 27452
rect 15528 27412 15534 27424
rect 15565 27421 15577 27424
rect 15611 27452 15623 27455
rect 16117 27455 16175 27461
rect 16117 27452 16129 27455
rect 15611 27424 16129 27452
rect 15611 27421 15623 27424
rect 15565 27415 15623 27421
rect 16117 27421 16129 27424
rect 16163 27421 16175 27455
rect 16117 27415 16175 27421
rect 11422 27344 11428 27396
rect 11480 27344 11486 27396
rect 12710 27384 12716 27396
rect 12650 27356 12716 27384
rect 12710 27344 12716 27356
rect 12768 27384 12774 27396
rect 16132 27384 16160 27415
rect 17034 27412 17040 27464
rect 17092 27452 17098 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 17092 27424 18337 27452
rect 17092 27412 17098 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18708 27448 18736 27492
rect 20530 27480 20536 27532
rect 20588 27480 20594 27532
rect 20622 27480 20628 27532
rect 20680 27480 20686 27532
rect 21910 27480 21916 27532
rect 21968 27480 21974 27532
rect 22738 27480 22744 27532
rect 22796 27520 22802 27532
rect 22796 27492 24716 27520
rect 22796 27480 22802 27492
rect 24688 27461 24716 27492
rect 24673 27455 24731 27461
rect 18708 27428 19012 27448
rect 18708 27420 19104 27428
rect 18984 27400 19104 27420
rect 24673 27421 24685 27455
rect 24719 27421 24731 27455
rect 24673 27415 24731 27421
rect 18230 27384 18236 27396
rect 12768 27356 13032 27384
rect 16132 27356 18236 27384
rect 12768 27344 12774 27356
rect 13004 27328 13032 27356
rect 18230 27344 18236 27356
rect 18288 27384 18294 27396
rect 18288 27356 18736 27384
rect 18288 27344 18294 27356
rect 10226 27276 10232 27328
rect 10284 27316 10290 27328
rect 12894 27316 12900 27328
rect 10284 27288 12900 27316
rect 10284 27276 10290 27288
rect 12894 27276 12900 27288
rect 12952 27276 12958 27328
rect 12986 27276 12992 27328
rect 13044 27316 13050 27328
rect 13265 27319 13323 27325
rect 13265 27316 13277 27319
rect 13044 27288 13277 27316
rect 13044 27276 13050 27288
rect 13265 27285 13277 27288
rect 13311 27316 13323 27319
rect 14090 27316 14096 27328
rect 13311 27288 14096 27316
rect 13311 27285 13323 27288
rect 13265 27279 13323 27285
rect 14090 27276 14096 27288
rect 14148 27276 14154 27328
rect 15010 27276 15016 27328
rect 15068 27316 15074 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 15068 27288 15117 27316
rect 15068 27276 15074 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 15105 27279 15163 27285
rect 15473 27319 15531 27325
rect 15473 27285 15485 27319
rect 15519 27316 15531 27319
rect 16390 27316 16396 27328
rect 15519 27288 16396 27316
rect 15519 27285 15531 27288
rect 15473 27279 15531 27285
rect 16390 27276 16396 27288
rect 16448 27276 16454 27328
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18598 27316 18604 27328
rect 18187 27288 18604 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18598 27276 18604 27288
rect 18656 27276 18662 27328
rect 18708 27316 18736 27356
rect 18969 27319 19027 27325
rect 18969 27316 18981 27319
rect 18708 27288 18981 27316
rect 18969 27285 18981 27288
rect 19015 27285 19027 27319
rect 19076 27316 19104 27400
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 22278 27344 22284 27396
rect 22336 27384 22342 27396
rect 22646 27384 22652 27396
rect 22336 27356 22652 27384
rect 22336 27344 22342 27356
rect 19797 27319 19855 27325
rect 19797 27316 19809 27319
rect 19076 27288 19809 27316
rect 18969 27279 19027 27285
rect 19797 27285 19809 27288
rect 19843 27316 19855 27319
rect 20441 27319 20499 27325
rect 20441 27316 20453 27319
rect 19843 27288 20453 27316
rect 19843 27285 19855 27288
rect 19797 27279 19855 27285
rect 20441 27285 20453 27288
rect 20487 27285 20499 27319
rect 22572 27316 22600 27356
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 24857 27387 24915 27393
rect 24857 27353 24869 27387
rect 24903 27384 24915 27387
rect 25038 27384 25044 27396
rect 24903 27356 25044 27384
rect 24903 27353 24915 27356
rect 24857 27347 24915 27353
rect 25038 27344 25044 27356
rect 25096 27344 25102 27396
rect 23014 27316 23020 27328
rect 22572 27288 23020 27316
rect 20441 27279 20499 27285
rect 23014 27276 23020 27288
rect 23072 27276 23078 27328
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 23661 27319 23719 27325
rect 23661 27316 23673 27319
rect 23164 27288 23673 27316
rect 23164 27276 23170 27288
rect 23661 27285 23673 27288
rect 23707 27285 23719 27319
rect 23661 27279 23719 27285
rect 25222 27276 25228 27328
rect 25280 27276 25286 27328
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 3191 27115 3249 27121
rect 3191 27081 3203 27115
rect 3237 27112 3249 27115
rect 3878 27112 3884 27124
rect 3237 27084 3884 27112
rect 3237 27081 3249 27084
rect 3191 27075 3249 27081
rect 3878 27072 3884 27084
rect 3936 27072 3942 27124
rect 6472 27084 10640 27112
rect 3120 26979 3178 26985
rect 3120 26945 3132 26979
rect 3166 26976 3178 26979
rect 3326 26976 3332 26988
rect 3166 26948 3332 26976
rect 3166 26945 3178 26948
rect 3120 26939 3178 26945
rect 3326 26936 3332 26948
rect 3384 26936 3390 26988
rect 3510 26936 3516 26988
rect 3568 26976 3574 26988
rect 3697 26979 3755 26985
rect 3697 26976 3709 26979
rect 3568 26948 3709 26976
rect 3568 26936 3574 26948
rect 3697 26945 3709 26948
rect 3743 26945 3755 26979
rect 3697 26939 3755 26945
rect 3881 26911 3939 26917
rect 3881 26877 3893 26911
rect 3927 26908 3939 26911
rect 4338 26908 4344 26920
rect 3927 26880 4344 26908
rect 3927 26877 3939 26880
rect 3881 26871 3939 26877
rect 4338 26868 4344 26880
rect 4396 26868 4402 26920
rect 4433 26911 4491 26917
rect 4433 26877 4445 26911
rect 4479 26908 4491 26911
rect 6472 26908 6500 27084
rect 7558 27004 7564 27056
rect 7616 27004 7622 27056
rect 10042 27004 10048 27056
rect 10100 27044 10106 27056
rect 10505 27047 10563 27053
rect 10505 27044 10517 27047
rect 10100 27016 10517 27044
rect 10100 27004 10106 27016
rect 10505 27013 10517 27016
rect 10551 27013 10563 27047
rect 10612 27044 10640 27084
rect 11514 27072 11520 27124
rect 11572 27112 11578 27124
rect 15105 27115 15163 27121
rect 15105 27112 15117 27115
rect 11572 27084 15117 27112
rect 11572 27072 11578 27084
rect 15105 27081 15117 27084
rect 15151 27081 15163 27115
rect 15105 27075 15163 27081
rect 15197 27115 15255 27121
rect 15197 27081 15209 27115
rect 15243 27112 15255 27115
rect 16574 27112 16580 27124
rect 15243 27084 16580 27112
rect 15243 27081 15255 27084
rect 15197 27075 15255 27081
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 17589 27115 17647 27121
rect 17589 27081 17601 27115
rect 17635 27112 17647 27115
rect 19981 27115 20039 27121
rect 19981 27112 19993 27115
rect 17635 27084 19993 27112
rect 17635 27081 17647 27084
rect 17589 27075 17647 27081
rect 19981 27081 19993 27084
rect 20027 27081 20039 27115
rect 19981 27075 20039 27081
rect 22554 27072 22560 27124
rect 22612 27112 22618 27124
rect 22738 27112 22744 27124
rect 22612 27084 22744 27112
rect 22612 27072 22618 27084
rect 22738 27072 22744 27084
rect 22796 27072 22802 27124
rect 24578 27112 24584 27124
rect 22848 27084 24584 27112
rect 13078 27044 13084 27056
rect 10612 27016 13084 27044
rect 10505 27007 10563 27013
rect 13078 27004 13084 27016
rect 13136 27004 13142 27056
rect 14090 27044 14096 27056
rect 14030 27016 14096 27044
rect 14090 27004 14096 27016
rect 14148 27004 14154 27056
rect 16390 27004 16396 27056
rect 16448 27044 16454 27056
rect 16448 27016 18092 27044
rect 16448 27004 16454 27016
rect 6546 26936 6552 26988
rect 6604 26936 6610 26988
rect 9122 26936 9128 26988
rect 9180 26936 9186 26988
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 12529 26979 12587 26985
rect 12529 26976 12541 26979
rect 11020 26948 12541 26976
rect 11020 26936 11026 26948
rect 12529 26945 12541 26948
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 18064 26976 18092 27016
rect 18138 27004 18144 27056
rect 18196 27044 18202 27056
rect 18414 27044 18420 27056
rect 18196 27016 18420 27044
rect 18196 27004 18202 27016
rect 18414 27004 18420 27016
rect 18472 27004 18478 27056
rect 21358 27044 21364 27056
rect 18524 27016 21364 27044
rect 18524 26976 18552 27016
rect 21358 27004 21364 27016
rect 21416 27004 21422 27056
rect 18064 26948 18552 26976
rect 19889 26979 19947 26985
rect 17957 26939 18015 26945
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 19935 26948 20729 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 22848 26976 22876 27084
rect 24578 27072 24584 27084
rect 24636 27072 24642 27124
rect 23014 27004 23020 27056
rect 23072 27044 23078 27056
rect 23566 27044 23572 27056
rect 23072 27016 23572 27044
rect 23072 27004 23078 27016
rect 23566 27004 23572 27016
rect 23624 27004 23630 27056
rect 24946 27004 24952 27056
rect 25004 27044 25010 27056
rect 25133 27047 25191 27053
rect 25133 27044 25145 27047
rect 25004 27016 25145 27044
rect 25004 27004 25010 27016
rect 25133 27013 25145 27016
rect 25179 27013 25191 27047
rect 25133 27007 25191 27013
rect 22419 26948 22876 26976
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 4479 26880 6500 26908
rect 6825 26911 6883 26917
rect 4479 26877 4491 26880
rect 4433 26871 4491 26877
rect 6825 26877 6837 26911
rect 6871 26908 6883 26911
rect 7834 26908 7840 26920
rect 6871 26880 7840 26908
rect 6871 26877 6883 26880
rect 6825 26871 6883 26877
rect 3694 26800 3700 26852
rect 3752 26840 3758 26852
rect 4448 26840 4476 26871
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 9217 26911 9275 26917
rect 9217 26908 9229 26911
rect 8720 26880 9229 26908
rect 8720 26868 8726 26880
rect 9217 26877 9229 26880
rect 9263 26877 9275 26911
rect 9217 26871 9275 26877
rect 9398 26868 9404 26920
rect 9456 26868 9462 26920
rect 12802 26868 12808 26920
rect 12860 26868 12866 26920
rect 12894 26868 12900 26920
rect 12952 26908 12958 26920
rect 15289 26911 15347 26917
rect 12952 26880 13860 26908
rect 12952 26868 12958 26880
rect 3752 26812 4476 26840
rect 3752 26800 3758 26812
rect 8294 26800 8300 26852
rect 8352 26840 8358 26852
rect 9674 26840 9680 26852
rect 8352 26812 9680 26840
rect 8352 26800 8358 26812
rect 9674 26800 9680 26812
rect 9732 26800 9738 26852
rect 10318 26800 10324 26852
rect 10376 26840 10382 26852
rect 10689 26843 10747 26849
rect 10689 26840 10701 26843
rect 10376 26812 10701 26840
rect 10376 26800 10382 26812
rect 10689 26809 10701 26812
rect 10735 26809 10747 26843
rect 13832 26840 13860 26880
rect 15289 26877 15301 26911
rect 15335 26877 15347 26911
rect 15289 26871 15347 26877
rect 15304 26840 15332 26871
rect 17402 26840 17408 26852
rect 13832 26812 15332 26840
rect 17144 26812 17408 26840
rect 10689 26803 10747 26809
rect 8757 26775 8815 26781
rect 8757 26741 8769 26775
rect 8803 26772 8815 26775
rect 10502 26772 10508 26784
rect 8803 26744 10508 26772
rect 8803 26741 8815 26744
rect 8757 26735 8815 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 11885 26775 11943 26781
rect 11885 26741 11897 26775
rect 11931 26772 11943 26775
rect 12986 26772 12992 26784
rect 11931 26744 12992 26772
rect 11931 26741 11943 26744
rect 11885 26735 11943 26741
rect 12986 26732 12992 26744
rect 13044 26732 13050 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14366 26772 14372 26784
rect 14323 26744 14372 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14366 26732 14372 26744
rect 14424 26732 14430 26784
rect 14737 26775 14795 26781
rect 14737 26741 14749 26775
rect 14783 26772 14795 26775
rect 17144 26772 17172 26812
rect 17402 26800 17408 26812
rect 17460 26800 17466 26852
rect 14783 26744 17172 26772
rect 17313 26775 17371 26781
rect 14783 26741 14795 26744
rect 14737 26735 14795 26741
rect 17313 26741 17325 26775
rect 17359 26772 17371 26775
rect 17972 26772 18000 26939
rect 18049 26911 18107 26917
rect 18049 26877 18061 26911
rect 18095 26908 18107 26911
rect 18138 26908 18144 26920
rect 18095 26880 18144 26908
rect 18095 26877 18107 26880
rect 18049 26871 18107 26877
rect 18138 26868 18144 26880
rect 18196 26868 18202 26920
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 19334 26908 19340 26920
rect 18279 26880 19340 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 19334 26868 19340 26880
rect 19392 26908 19398 26920
rect 19794 26908 19800 26920
rect 19392 26880 19800 26908
rect 19392 26868 19398 26880
rect 19794 26868 19800 26880
rect 19852 26868 19858 26920
rect 20165 26911 20223 26917
rect 20165 26877 20177 26911
rect 20211 26908 20223 26911
rect 21174 26908 21180 26920
rect 20211 26880 21180 26908
rect 20211 26877 20223 26880
rect 20165 26871 20223 26877
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 21450 26868 21456 26920
rect 21508 26908 21514 26920
rect 22002 26908 22008 26920
rect 21508 26880 22008 26908
rect 21508 26868 21514 26880
rect 22002 26868 22008 26880
rect 22060 26908 22066 26920
rect 22833 26911 22891 26917
rect 22833 26908 22845 26911
rect 22060 26880 22845 26908
rect 22060 26868 22066 26880
rect 22833 26877 22845 26880
rect 22879 26877 22891 26911
rect 23109 26911 23167 26917
rect 23109 26908 23121 26911
rect 22833 26871 22891 26877
rect 22940 26880 23121 26908
rect 20622 26800 20628 26852
rect 20680 26840 20686 26852
rect 22554 26840 22560 26852
rect 20680 26812 22560 26840
rect 20680 26800 20686 26812
rect 22554 26800 22560 26812
rect 22612 26840 22618 26852
rect 22940 26840 22968 26880
rect 23109 26877 23121 26880
rect 23155 26877 23167 26911
rect 23109 26871 23167 26877
rect 23198 26868 23204 26920
rect 23256 26908 23262 26920
rect 25317 26911 25375 26917
rect 25317 26908 25329 26911
rect 23256 26880 25329 26908
rect 23256 26868 23262 26880
rect 25317 26877 25329 26880
rect 25363 26877 25375 26911
rect 25317 26871 25375 26877
rect 22612 26812 22968 26840
rect 22612 26800 22618 26812
rect 18322 26772 18328 26784
rect 17359 26744 18328 26772
rect 17359 26741 17371 26744
rect 17313 26735 17371 26741
rect 18322 26732 18328 26744
rect 18380 26732 18386 26784
rect 19518 26732 19524 26784
rect 19576 26732 19582 26784
rect 22189 26775 22247 26781
rect 22189 26741 22201 26775
rect 22235 26772 22247 26775
rect 23842 26772 23848 26784
rect 22235 26744 23848 26772
rect 22235 26741 22247 26744
rect 22189 26735 22247 26741
rect 23842 26732 23848 26744
rect 23900 26732 23906 26784
rect 24578 26732 24584 26784
rect 24636 26732 24642 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 4062 26528 4068 26580
rect 4120 26528 4126 26580
rect 8570 26528 8576 26580
rect 8628 26568 8634 26580
rect 11701 26571 11759 26577
rect 11701 26568 11713 26571
rect 8628 26540 11713 26568
rect 8628 26528 8634 26540
rect 11701 26537 11713 26540
rect 11747 26537 11759 26571
rect 11701 26531 11759 26537
rect 11716 26500 11744 26531
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17129 26571 17187 26577
rect 17129 26568 17141 26571
rect 16724 26540 17141 26568
rect 16724 26528 16730 26540
rect 17129 26537 17141 26540
rect 17175 26568 17187 26571
rect 17770 26568 17776 26580
rect 17175 26540 17776 26568
rect 17175 26537 17187 26540
rect 17129 26531 17187 26537
rect 17770 26528 17776 26540
rect 17828 26528 17834 26580
rect 22186 26528 22192 26580
rect 22244 26568 22250 26580
rect 22373 26571 22431 26577
rect 22373 26568 22385 26571
rect 22244 26540 22385 26568
rect 22244 26528 22250 26540
rect 22373 26537 22385 26540
rect 22419 26537 22431 26571
rect 22373 26531 22431 26537
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 24578 26568 24584 26580
rect 22704 26540 24584 26568
rect 22704 26528 22710 26540
rect 24578 26528 24584 26540
rect 24636 26528 24642 26580
rect 14826 26500 14832 26512
rect 11716 26472 14832 26500
rect 14826 26460 14832 26472
rect 14884 26460 14890 26512
rect 17494 26460 17500 26512
rect 17552 26500 17558 26512
rect 17862 26500 17868 26512
rect 17552 26472 17868 26500
rect 17552 26460 17558 26472
rect 17862 26460 17868 26472
rect 17920 26460 17926 26512
rect 19429 26503 19487 26509
rect 19429 26469 19441 26503
rect 19475 26500 19487 26503
rect 19702 26500 19708 26512
rect 19475 26472 19708 26500
rect 19475 26469 19487 26472
rect 19429 26463 19487 26469
rect 19702 26460 19708 26472
rect 19760 26460 19766 26512
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22833 26503 22891 26509
rect 22833 26500 22845 26503
rect 22612 26472 22845 26500
rect 22612 26460 22618 26472
rect 22833 26469 22845 26472
rect 22879 26469 22891 26503
rect 22833 26463 22891 26469
rect 23566 26460 23572 26512
rect 23624 26500 23630 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23624 26472 23857 26500
rect 23624 26460 23630 26472
rect 23845 26469 23857 26472
rect 23891 26500 23903 26503
rect 25133 26503 25191 26509
rect 25133 26500 25145 26503
rect 23891 26472 25145 26500
rect 23891 26469 23903 26472
rect 23845 26463 23903 26469
rect 25133 26469 25145 26472
rect 25179 26500 25191 26503
rect 25222 26500 25228 26512
rect 25179 26472 25228 26500
rect 25179 26469 25191 26472
rect 25133 26463 25191 26469
rect 25222 26460 25228 26472
rect 25280 26460 25286 26512
rect 6454 26392 6460 26444
rect 6512 26392 6518 26444
rect 6733 26435 6791 26441
rect 6733 26401 6745 26435
rect 6779 26432 6791 26435
rect 8294 26432 8300 26444
rect 6779 26404 8300 26432
rect 6779 26401 6791 26404
rect 6733 26395 6791 26401
rect 8294 26392 8300 26404
rect 8352 26392 8358 26444
rect 9122 26392 9128 26444
rect 9180 26392 9186 26444
rect 10226 26392 10232 26444
rect 10284 26392 10290 26444
rect 11238 26392 11244 26444
rect 11296 26432 11302 26444
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11296 26404 12725 26432
rect 11296 26392 11302 26404
rect 12713 26401 12725 26404
rect 12759 26401 12771 26435
rect 12713 26395 12771 26401
rect 13538 26392 13544 26444
rect 13596 26432 13602 26444
rect 13906 26432 13912 26444
rect 13596 26404 13912 26432
rect 13596 26392 13602 26404
rect 13906 26392 13912 26404
rect 13964 26392 13970 26444
rect 15657 26435 15715 26441
rect 15657 26401 15669 26435
rect 15703 26432 15715 26435
rect 17512 26432 17540 26460
rect 15703 26404 17540 26432
rect 15703 26401 15715 26404
rect 15657 26395 15715 26401
rect 18966 26392 18972 26444
rect 19024 26432 19030 26444
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 19024 26404 19901 26432
rect 19024 26392 19030 26404
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 20162 26432 20168 26444
rect 20119 26404 20168 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 21450 26432 21456 26444
rect 20680 26404 21456 26432
rect 20680 26392 20686 26404
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 21634 26392 21640 26444
rect 21692 26432 21698 26444
rect 23293 26435 23351 26441
rect 23293 26432 23305 26435
rect 21692 26404 23305 26432
rect 21692 26392 21698 26404
rect 23293 26401 23305 26404
rect 23339 26401 23351 26435
rect 23293 26395 23351 26401
rect 23385 26435 23443 26441
rect 23385 26401 23397 26435
rect 23431 26432 23443 26435
rect 24578 26432 24584 26444
rect 23431 26404 24584 26432
rect 23431 26401 23443 26404
rect 23385 26395 23443 26401
rect 24578 26392 24584 26404
rect 24636 26392 24642 26444
rect 1765 26367 1823 26373
rect 1765 26333 1777 26367
rect 1811 26364 1823 26367
rect 2038 26364 2044 26376
rect 1811 26336 2044 26364
rect 1811 26333 1823 26336
rect 1765 26327 1823 26333
rect 2038 26324 2044 26336
rect 2096 26324 2102 26376
rect 9950 26324 9956 26376
rect 10008 26324 10014 26376
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26364 12679 26367
rect 14274 26364 14280 26376
rect 12667 26336 14280 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 14274 26324 14280 26336
rect 14332 26324 14338 26376
rect 15378 26324 15384 26376
rect 15436 26324 15442 26376
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20254 26364 20260 26376
rect 19843 26336 20260 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20254 26324 20260 26336
rect 20312 26324 20318 26376
rect 22278 26364 22284 26376
rect 22034 26336 22284 26364
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 24210 26324 24216 26376
rect 24268 26364 24274 26376
rect 24857 26367 24915 26373
rect 24857 26364 24869 26367
rect 24268 26336 24869 26364
rect 24268 26324 24274 26336
rect 24857 26333 24869 26336
rect 24903 26333 24915 26367
rect 24857 26327 24915 26333
rect 2774 26256 2780 26308
rect 2832 26256 2838 26308
rect 7466 26256 7472 26308
rect 7524 26256 7530 26308
rect 8662 26256 8668 26308
rect 8720 26256 8726 26308
rect 8754 26256 8760 26308
rect 8812 26296 8818 26308
rect 8812 26268 10718 26296
rect 8812 26256 8818 26268
rect 13354 26256 13360 26308
rect 13412 26296 13418 26308
rect 13538 26296 13544 26308
rect 13412 26268 13544 26296
rect 13412 26256 13418 26268
rect 13538 26256 13544 26268
rect 13596 26256 13602 26308
rect 15194 26256 15200 26308
rect 15252 26256 15258 26308
rect 17681 26299 17739 26305
rect 17681 26296 17693 26299
rect 16882 26268 17693 26296
rect 7650 26188 7656 26240
rect 7708 26228 7714 26240
rect 8205 26231 8263 26237
rect 8205 26228 8217 26231
rect 7708 26200 8217 26228
rect 7708 26188 7714 26200
rect 8205 26197 8217 26200
rect 8251 26197 8263 26231
rect 8205 26191 8263 26197
rect 12158 26188 12164 26240
rect 12216 26188 12222 26240
rect 12526 26188 12532 26240
rect 12584 26188 12590 26240
rect 14090 26188 14096 26240
rect 14148 26228 14154 26240
rect 14461 26231 14519 26237
rect 14461 26228 14473 26231
rect 14148 26200 14473 26228
rect 14148 26188 14154 26200
rect 14461 26197 14473 26200
rect 14507 26228 14519 26231
rect 14826 26228 14832 26240
rect 14507 26200 14832 26228
rect 14507 26197 14519 26200
rect 14461 26191 14519 26197
rect 14826 26188 14832 26200
rect 14884 26228 14890 26240
rect 15212 26228 15240 26256
rect 16960 26228 16988 26268
rect 17681 26265 17693 26268
rect 17727 26296 17739 26299
rect 17770 26296 17776 26308
rect 17727 26268 17776 26296
rect 17727 26265 17739 26268
rect 17681 26259 17739 26265
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 20901 26299 20959 26305
rect 20901 26265 20913 26299
rect 20947 26296 20959 26299
rect 21174 26296 21180 26308
rect 20947 26268 21180 26296
rect 20947 26265 20959 26268
rect 20901 26259 20959 26265
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 23201 26299 23259 26305
rect 23201 26296 23213 26299
rect 22204 26268 23213 26296
rect 14884 26200 16988 26228
rect 14884 26188 14890 26200
rect 21818 26188 21824 26240
rect 21876 26228 21882 26240
rect 22204 26228 22232 26268
rect 23201 26265 23213 26268
rect 23247 26265 23259 26299
rect 23201 26259 23259 26265
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 24673 26299 24731 26305
rect 24673 26296 24685 26299
rect 24544 26268 24685 26296
rect 24544 26256 24550 26268
rect 24673 26265 24685 26268
rect 24719 26265 24731 26299
rect 24673 26259 24731 26265
rect 21876 26200 22232 26228
rect 21876 26188 21882 26200
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 1762 25984 1768 26036
rect 1820 26024 1826 26036
rect 2133 26027 2191 26033
rect 2133 26024 2145 26027
rect 1820 25996 2145 26024
rect 1820 25984 1826 25996
rect 2133 25993 2145 25996
rect 2179 25993 2191 26027
rect 2133 25987 2191 25993
rect 7558 25984 7564 26036
rect 7616 26024 7622 26036
rect 8573 26027 8631 26033
rect 8573 26024 8585 26027
rect 7616 25996 8585 26024
rect 7616 25984 7622 25996
rect 8573 25993 8585 25996
rect 8619 26024 8631 26027
rect 8754 26024 8760 26036
rect 8619 25996 8760 26024
rect 8619 25993 8631 25996
rect 8573 25987 8631 25993
rect 8754 25984 8760 25996
rect 8812 25984 8818 26036
rect 9217 26027 9275 26033
rect 9217 25993 9229 26027
rect 9263 25993 9275 26027
rect 9217 25987 9275 25993
rect 3510 25916 3516 25968
rect 3568 25956 3574 25968
rect 4062 25956 4068 25968
rect 3568 25928 4068 25956
rect 3568 25916 3574 25928
rect 4062 25916 4068 25928
rect 4120 25956 4126 25968
rect 9232 25956 9260 25987
rect 10502 25984 10508 26036
rect 10560 26024 10566 26036
rect 10781 26027 10839 26033
rect 10781 26024 10793 26027
rect 10560 25996 10793 26024
rect 10560 25984 10566 25996
rect 10781 25993 10793 25996
rect 10827 25993 10839 26027
rect 10781 25987 10839 25993
rect 10870 25984 10876 26036
rect 10928 25984 10934 26036
rect 15378 26024 15384 26036
rect 12728 25996 15384 26024
rect 12526 25956 12532 25968
rect 4120 25928 4200 25956
rect 9232 25928 12532 25956
rect 4120 25916 4126 25928
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25888 2375 25891
rect 2866 25888 2872 25900
rect 2363 25860 2872 25888
rect 2363 25857 2375 25860
rect 2317 25851 2375 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 4172 25897 4200 25928
rect 12526 25916 12532 25928
rect 12584 25916 12590 25968
rect 3053 25891 3111 25897
rect 3053 25857 3065 25891
rect 3099 25888 3111 25891
rect 4157 25891 4215 25897
rect 3099 25860 4108 25888
rect 3099 25857 3111 25860
rect 3053 25851 3111 25857
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 3237 25823 3295 25829
rect 3237 25820 3249 25823
rect 2832 25792 3249 25820
rect 2832 25780 2838 25792
rect 3237 25789 3249 25792
rect 3283 25820 3295 25823
rect 3602 25820 3608 25832
rect 3283 25792 3608 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 4080 25820 4108 25860
rect 4157 25857 4169 25891
rect 4203 25857 4215 25891
rect 4157 25851 4215 25857
rect 5442 25848 5448 25900
rect 5500 25888 5506 25900
rect 8478 25888 8484 25900
rect 5500 25860 8484 25888
rect 5500 25848 5506 25860
rect 8478 25848 8484 25860
rect 8536 25888 8542 25900
rect 8849 25891 8907 25897
rect 8849 25888 8861 25891
rect 8536 25860 8861 25888
rect 8536 25848 8542 25860
rect 8849 25857 8861 25860
rect 8895 25857 8907 25891
rect 8849 25851 8907 25857
rect 6178 25820 6184 25832
rect 4080 25792 6184 25820
rect 6178 25780 6184 25792
rect 6236 25780 6242 25832
rect 7834 25780 7840 25832
rect 7892 25820 7898 25832
rect 8021 25823 8079 25829
rect 8021 25820 8033 25823
rect 7892 25792 8033 25820
rect 7892 25780 7898 25792
rect 8021 25789 8033 25792
rect 8067 25789 8079 25823
rect 8864 25820 8892 25851
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 12728 25897 12756 25996
rect 15378 25984 15384 25996
rect 15436 25984 15442 26036
rect 15562 25984 15568 26036
rect 15620 26024 15626 26036
rect 15841 26027 15899 26033
rect 15841 26024 15853 26027
rect 15620 25996 15853 26024
rect 15620 25984 15626 25996
rect 15841 25993 15853 25996
rect 15887 25993 15899 26027
rect 18690 26024 18696 26036
rect 15841 25987 15899 25993
rect 17236 25996 18696 26024
rect 14826 25956 14832 25968
rect 14214 25928 14832 25956
rect 14826 25916 14832 25928
rect 14884 25916 14890 25968
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9456 25860 9597 25888
rect 9456 25848 9462 25860
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 12713 25891 12771 25897
rect 12713 25857 12725 25891
rect 12759 25857 12771 25891
rect 12713 25851 12771 25857
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25888 15807 25891
rect 17236 25888 17264 25996
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 19334 25984 19340 26036
rect 19392 25984 19398 26036
rect 19518 25984 19524 26036
rect 19576 26024 19582 26036
rect 20257 26027 20315 26033
rect 20257 26024 20269 26027
rect 19576 25996 20269 26024
rect 19576 25984 19582 25996
rect 20257 25993 20269 25996
rect 20303 25993 20315 26027
rect 20257 25987 20315 25993
rect 20346 25984 20352 26036
rect 20404 25984 20410 26036
rect 20993 26027 21051 26033
rect 20993 25993 21005 26027
rect 21039 26024 21051 26027
rect 21358 26024 21364 26036
rect 21039 25996 21364 26024
rect 21039 25993 21051 25996
rect 20993 25987 21051 25993
rect 21008 25956 21036 25987
rect 21358 25984 21364 25996
rect 21416 26024 21422 26036
rect 22278 26024 22284 26036
rect 21416 25996 22284 26024
rect 21416 25984 21422 25996
rect 22278 25984 22284 25996
rect 22336 25984 22342 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 19306 25928 21036 25956
rect 15795 25860 17264 25888
rect 17589 25891 17647 25897
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 17589 25857 17601 25891
rect 17635 25857 17647 25891
rect 19306 25888 19334 25928
rect 21542 25916 21548 25968
rect 21600 25956 21606 25968
rect 23293 25959 23351 25965
rect 23293 25956 23305 25959
rect 21600 25928 23305 25956
rect 21600 25916 21606 25928
rect 23293 25925 23305 25928
rect 23339 25925 23351 25959
rect 23293 25919 23351 25925
rect 25130 25916 25136 25968
rect 25188 25956 25194 25968
rect 25406 25956 25412 25968
rect 25188 25928 25412 25956
rect 25188 25916 25194 25928
rect 25406 25916 25412 25928
rect 25464 25916 25470 25968
rect 22186 25888 22192 25900
rect 18998 25874 19334 25888
rect 17589 25851 17647 25857
rect 18984 25860 19334 25874
rect 20548 25860 22192 25888
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 8864 25792 9689 25820
rect 8021 25783 8079 25789
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 9769 25823 9827 25829
rect 9769 25789 9781 25823
rect 9815 25789 9827 25823
rect 9769 25783 9827 25789
rect 3418 25712 3424 25764
rect 3476 25712 3482 25764
rect 3620 25752 3648 25780
rect 4617 25755 4675 25761
rect 4617 25752 4629 25755
rect 3620 25724 4629 25752
rect 4617 25721 4629 25724
rect 4663 25721 4675 25755
rect 4617 25715 4675 25721
rect 8570 25712 8576 25764
rect 8628 25752 8634 25764
rect 9784 25752 9812 25783
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10965 25823 11023 25829
rect 10965 25820 10977 25823
rect 9916 25792 10977 25820
rect 9916 25780 9922 25792
rect 10965 25789 10977 25792
rect 11011 25789 11023 25823
rect 10965 25783 11023 25789
rect 11790 25780 11796 25832
rect 11848 25820 11854 25832
rect 11977 25823 12035 25829
rect 11977 25820 11989 25823
rect 11848 25792 11989 25820
rect 11848 25780 11854 25792
rect 11977 25789 11989 25792
rect 12023 25789 12035 25823
rect 11977 25783 12035 25789
rect 12989 25823 13047 25829
rect 12989 25789 13001 25823
rect 13035 25820 13047 25823
rect 14366 25820 14372 25832
rect 13035 25792 14372 25820
rect 13035 25789 13047 25792
rect 12989 25783 13047 25789
rect 14366 25780 14372 25792
rect 14424 25780 14430 25832
rect 14458 25780 14464 25832
rect 14516 25780 14522 25832
rect 16022 25780 16028 25832
rect 16080 25780 16086 25832
rect 8628 25724 9812 25752
rect 8628 25712 8634 25724
rect 4246 25644 4252 25696
rect 4304 25644 4310 25696
rect 10413 25687 10471 25693
rect 10413 25653 10425 25687
rect 10459 25684 10471 25687
rect 11330 25684 11336 25696
rect 10459 25656 11336 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 11330 25644 11336 25656
rect 11388 25644 11394 25696
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 14476 25684 14504 25780
rect 15470 25712 15476 25764
rect 15528 25752 15534 25764
rect 17604 25752 17632 25851
rect 17862 25780 17868 25832
rect 17920 25780 17926 25832
rect 18230 25780 18236 25832
rect 18288 25820 18294 25832
rect 18984 25820 19012 25860
rect 20548 25829 20576 25860
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25888 22431 25891
rect 23382 25888 23388 25900
rect 22419 25860 23388 25888
rect 22419 25857 22431 25860
rect 22373 25851 22431 25857
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 23842 25848 23848 25900
rect 23900 25888 23906 25900
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 23900 25860 23949 25888
rect 23900 25848 23906 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 18288 25792 19012 25820
rect 20533 25823 20591 25829
rect 18288 25780 18294 25792
rect 20533 25789 20545 25823
rect 20579 25789 20591 25823
rect 20533 25783 20591 25789
rect 21269 25823 21327 25829
rect 21269 25789 21281 25823
rect 21315 25820 21327 25823
rect 21634 25820 21640 25832
rect 21315 25792 21640 25820
rect 21315 25789 21327 25792
rect 21269 25783 21327 25789
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22278 25780 22284 25832
rect 22336 25820 22342 25832
rect 22557 25823 22615 25829
rect 22557 25820 22569 25823
rect 22336 25792 22569 25820
rect 22336 25780 22342 25792
rect 22557 25789 22569 25792
rect 22603 25789 22615 25823
rect 22557 25783 22615 25789
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 15528 25724 17632 25752
rect 15528 25712 15534 25724
rect 18966 25712 18972 25764
rect 19024 25752 19030 25764
rect 19889 25755 19947 25761
rect 19889 25752 19901 25755
rect 19024 25724 19901 25752
rect 19024 25712 19030 25724
rect 19889 25721 19901 25724
rect 19935 25721 19947 25755
rect 19889 25715 19947 25721
rect 22094 25712 22100 25764
rect 22152 25752 22158 25764
rect 22830 25752 22836 25764
rect 22152 25724 22836 25752
rect 22152 25712 22158 25724
rect 22830 25712 22836 25724
rect 22888 25712 22894 25764
rect 23477 25755 23535 25761
rect 23477 25721 23489 25755
rect 23523 25752 23535 25755
rect 23750 25752 23756 25764
rect 23523 25724 23756 25752
rect 23523 25721 23535 25724
rect 23477 25715 23535 25721
rect 23750 25712 23756 25724
rect 23808 25712 23814 25764
rect 11480 25656 14504 25684
rect 11480 25644 11486 25656
rect 15194 25644 15200 25696
rect 15252 25684 15258 25696
rect 15381 25687 15439 25693
rect 15381 25684 15393 25687
rect 15252 25656 15393 25684
rect 15252 25644 15258 25656
rect 15381 25653 15393 25656
rect 15427 25653 15439 25687
rect 15381 25647 15439 25653
rect 21174 25644 21180 25696
rect 21232 25684 21238 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21232 25656 22017 25684
rect 21232 25644 21238 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 7088 25483 7146 25489
rect 7088 25449 7100 25483
rect 7134 25480 7146 25483
rect 7466 25480 7472 25492
rect 7134 25452 7472 25480
rect 7134 25449 7146 25452
rect 7088 25443 7146 25449
rect 7466 25440 7472 25452
rect 7524 25480 7530 25492
rect 7650 25480 7656 25492
rect 7524 25452 7656 25480
rect 7524 25440 7530 25452
rect 7650 25440 7656 25452
rect 7708 25440 7714 25492
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 8941 25483 8999 25489
rect 8941 25480 8953 25483
rect 8812 25452 8953 25480
rect 8812 25440 8818 25452
rect 8941 25449 8953 25452
rect 8987 25480 8999 25483
rect 9030 25480 9036 25492
rect 8987 25452 9036 25480
rect 8987 25449 8999 25452
rect 8941 25443 8999 25449
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 11425 25483 11483 25489
rect 11425 25449 11437 25483
rect 11471 25480 11483 25483
rect 11514 25480 11520 25492
rect 11471 25452 11520 25480
rect 11471 25449 11483 25452
rect 11425 25443 11483 25449
rect 11514 25440 11520 25452
rect 11572 25440 11578 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 14737 25483 14795 25489
rect 12492 25452 12572 25480
rect 12492 25440 12498 25452
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7650 25344 7656 25356
rect 6871 25316 7656 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8772 25344 8800 25440
rect 10045 25415 10103 25421
rect 10045 25381 10057 25415
rect 10091 25412 10103 25415
rect 10091 25384 12434 25412
rect 10091 25381 10103 25384
rect 10045 25375 10103 25381
rect 8220 25316 8800 25344
rect 4062 25285 4068 25288
rect 4040 25279 4068 25285
rect 4040 25245 4052 25279
rect 4040 25239 4068 25245
rect 4062 25236 4068 25239
rect 4120 25236 4126 25288
rect 8220 25262 8248 25316
rect 9398 25304 9404 25356
rect 9456 25304 9462 25356
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 10597 25347 10655 25353
rect 10597 25344 10609 25347
rect 9732 25316 10609 25344
rect 9732 25304 9738 25316
rect 10597 25313 10609 25316
rect 10643 25313 10655 25347
rect 10597 25307 10655 25313
rect 11422 25304 11428 25356
rect 11480 25344 11486 25356
rect 11977 25347 12035 25353
rect 11977 25344 11989 25347
rect 11480 25316 11989 25344
rect 11480 25304 11486 25316
rect 11977 25313 11989 25316
rect 12023 25313 12035 25347
rect 11977 25307 12035 25313
rect 8386 25236 8392 25288
rect 8444 25276 8450 25288
rect 10413 25279 10471 25285
rect 10413 25276 10425 25279
rect 8444 25248 10425 25276
rect 8444 25236 8450 25248
rect 10413 25245 10425 25248
rect 10459 25245 10471 25279
rect 10413 25239 10471 25245
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10778 25276 10784 25288
rect 10551 25248 10784 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 12406 25208 12434 25384
rect 12544 25288 12572 25452
rect 14737 25449 14749 25483
rect 14783 25480 14795 25483
rect 16758 25480 16764 25492
rect 14783 25452 16764 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 17770 25440 17776 25492
rect 17828 25480 17834 25492
rect 18049 25483 18107 25489
rect 18049 25480 18061 25483
rect 17828 25452 18061 25480
rect 17828 25440 17834 25452
rect 18049 25449 18061 25452
rect 18095 25480 18107 25483
rect 18230 25480 18236 25492
rect 18095 25452 18236 25480
rect 18095 25449 18107 25452
rect 18049 25443 18107 25449
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 22462 25440 22468 25492
rect 22520 25480 22526 25492
rect 23109 25483 23167 25489
rect 23109 25480 23121 25483
rect 22520 25452 23121 25480
rect 22520 25440 22526 25452
rect 23109 25449 23121 25452
rect 23155 25449 23167 25483
rect 23109 25443 23167 25449
rect 23382 25440 23388 25492
rect 23440 25440 23446 25492
rect 25222 25440 25228 25492
rect 25280 25440 25286 25492
rect 25498 25440 25504 25492
rect 25556 25440 25562 25492
rect 22097 25415 22155 25421
rect 15304 25384 16068 25412
rect 12802 25304 12808 25356
rect 12860 25344 12866 25356
rect 13173 25347 13231 25353
rect 13173 25344 13185 25347
rect 12860 25316 13185 25344
rect 12860 25304 12866 25316
rect 13173 25313 13185 25316
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 13630 25304 13636 25356
rect 13688 25304 13694 25356
rect 15304 25353 15332 25384
rect 15289 25347 15347 25353
rect 15289 25313 15301 25347
rect 15335 25313 15347 25347
rect 15289 25307 15347 25313
rect 15378 25304 15384 25356
rect 15436 25344 15442 25356
rect 15933 25347 15991 25353
rect 15933 25344 15945 25347
rect 15436 25316 15945 25344
rect 15436 25304 15442 25316
rect 15933 25313 15945 25316
rect 15979 25313 15991 25347
rect 16040 25344 16068 25384
rect 22097 25381 22109 25415
rect 22143 25412 22155 25415
rect 24946 25412 24952 25424
rect 22143 25384 24952 25412
rect 22143 25381 22155 25384
rect 22097 25375 22155 25381
rect 24946 25372 24952 25384
rect 25004 25372 25010 25424
rect 16209 25347 16267 25353
rect 16209 25344 16221 25347
rect 16040 25316 16221 25344
rect 15933 25307 15991 25313
rect 16209 25313 16221 25316
rect 16255 25344 16267 25347
rect 16666 25344 16672 25356
rect 16255 25316 16672 25344
rect 16255 25313 16267 25316
rect 16209 25307 16267 25313
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 19058 25304 19064 25356
rect 19116 25344 19122 25356
rect 19889 25347 19947 25353
rect 19889 25344 19901 25347
rect 19116 25316 19901 25344
rect 19116 25304 19122 25316
rect 19889 25313 19901 25316
rect 19935 25313 19947 25347
rect 19889 25307 19947 25313
rect 20070 25304 20076 25356
rect 20128 25304 20134 25356
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 22557 25347 22615 25353
rect 22557 25344 22569 25347
rect 21140 25316 22569 25344
rect 21140 25304 21146 25316
rect 22557 25313 22569 25316
rect 22603 25313 22615 25347
rect 22557 25307 22615 25313
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 22741 25347 22799 25353
rect 22741 25344 22753 25347
rect 22704 25316 22753 25344
rect 22704 25304 22710 25316
rect 22741 25313 22753 25316
rect 22787 25344 22799 25347
rect 23198 25344 23204 25356
rect 22787 25316 23204 25344
rect 22787 25313 22799 25316
rect 22741 25307 22799 25313
rect 23198 25304 23204 25316
rect 23256 25304 23262 25356
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 13078 25236 13084 25288
rect 13136 25276 13142 25288
rect 13648 25276 13676 25304
rect 13136 25248 13676 25276
rect 13136 25236 13142 25248
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19484 25248 19809 25276
rect 19484 25236 19490 25248
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 21634 25236 21640 25288
rect 21692 25276 21698 25288
rect 22465 25279 22523 25285
rect 22465 25276 22477 25279
rect 21692 25248 22477 25276
rect 21692 25236 21698 25248
rect 22465 25245 22477 25248
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 22830 25236 22836 25288
rect 22888 25276 22894 25288
rect 24673 25279 24731 25285
rect 24673 25276 24685 25279
rect 22888 25248 24685 25276
rect 22888 25236 22894 25248
rect 24673 25245 24685 25248
rect 24719 25245 24731 25279
rect 24673 25239 24731 25245
rect 13630 25208 13636 25220
rect 8496 25180 9904 25208
rect 12406 25180 13636 25208
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 4111 25143 4169 25149
rect 4111 25140 4123 25143
rect 4028 25112 4123 25140
rect 4028 25100 4034 25112
rect 4111 25109 4123 25112
rect 4157 25109 4169 25143
rect 4111 25103 4169 25109
rect 6638 25100 6644 25152
rect 6696 25140 6702 25152
rect 8496 25140 8524 25180
rect 6696 25112 8524 25140
rect 6696 25100 6702 25112
rect 8570 25100 8576 25152
rect 8628 25100 8634 25152
rect 9876 25140 9904 25180
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 17770 25208 17776 25220
rect 17434 25180 17776 25208
rect 17770 25168 17776 25180
rect 17828 25168 17834 25220
rect 22370 25168 22376 25220
rect 22428 25208 22434 25220
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 22428 25180 23857 25208
rect 22428 25168 22434 25180
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 23845 25171 23903 25177
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 9876 25112 11069 25140
rect 11057 25109 11069 25112
rect 11103 25140 11115 25143
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 11103 25112 11897 25140
rect 11103 25109 11115 25112
rect 11057 25103 11115 25109
rect 11885 25109 11897 25112
rect 11931 25140 11943 25143
rect 11974 25140 11980 25152
rect 11931 25112 11980 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 12989 25143 13047 25149
rect 12989 25140 13001 25143
rect 12860 25112 13001 25140
rect 12860 25100 12866 25112
rect 12989 25109 13001 25112
rect 13035 25109 13047 25143
rect 12989 25103 13047 25109
rect 15102 25100 15108 25152
rect 15160 25100 15166 25152
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 16850 25140 16856 25152
rect 15243 25112 16856 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 17681 25143 17739 25149
rect 17681 25140 17693 25143
rect 17092 25112 17693 25140
rect 17092 25100 17098 25112
rect 17681 25109 17693 25112
rect 17727 25140 17739 25143
rect 17862 25140 17868 25152
rect 17727 25112 17868 25140
rect 17727 25109 17739 25112
rect 17681 25103 17739 25109
rect 17862 25100 17868 25112
rect 17920 25100 17926 25152
rect 18233 25143 18291 25149
rect 18233 25109 18245 25143
rect 18279 25140 18291 25143
rect 18322 25140 18328 25152
rect 18279 25112 18328 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 18506 25100 18512 25152
rect 18564 25140 18570 25152
rect 18690 25140 18696 25152
rect 18564 25112 18696 25140
rect 18564 25100 18570 25112
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 19426 25100 19432 25152
rect 19484 25100 19490 25152
rect 23934 25100 23940 25152
rect 23992 25100 23998 25152
rect 24026 25100 24032 25152
rect 24084 25140 24090 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 24084 25112 24777 25140
rect 24084 25100 24090 25112
rect 24765 25109 24777 25112
rect 24811 25109 24823 25143
rect 24765 25103 24823 25109
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 4246 24896 4252 24948
rect 4304 24936 4310 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 4304 24908 5457 24936
rect 4304 24896 4310 24908
rect 5445 24905 5457 24908
rect 5491 24905 5503 24939
rect 5445 24899 5503 24905
rect 7834 24896 7840 24948
rect 7892 24936 7898 24948
rect 8021 24939 8079 24945
rect 8021 24936 8033 24939
rect 7892 24908 8033 24936
rect 7892 24896 7898 24908
rect 8021 24905 8033 24908
rect 8067 24905 8079 24939
rect 8021 24899 8079 24905
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 15197 24939 15255 24945
rect 15197 24936 15209 24939
rect 12676 24908 15209 24936
rect 12676 24896 12682 24908
rect 15197 24905 15209 24908
rect 15243 24905 15255 24939
rect 15197 24899 15255 24905
rect 16850 24896 16856 24948
rect 16908 24896 16914 24948
rect 17678 24896 17684 24948
rect 17736 24936 17742 24948
rect 18506 24936 18512 24948
rect 17736 24908 18512 24936
rect 17736 24896 17742 24908
rect 18506 24896 18512 24908
rect 18564 24896 18570 24948
rect 19886 24896 19892 24948
rect 19944 24936 19950 24948
rect 20625 24939 20683 24945
rect 20625 24936 20637 24939
rect 19944 24908 20637 24936
rect 19944 24896 19950 24908
rect 20625 24905 20637 24908
rect 20671 24905 20683 24939
rect 20625 24899 20683 24905
rect 7466 24828 7472 24880
rect 7524 24868 7530 24880
rect 9217 24871 9275 24877
rect 7524 24840 8340 24868
rect 7524 24828 7530 24840
rect 5810 24800 5816 24812
rect 5106 24772 5816 24800
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 7374 24760 7380 24812
rect 7432 24760 7438 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 8312 24800 8340 24840
rect 9217 24837 9229 24871
rect 9263 24868 9275 24871
rect 12069 24871 12127 24877
rect 9263 24840 10088 24868
rect 9263 24837 9275 24840
rect 9217 24831 9275 24837
rect 10060 24809 10088 24840
rect 12069 24837 12081 24871
rect 12115 24868 12127 24871
rect 12805 24871 12863 24877
rect 12115 24840 12756 24868
rect 12115 24837 12127 24840
rect 12069 24831 12127 24837
rect 10045 24803 10103 24809
rect 7800 24772 8248 24800
rect 8312 24772 9444 24800
rect 7800 24760 7806 24772
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24732 3755 24735
rect 3973 24735 4031 24741
rect 3743 24704 3832 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 3804 24596 3832 24704
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 5994 24732 6000 24744
rect 4019 24704 6000 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 5994 24692 6000 24704
rect 6052 24692 6058 24744
rect 7392 24732 7420 24760
rect 8110 24732 8116 24744
rect 7392 24704 8116 24732
rect 8110 24692 8116 24704
rect 8168 24692 8174 24744
rect 8220 24741 8248 24772
rect 8205 24735 8263 24741
rect 8205 24701 8217 24735
rect 8251 24701 8263 24735
rect 8205 24695 8263 24701
rect 9306 24692 9312 24744
rect 9364 24692 9370 24744
rect 9416 24741 9444 24772
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24800 12219 24803
rect 12434 24800 12440 24812
rect 12207 24772 12440 24800
rect 12207 24769 12219 24772
rect 12161 24763 12219 24769
rect 12434 24760 12440 24772
rect 12492 24760 12498 24812
rect 12728 24800 12756 24840
rect 12805 24837 12817 24871
rect 12851 24868 12863 24871
rect 12894 24868 12900 24880
rect 12851 24840 12900 24868
rect 12851 24837 12863 24840
rect 12805 24831 12863 24837
rect 12894 24828 12900 24840
rect 12952 24868 12958 24880
rect 13078 24868 13084 24880
rect 12952 24840 13084 24868
rect 12952 24828 12958 24840
rect 13078 24828 13084 24840
rect 13136 24828 13142 24880
rect 14936 24840 15424 24868
rect 13173 24803 13231 24809
rect 12728 24772 13032 24800
rect 13004 24744 13032 24772
rect 13173 24769 13185 24803
rect 13219 24800 13231 24803
rect 13538 24800 13544 24812
rect 13219 24772 13544 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 13814 24760 13820 24812
rect 13872 24760 13878 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14108 24772 14565 24800
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 10134 24692 10140 24744
rect 10192 24732 10198 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 10192 24704 12265 24732
rect 10192 24692 10198 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 12986 24692 12992 24744
rect 13044 24692 13050 24744
rect 13556 24732 13584 24760
rect 14108 24741 14136 24772
rect 14553 24769 14565 24772
rect 14599 24800 14611 24803
rect 14936 24800 14964 24840
rect 14599 24772 14964 24800
rect 14599 24769 14611 24772
rect 14553 24763 14611 24769
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 15068 24772 15301 24800
rect 15068 24760 15074 24772
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15396 24800 15424 24840
rect 16390 24828 16396 24880
rect 16448 24868 16454 24880
rect 17126 24868 17132 24880
rect 16448 24840 17132 24868
rect 16448 24828 16454 24840
rect 17126 24828 17132 24840
rect 17184 24868 17190 24880
rect 17221 24871 17279 24877
rect 17221 24868 17233 24871
rect 17184 24840 17233 24868
rect 17184 24828 17190 24840
rect 17221 24837 17233 24840
rect 17267 24837 17279 24871
rect 17221 24831 17279 24837
rect 23198 24828 23204 24880
rect 23256 24828 23262 24880
rect 24486 24868 24492 24880
rect 24426 24840 24492 24868
rect 24486 24828 24492 24840
rect 24544 24868 24550 24880
rect 25222 24868 25228 24880
rect 24544 24840 25228 24868
rect 24544 24828 24550 24840
rect 25222 24828 25228 24840
rect 25280 24828 25286 24880
rect 15396 24772 16436 24800
rect 15289 24763 15347 24769
rect 13909 24735 13967 24741
rect 13909 24732 13921 24735
rect 13556 24704 13921 24732
rect 13909 24701 13921 24704
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 14093 24735 14151 24741
rect 14093 24701 14105 24735
rect 14139 24701 14151 24735
rect 14093 24695 14151 24701
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 15381 24735 15439 24741
rect 15381 24732 15393 24735
rect 14424 24704 15393 24732
rect 14424 24692 14430 24704
rect 15381 24701 15393 24704
rect 15427 24701 15439 24735
rect 16408 24732 16436 24772
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 18322 24800 18328 24812
rect 17920 24772 18328 24800
rect 17920 24760 17926 24772
rect 18322 24760 18328 24772
rect 18380 24800 18386 24812
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 18380 24772 18429 24800
rect 18380 24760 18386 24772
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 18874 24760 18880 24812
rect 18932 24760 18938 24812
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 22830 24800 22836 24812
rect 20680 24772 22836 24800
rect 20680 24760 20686 24772
rect 22830 24760 22836 24772
rect 22888 24800 22894 24812
rect 22925 24803 22983 24809
rect 22925 24800 22937 24803
rect 22888 24772 22937 24800
rect 22888 24760 22894 24772
rect 22925 24769 22937 24772
rect 22971 24769 22983 24803
rect 22925 24763 22983 24769
rect 25317 24803 25375 24809
rect 25317 24769 25329 24803
rect 25363 24800 25375 24803
rect 25498 24800 25504 24812
rect 25363 24772 25504 24800
rect 25363 24769 25375 24772
rect 25317 24763 25375 24769
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 17494 24732 17500 24744
rect 16408 24704 17500 24732
rect 15381 24695 15439 24701
rect 17494 24692 17500 24704
rect 17552 24692 17558 24744
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18601 24735 18659 24741
rect 18601 24732 18613 24735
rect 17828 24704 18613 24732
rect 17828 24692 17834 24704
rect 18601 24701 18613 24704
rect 18647 24732 18659 24735
rect 18782 24732 18788 24744
rect 18647 24704 18788 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 18782 24692 18788 24704
rect 18840 24692 18846 24744
rect 18892 24732 18920 24760
rect 20530 24732 20536 24744
rect 18892 24704 20536 24732
rect 20530 24692 20536 24704
rect 20588 24732 20594 24744
rect 20717 24735 20775 24741
rect 20717 24732 20729 24735
rect 20588 24704 20729 24732
rect 20588 24692 20594 24704
rect 20717 24701 20729 24704
rect 20763 24701 20775 24735
rect 20717 24695 20775 24701
rect 20809 24735 20867 24741
rect 20809 24701 20821 24735
rect 20855 24701 20867 24735
rect 20809 24695 20867 24701
rect 7653 24667 7711 24673
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8386 24664 8392 24676
rect 7699 24636 8392 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8386 24624 8392 24636
rect 8444 24624 8450 24676
rect 11701 24667 11759 24673
rect 11701 24664 11713 24667
rect 8496 24636 11713 24664
rect 3970 24596 3976 24608
rect 3804 24568 3976 24596
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 5810 24556 5816 24608
rect 5868 24556 5874 24608
rect 7742 24556 7748 24608
rect 7800 24596 7806 24608
rect 8496 24596 8524 24636
rect 11701 24633 11713 24636
rect 11747 24633 11759 24667
rect 11701 24627 11759 24633
rect 12618 24624 12624 24676
rect 12676 24664 12682 24676
rect 13449 24667 13507 24673
rect 12676 24636 13032 24664
rect 12676 24624 12682 24636
rect 7800 24568 8524 24596
rect 8849 24599 8907 24605
rect 7800 24556 7806 24568
rect 8849 24565 8861 24599
rect 8895 24596 8907 24599
rect 11146 24596 11152 24608
rect 8895 24568 11152 24596
rect 8895 24565 8907 24568
rect 8849 24559 8907 24565
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 12250 24556 12256 24608
rect 12308 24596 12314 24608
rect 12894 24596 12900 24608
rect 12308 24568 12900 24596
rect 12308 24556 12314 24568
rect 12894 24556 12900 24568
rect 12952 24556 12958 24608
rect 13004 24596 13032 24636
rect 13449 24633 13461 24667
rect 13495 24664 13507 24667
rect 15102 24664 15108 24676
rect 13495 24636 15108 24664
rect 13495 24633 13507 24636
rect 13449 24627 13507 24633
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 18874 24664 18880 24676
rect 16316 24636 18880 24664
rect 13722 24596 13728 24608
rect 13004 24568 13728 24596
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14829 24599 14887 24605
rect 14829 24565 14841 24599
rect 14875 24596 14887 24599
rect 16316 24596 16344 24636
rect 18874 24624 18880 24636
rect 18932 24624 18938 24676
rect 20438 24624 20444 24676
rect 20496 24664 20502 24676
rect 20622 24664 20628 24676
rect 20496 24636 20628 24664
rect 20496 24624 20502 24636
rect 20622 24624 20628 24636
rect 20680 24664 20686 24676
rect 20824 24664 20852 24695
rect 24670 24692 24676 24744
rect 24728 24692 24734 24744
rect 20680 24636 20852 24664
rect 20680 24624 20686 24636
rect 25130 24624 25136 24676
rect 25188 24624 25194 24676
rect 14875 24568 16344 24596
rect 14875 24565 14887 24568
rect 14829 24559 14887 24565
rect 16390 24556 16396 24608
rect 16448 24556 16454 24608
rect 18049 24599 18107 24605
rect 18049 24565 18061 24599
rect 18095 24596 18107 24599
rect 18506 24596 18512 24608
rect 18095 24568 18512 24596
rect 18095 24565 18107 24568
rect 18049 24559 18107 24565
rect 18506 24556 18512 24568
rect 18564 24556 18570 24608
rect 20257 24599 20315 24605
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 23382 24596 23388 24608
rect 20303 24568 23388 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 3237 24395 3295 24401
rect 3237 24361 3249 24395
rect 3283 24361 3295 24395
rect 3237 24355 3295 24361
rect 3252 24324 3280 24355
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3421 24395 3479 24401
rect 3421 24392 3433 24395
rect 3384 24364 3433 24392
rect 3384 24352 3390 24364
rect 3421 24361 3433 24364
rect 3467 24361 3479 24395
rect 4430 24392 4436 24404
rect 3421 24355 3479 24361
rect 3528 24364 4436 24392
rect 3528 24324 3556 24364
rect 4430 24352 4436 24364
rect 4488 24392 4494 24404
rect 5721 24395 5779 24401
rect 5721 24392 5733 24395
rect 4488 24364 5733 24392
rect 4488 24352 4494 24364
rect 5721 24361 5733 24364
rect 5767 24361 5779 24395
rect 5721 24355 5779 24361
rect 6178 24352 6184 24404
rect 6236 24352 6242 24404
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 8757 24395 8815 24401
rect 8757 24392 8769 24395
rect 8536 24364 8769 24392
rect 8536 24352 8542 24364
rect 8757 24361 8769 24364
rect 8803 24392 8815 24395
rect 9306 24392 9312 24404
rect 8803 24364 9312 24392
rect 8803 24361 8815 24364
rect 8757 24355 8815 24361
rect 9306 24352 9312 24364
rect 9364 24352 9370 24404
rect 10226 24352 10232 24404
rect 10284 24392 10290 24404
rect 13633 24395 13691 24401
rect 10284 24364 11468 24392
rect 10284 24352 10290 24364
rect 3252 24296 3556 24324
rect 6362 24284 6368 24336
rect 6420 24284 6426 24336
rect 8570 24284 8576 24336
rect 8628 24324 8634 24336
rect 8628 24296 11376 24324
rect 8628 24284 8634 24296
rect 4246 24216 4252 24268
rect 4304 24216 4310 24268
rect 6380 24256 6408 24284
rect 9858 24256 9864 24268
rect 6380 24228 9864 24256
rect 9858 24216 9864 24228
rect 9916 24216 9922 24268
rect 10045 24259 10103 24265
rect 10045 24225 10057 24259
rect 10091 24256 10103 24259
rect 11054 24256 11060 24268
rect 10091 24228 11060 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11348 24265 11376 24296
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24225 11391 24259
rect 11440 24256 11468 24364
rect 13633 24361 13645 24395
rect 13679 24392 13691 24395
rect 15378 24392 15384 24404
rect 13679 24364 15384 24392
rect 13679 24361 13691 24364
rect 13633 24355 13691 24361
rect 12158 24284 12164 24336
rect 12216 24324 12222 24336
rect 13722 24324 13728 24336
rect 12216 24296 13728 24324
rect 12216 24284 12222 24296
rect 13722 24284 13728 24296
rect 13780 24284 13786 24336
rect 12529 24259 12587 24265
rect 12529 24256 12541 24259
rect 11440 24228 12541 24256
rect 11333 24219 11391 24225
rect 12529 24225 12541 24228
rect 12575 24225 12587 24259
rect 12529 24219 12587 24225
rect 12802 24216 12808 24268
rect 12860 24256 12866 24268
rect 13173 24259 13231 24265
rect 13173 24256 13185 24259
rect 12860 24228 13185 24256
rect 12860 24216 12866 24228
rect 13173 24225 13185 24228
rect 13219 24225 13231 24259
rect 13832 24256 13860 24364
rect 15378 24352 15384 24364
rect 15436 24392 15442 24404
rect 15930 24392 15936 24404
rect 15436 24364 15936 24392
rect 15436 24352 15442 24364
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 17589 24395 17647 24401
rect 17589 24361 17601 24395
rect 17635 24392 17647 24395
rect 20714 24392 20720 24404
rect 17635 24364 20720 24392
rect 17635 24361 17647 24364
rect 17589 24355 17647 24361
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 24670 24284 24676 24336
rect 24728 24324 24734 24336
rect 24728 24296 25176 24324
rect 24728 24284 24734 24296
rect 13173 24219 13231 24225
rect 13740 24228 13860 24256
rect 16853 24259 16911 24265
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2774 24188 2780 24200
rect 2271 24160 2780 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 2961 24191 3019 24197
rect 2961 24157 2973 24191
rect 3007 24188 3019 24191
rect 3510 24188 3516 24200
rect 3007 24160 3516 24188
rect 3007 24157 3019 24160
rect 2961 24151 3019 24157
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24120 2743 24123
rect 2976 24120 3004 24151
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 3970 24148 3976 24200
rect 4028 24148 4034 24200
rect 6365 24191 6423 24197
rect 6365 24157 6377 24191
rect 6411 24188 6423 24191
rect 7098 24188 7104 24200
rect 6411 24160 7104 24188
rect 6411 24157 6423 24160
rect 6365 24151 6423 24157
rect 7098 24148 7104 24160
rect 7156 24148 7162 24200
rect 11146 24148 11152 24200
rect 11204 24148 11210 24200
rect 11241 24191 11299 24197
rect 11241 24157 11253 24191
rect 11287 24188 11299 24191
rect 12618 24188 12624 24200
rect 11287 24160 12624 24188
rect 11287 24157 11299 24160
rect 11241 24151 11299 24157
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 2731 24092 3004 24120
rect 3528 24120 3556 24148
rect 4522 24120 4528 24132
rect 3528 24092 4528 24120
rect 2731 24089 2743 24092
rect 2685 24083 2743 24089
rect 4522 24080 4528 24092
rect 4580 24080 4586 24132
rect 5810 24120 5816 24132
rect 5474 24092 5816 24120
rect 5810 24080 5816 24092
rect 5868 24120 5874 24132
rect 6546 24120 6552 24132
rect 5868 24092 6552 24120
rect 5868 24080 5874 24092
rect 6546 24080 6552 24092
rect 6604 24120 6610 24132
rect 6733 24123 6791 24129
rect 6733 24120 6745 24123
rect 6604 24092 6745 24120
rect 6604 24080 6610 24092
rect 6733 24089 6745 24092
rect 6779 24120 6791 24123
rect 9030 24120 9036 24132
rect 6779 24092 9036 24120
rect 6779 24089 6791 24092
rect 6733 24083 6791 24089
rect 9030 24080 9036 24092
rect 9088 24080 9094 24132
rect 9861 24123 9919 24129
rect 9861 24089 9873 24123
rect 9907 24089 9919 24123
rect 9861 24083 9919 24089
rect 12345 24123 12403 24129
rect 12345 24089 12357 24123
rect 12391 24120 12403 24123
rect 13740 24120 13768 24228
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 16942 24256 16948 24268
rect 16899 24228 16948 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 17034 24216 17040 24268
rect 17092 24216 17098 24268
rect 17310 24216 17316 24268
rect 17368 24256 17374 24268
rect 18233 24259 18291 24265
rect 18233 24256 18245 24259
rect 17368 24228 18245 24256
rect 17368 24216 17374 24228
rect 18233 24225 18245 24228
rect 18279 24225 18291 24259
rect 18233 24219 18291 24225
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 22830 24256 22836 24268
rect 19751 24228 22836 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 23845 24259 23903 24265
rect 23845 24225 23857 24259
rect 23891 24256 23903 24259
rect 24854 24256 24860 24268
rect 23891 24228 24860 24256
rect 23891 24225 23903 24228
rect 23845 24219 23903 24225
rect 24854 24216 24860 24228
rect 24912 24216 24918 24268
rect 25148 24265 25176 24296
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 17773 24191 17831 24197
rect 17773 24157 17785 24191
rect 17819 24157 17831 24191
rect 17773 24151 17831 24157
rect 12391 24092 13768 24120
rect 12391 24089 12403 24092
rect 12345 24083 12403 24089
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 2041 24055 2099 24061
rect 2041 24052 2053 24055
rect 1912 24024 2053 24052
rect 1912 24012 1918 24024
rect 2041 24021 2053 24024
rect 2087 24021 2099 24055
rect 2041 24015 2099 24021
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8812 24024 9413 24052
rect 8812 24012 8818 24024
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 9766 24012 9772 24064
rect 9824 24012 9830 24064
rect 9876 24052 9904 24083
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 14277 24123 14335 24129
rect 14277 24120 14289 24123
rect 13872 24092 14289 24120
rect 13872 24080 13878 24092
rect 14277 24089 14289 24092
rect 14323 24089 14335 24123
rect 14277 24083 14335 24089
rect 14734 24080 14740 24132
rect 14792 24120 14798 24132
rect 17788 24120 17816 24151
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21784 24160 22017 24188
rect 21784 24148 21790 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24188 22799 24191
rect 23290 24188 23296 24200
rect 22787 24160 23296 24188
rect 22787 24157 22799 24160
rect 22741 24151 22799 24157
rect 23290 24148 23296 24160
rect 23348 24148 23354 24200
rect 24394 24148 24400 24200
rect 24452 24188 24458 24200
rect 25041 24191 25099 24197
rect 25041 24188 25053 24191
rect 24452 24160 25053 24188
rect 24452 24148 24458 24160
rect 25041 24157 25053 24160
rect 25087 24157 25099 24191
rect 25041 24151 25099 24157
rect 14792 24092 17816 24120
rect 14792 24080 14798 24092
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19886 24120 19892 24132
rect 18840 24092 19892 24120
rect 18840 24080 18846 24092
rect 19886 24080 19892 24092
rect 19944 24120 19950 24132
rect 19981 24123 20039 24129
rect 19981 24120 19993 24123
rect 19944 24092 19993 24120
rect 19944 24080 19950 24092
rect 19981 24089 19993 24092
rect 20027 24089 20039 24123
rect 21358 24120 21364 24132
rect 21206 24092 21364 24120
rect 19981 24083 20039 24089
rect 21358 24080 21364 24092
rect 21416 24080 21422 24132
rect 24946 24080 24952 24132
rect 25004 24080 25010 24132
rect 10413 24055 10471 24061
rect 10413 24052 10425 24055
rect 9876 24024 10425 24052
rect 10413 24021 10425 24024
rect 10459 24052 10471 24055
rect 10686 24052 10692 24064
rect 10459 24024 10692 24052
rect 10459 24021 10471 24024
rect 10413 24015 10471 24021
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 10781 24055 10839 24061
rect 10781 24021 10793 24055
rect 10827 24052 10839 24055
rect 10962 24052 10968 24064
rect 10827 24024 10968 24052
rect 10827 24021 10839 24024
rect 10781 24015 10839 24021
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 11974 24012 11980 24064
rect 12032 24012 12038 24064
rect 12066 24012 12072 24064
rect 12124 24052 12130 24064
rect 12437 24055 12495 24061
rect 12437 24052 12449 24055
rect 12124 24024 12449 24052
rect 12124 24012 12130 24024
rect 12437 24021 12449 24024
rect 12483 24021 12495 24055
rect 12437 24015 12495 24021
rect 16393 24055 16451 24061
rect 16393 24021 16405 24055
rect 16439 24052 16451 24055
rect 16666 24052 16672 24064
rect 16439 24024 16672 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 18049 24055 18107 24061
rect 18049 24052 18061 24055
rect 17552 24024 18061 24052
rect 17552 24012 17558 24024
rect 18049 24021 18061 24024
rect 18095 24021 18107 24055
rect 18049 24015 18107 24021
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 21453 24055 21511 24061
rect 21453 24052 21465 24055
rect 20312 24024 21465 24052
rect 20312 24012 20318 24024
rect 21453 24021 21465 24024
rect 21499 24021 21511 24055
rect 21453 24015 21511 24021
rect 22094 24012 22100 24064
rect 22152 24012 22158 24064
rect 22370 24012 22376 24064
rect 22428 24052 22434 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 22428 24024 24593 24052
rect 22428 24012 22434 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 5994 23808 6000 23860
rect 6052 23808 6058 23860
rect 6457 23851 6515 23857
rect 6457 23817 6469 23851
rect 6503 23848 6515 23851
rect 6546 23848 6552 23860
rect 6503 23820 6552 23848
rect 6503 23817 6515 23820
rect 6457 23811 6515 23817
rect 6472 23780 6500 23811
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 7650 23808 7656 23860
rect 7708 23848 7714 23860
rect 9950 23848 9956 23860
rect 7708 23820 9956 23848
rect 7708 23808 7714 23820
rect 9950 23808 9956 23820
rect 10008 23848 10014 23860
rect 10686 23848 10692 23860
rect 10008 23820 10692 23848
rect 10008 23808 10014 23820
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 11793 23851 11851 23857
rect 11793 23848 11805 23851
rect 11296 23820 11805 23848
rect 11296 23808 11302 23820
rect 11793 23817 11805 23820
rect 11839 23848 11851 23851
rect 12066 23848 12072 23860
rect 11839 23820 12072 23848
rect 11839 23817 11851 23820
rect 11793 23811 11851 23817
rect 12066 23808 12072 23820
rect 12124 23808 12130 23860
rect 12342 23808 12348 23860
rect 12400 23848 12406 23860
rect 12437 23851 12495 23857
rect 12437 23848 12449 23851
rect 12400 23820 12449 23848
rect 12400 23808 12406 23820
rect 12437 23817 12449 23820
rect 12483 23848 12495 23851
rect 13538 23848 13544 23860
rect 12483 23820 13544 23848
rect 12483 23817 12495 23820
rect 12437 23811 12495 23817
rect 13538 23808 13544 23820
rect 13596 23808 13602 23860
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 18690 23848 18696 23860
rect 13964 23820 18696 23848
rect 13964 23808 13970 23820
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 19886 23808 19892 23860
rect 19944 23848 19950 23860
rect 19944 23820 20484 23848
rect 19944 23808 19950 23820
rect 5750 23752 6500 23780
rect 1762 23672 1768 23724
rect 1820 23672 1826 23724
rect 7668 23721 7696 23808
rect 9766 23740 9772 23792
rect 9824 23780 9830 23792
rect 9861 23783 9919 23789
rect 9861 23780 9873 23783
rect 9824 23752 9873 23780
rect 9824 23740 9830 23752
rect 9861 23749 9873 23752
rect 9907 23749 9919 23783
rect 9861 23743 9919 23749
rect 10502 23740 10508 23792
rect 10560 23780 10566 23792
rect 11256 23780 11284 23808
rect 10560 23752 11284 23780
rect 10560 23740 10566 23752
rect 7653 23715 7711 23721
rect 7653 23681 7665 23715
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 10321 23715 10379 23721
rect 10321 23712 10333 23715
rect 9088 23684 10333 23712
rect 9088 23672 9094 23684
rect 10321 23681 10333 23684
rect 10367 23712 10379 23715
rect 11238 23712 11244 23724
rect 10367 23684 11244 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 11238 23672 11244 23684
rect 11296 23672 11302 23724
rect 20456 23712 20484 23820
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 20588 23820 25145 23848
rect 20588 23808 20594 23820
rect 25133 23817 25145 23820
rect 25179 23817 25191 23851
rect 25133 23811 25191 23817
rect 20622 23740 20628 23792
rect 20680 23780 20686 23792
rect 23201 23783 23259 23789
rect 23201 23780 23213 23783
rect 20680 23752 23213 23780
rect 20680 23740 20686 23752
rect 23201 23749 23213 23752
rect 23247 23780 23259 23783
rect 23474 23780 23480 23792
rect 23247 23752 23480 23780
rect 23247 23749 23259 23752
rect 23201 23743 23259 23749
rect 23474 23740 23480 23752
rect 23532 23740 23538 23792
rect 24486 23780 24492 23792
rect 24426 23752 24492 23780
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 21177 23715 21235 23721
rect 1302 23604 1308 23656
rect 1360 23644 1366 23656
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 1360 23616 2053 23644
rect 1360 23604 1366 23616
rect 2041 23613 2053 23616
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4249 23647 4307 23653
rect 4249 23644 4261 23647
rect 4028 23616 4261 23644
rect 4028 23604 4034 23616
rect 4249 23613 4261 23616
rect 4295 23613 4307 23647
rect 4249 23607 4307 23613
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 7558 23644 7564 23656
rect 4571 23616 7564 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 4264 23508 4292 23607
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7929 23647 7987 23653
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 8570 23644 8576 23656
rect 7975 23616 8576 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 10870 23604 10876 23656
rect 10928 23604 10934 23656
rect 11698 23604 11704 23656
rect 11756 23644 11762 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 11756 23616 12173 23644
rect 11756 23604 11762 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12492 23616 12541 23644
rect 12492 23604 12498 23616
rect 12529 23613 12541 23616
rect 12575 23644 12587 23647
rect 13446 23644 13452 23656
rect 12575 23616 13452 23644
rect 12575 23613 12587 23616
rect 12529 23607 12587 23613
rect 13446 23604 13452 23616
rect 13504 23604 13510 23656
rect 17034 23604 17040 23656
rect 17092 23604 17098 23656
rect 18598 23604 18604 23656
rect 18656 23644 18662 23656
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 18656 23616 18797 23644
rect 18656 23604 18662 23616
rect 18785 23613 18797 23616
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19794 23644 19800 23656
rect 19107 23616 19800 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 19794 23604 19800 23616
rect 19852 23604 19858 23656
rect 20180 23644 20208 23698
rect 20456 23684 20944 23712
rect 20180 23616 20576 23644
rect 9950 23536 9956 23588
rect 10008 23576 10014 23588
rect 11609 23579 11667 23585
rect 11609 23576 11621 23579
rect 10008 23548 11621 23576
rect 10008 23536 10014 23548
rect 11609 23545 11621 23548
rect 11655 23576 11667 23579
rect 16482 23576 16488 23588
rect 11655 23548 16488 23576
rect 11655 23545 11667 23548
rect 11609 23539 11667 23545
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 20548 23576 20576 23616
rect 20806 23604 20812 23656
rect 20864 23604 20870 23656
rect 20916 23644 20944 23684
rect 21177 23681 21189 23715
rect 21223 23712 21235 23715
rect 21358 23712 21364 23724
rect 21223 23684 21364 23712
rect 21223 23681 21235 23684
rect 21177 23675 21235 23681
rect 21358 23672 21364 23684
rect 21416 23712 21422 23724
rect 21545 23715 21603 23721
rect 21545 23712 21557 23715
rect 21416 23684 21557 23712
rect 21416 23672 21422 23684
rect 21545 23681 21557 23684
rect 21591 23681 21603 23715
rect 21545 23675 21603 23681
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 22830 23712 22836 23724
rect 22060 23684 22836 23712
rect 22060 23672 22066 23684
rect 22830 23672 22836 23684
rect 22888 23712 22894 23724
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 22888 23684 22937 23712
rect 22888 23672 22894 23684
rect 22925 23681 22937 23684
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 25314 23672 25320 23724
rect 25372 23672 25378 23724
rect 20916 23616 24348 23644
rect 24320 23588 24348 23616
rect 21358 23576 21364 23588
rect 20548 23548 21364 23576
rect 21358 23536 21364 23548
rect 21416 23536 21422 23588
rect 24302 23536 24308 23588
rect 24360 23536 24366 23588
rect 5718 23508 5724 23520
rect 4264 23480 5724 23508
rect 5718 23468 5724 23480
rect 5776 23468 5782 23520
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 9401 23511 9459 23517
rect 9401 23508 9413 23511
rect 6880 23480 9413 23508
rect 6880 23468 6886 23480
rect 9401 23477 9413 23480
rect 9447 23508 9459 23511
rect 10134 23508 10140 23520
rect 9447 23480 10140 23508
rect 9447 23477 9459 23480
rect 9401 23471 9459 23477
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 11790 23508 11796 23520
rect 10836 23480 11796 23508
rect 10836 23468 10842 23480
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 17494 23468 17500 23520
rect 17552 23508 17558 23520
rect 20806 23508 20812 23520
rect 17552 23480 20812 23508
rect 17552 23468 17558 23480
rect 20806 23468 20812 23480
rect 20864 23468 20870 23520
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24670 23508 24676 23520
rect 23716 23480 24676 23508
rect 23716 23468 23722 23480
rect 24670 23468 24676 23480
rect 24728 23468 24734 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 2038 23264 2044 23316
rect 2096 23264 2102 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2924 23276 3157 23304
rect 2924 23264 2930 23276
rect 3145 23273 3157 23276
rect 3191 23273 3203 23307
rect 3145 23267 3203 23273
rect 7558 23264 7564 23316
rect 7616 23264 7622 23316
rect 7929 23307 7987 23313
rect 7929 23273 7941 23307
rect 7975 23304 7987 23307
rect 9030 23304 9036 23316
rect 7975 23276 9036 23304
rect 7975 23273 7987 23276
rect 7929 23267 7987 23273
rect 2866 23128 2872 23180
rect 2924 23168 2930 23180
rect 2961 23171 3019 23177
rect 2961 23168 2973 23171
rect 2924 23140 2973 23168
rect 2924 23128 2930 23140
rect 2961 23137 2973 23140
rect 3007 23168 3019 23171
rect 3326 23168 3332 23180
rect 3007 23140 3332 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 5718 23128 5724 23180
rect 5776 23168 5782 23180
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5776 23140 5825 23168
rect 5776 23128 5782 23140
rect 5813 23137 5825 23140
rect 5859 23168 5871 23171
rect 6454 23168 6460 23180
rect 5859 23140 6460 23168
rect 5859 23137 5871 23140
rect 5813 23131 5871 23137
rect 6454 23128 6460 23140
rect 6512 23128 6518 23180
rect 7834 23168 7840 23180
rect 7208 23140 7840 23168
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 2823 23072 3924 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 2240 23032 2268 23063
rect 3786 23032 3792 23044
rect 2240 23004 3792 23032
rect 3786 22992 3792 23004
rect 3844 22992 3850 23044
rect 3896 23032 3924 23072
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4100 23103 4158 23109
rect 4100 23100 4112 23103
rect 4028 23072 4112 23100
rect 4028 23060 4034 23072
rect 4100 23069 4112 23072
rect 4146 23069 4158 23103
rect 4100 23063 4158 23069
rect 4203 23103 4261 23109
rect 4203 23069 4215 23103
rect 4249 23100 4261 23103
rect 4338 23100 4344 23112
rect 4249 23072 4344 23100
rect 4249 23069 4261 23072
rect 4203 23063 4261 23069
rect 4338 23060 4344 23072
rect 4396 23060 4402 23112
rect 7208 23086 7236 23140
rect 7834 23128 7840 23140
rect 7892 23168 7898 23180
rect 7944 23168 7972 23267
rect 9030 23264 9036 23276
rect 9088 23264 9094 23316
rect 14642 23264 14648 23316
rect 14700 23304 14706 23316
rect 16022 23304 16028 23316
rect 14700 23276 16028 23304
rect 14700 23264 14706 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 20438 23304 20444 23316
rect 20128 23276 20444 23304
rect 20128 23264 20134 23276
rect 20438 23264 20444 23276
rect 20496 23304 20502 23316
rect 21177 23307 21235 23313
rect 21177 23304 21189 23307
rect 20496 23276 21189 23304
rect 20496 23264 20502 23276
rect 21177 23273 21189 23276
rect 21223 23273 21235 23307
rect 21177 23267 21235 23273
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 21453 23307 21511 23313
rect 21453 23304 21465 23307
rect 21416 23276 21465 23304
rect 21416 23264 21422 23276
rect 21453 23273 21465 23276
rect 21499 23273 21511 23307
rect 21453 23267 21511 23273
rect 18233 23239 18291 23245
rect 18233 23205 18245 23239
rect 18279 23236 18291 23239
rect 19334 23236 19340 23248
rect 18279 23208 19340 23236
rect 18279 23205 18291 23208
rect 18233 23199 18291 23205
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 24670 23196 24676 23248
rect 24728 23236 24734 23248
rect 24728 23208 25176 23236
rect 24728 23196 24734 23208
rect 7892 23140 7972 23168
rect 11977 23171 12035 23177
rect 7892 23128 7898 23140
rect 11977 23137 11989 23171
rect 12023 23168 12035 23171
rect 12158 23168 12164 23180
rect 12023 23140 12164 23168
rect 12023 23137 12035 23140
rect 11977 23131 12035 23137
rect 12158 23128 12164 23140
rect 12216 23128 12222 23180
rect 12713 23171 12771 23177
rect 12713 23137 12725 23171
rect 12759 23168 12771 23171
rect 13538 23168 13544 23180
rect 12759 23140 13544 23168
rect 12759 23137 12771 23140
rect 12713 23131 12771 23137
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 14274 23128 14280 23180
rect 14332 23168 14338 23180
rect 15286 23168 15292 23180
rect 14332 23140 15292 23168
rect 14332 23128 14338 23140
rect 15286 23128 15292 23140
rect 15344 23168 15350 23180
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 15344 23140 16497 23168
rect 15344 23128 15350 23140
rect 16485 23137 16497 23140
rect 16531 23168 16543 23171
rect 18598 23168 18604 23180
rect 16531 23140 18604 23168
rect 16531 23137 16543 23140
rect 16485 23131 16543 23137
rect 18598 23128 18604 23140
rect 18656 23168 18662 23180
rect 25148 23177 25176 23208
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 18656 23140 19441 23168
rect 18656 23128 18662 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 25133 23171 25191 23177
rect 22051 23140 24992 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 9950 23060 9956 23112
rect 10008 23060 10014 23112
rect 10870 23060 10876 23112
rect 10928 23100 10934 23112
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 10928 23072 11713 23100
rect 10928 23060 10934 23072
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 12529 23103 12587 23109
rect 12529 23100 12541 23103
rect 11701 23063 11759 23069
rect 11808 23072 12541 23100
rect 5074 23032 5080 23044
rect 3896 23004 5080 23032
rect 5074 22992 5080 23004
rect 5132 22992 5138 23044
rect 6089 23035 6147 23041
rect 6089 23001 6101 23035
rect 6135 23001 6147 23035
rect 6089 22995 6147 23001
rect 3326 22924 3332 22976
rect 3384 22964 3390 22976
rect 5442 22964 5448 22976
rect 3384 22936 5448 22964
rect 3384 22924 3390 22936
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 6104 22964 6132 22995
rect 10686 22992 10692 23044
rect 10744 22992 10750 23044
rect 10778 22992 10784 23044
rect 10836 23032 10842 23044
rect 11808 23032 11836 23072
rect 12529 23069 12541 23072
rect 12575 23100 12587 23103
rect 13449 23103 13507 23109
rect 13449 23100 13461 23103
rect 12575 23072 13461 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 13449 23069 13461 23072
rect 13495 23069 13507 23103
rect 16390 23100 16396 23112
rect 15686 23072 16396 23100
rect 13449 23063 13507 23069
rect 16390 23060 16396 23072
rect 16448 23060 16454 23112
rect 22738 23060 22744 23112
rect 22796 23060 22802 23112
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24964 23109 24992 23140
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 10836 23004 11836 23032
rect 10836 22992 10842 23004
rect 12434 22992 12440 23044
rect 12492 23032 12498 23044
rect 13357 23035 13415 23041
rect 12492 23004 13032 23032
rect 12492 22992 12498 23004
rect 7466 22964 7472 22976
rect 6104 22936 7472 22964
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 9766 22924 9772 22976
rect 9824 22964 9830 22976
rect 11333 22967 11391 22973
rect 11333 22964 11345 22967
rect 9824 22936 11345 22964
rect 9824 22924 9830 22936
rect 11333 22933 11345 22936
rect 11379 22933 11391 22967
rect 11333 22927 11391 22933
rect 11698 22924 11704 22976
rect 11756 22964 11762 22976
rect 11793 22967 11851 22973
rect 11793 22964 11805 22967
rect 11756 22936 11805 22964
rect 11756 22924 11762 22936
rect 11793 22933 11805 22936
rect 11839 22964 11851 22967
rect 12250 22964 12256 22976
rect 11839 22936 12256 22964
rect 11839 22933 11851 22936
rect 11793 22927 11851 22933
rect 12250 22924 12256 22936
rect 12308 22924 12314 22976
rect 13004 22973 13032 23004
rect 13357 23001 13369 23035
rect 13403 23032 13415 23035
rect 13906 23032 13912 23044
rect 13403 23004 13912 23032
rect 13403 23001 13415 23004
rect 13357 22995 13415 23001
rect 13906 22992 13912 23004
rect 13964 22992 13970 23044
rect 14553 23035 14611 23041
rect 14553 23001 14565 23035
rect 14599 23001 14611 23035
rect 14553 22995 14611 23001
rect 12989 22967 13047 22973
rect 12989 22933 13001 22967
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 14568 22964 14596 22995
rect 15930 22992 15936 23044
rect 15988 23032 15994 23044
rect 16761 23035 16819 23041
rect 16761 23032 16773 23035
rect 15988 23004 16773 23032
rect 15988 22992 15994 23004
rect 16761 23001 16773 23004
rect 16807 23001 16819 23035
rect 17986 23004 18644 23032
rect 16761 22995 16819 23001
rect 16206 22964 16212 22976
rect 13136 22936 16212 22964
rect 13136 22924 13142 22936
rect 16206 22924 16212 22936
rect 16264 22924 16270 22976
rect 16390 22924 16396 22976
rect 16448 22964 16454 22976
rect 18064 22964 18092 23004
rect 18616 22973 18644 23004
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 19705 23035 19763 23041
rect 19705 23032 19717 23035
rect 19392 23004 19717 23032
rect 19392 22992 19398 23004
rect 19705 23001 19717 23004
rect 19751 23032 19763 23035
rect 19978 23032 19984 23044
rect 19751 23004 19984 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 21358 23032 21364 23044
rect 20930 23004 21364 23032
rect 16448 22936 18092 22964
rect 18601 22967 18659 22973
rect 16448 22924 16454 22936
rect 18601 22933 18613 22967
rect 18647 22964 18659 22967
rect 21008 22964 21036 23004
rect 21358 22992 21364 23004
rect 21416 22992 21422 23044
rect 23382 22992 23388 23044
rect 23440 23032 23446 23044
rect 25041 23035 25099 23041
rect 25041 23032 25053 23035
rect 23440 23004 25053 23032
rect 23440 22992 23446 23004
rect 25041 23001 25053 23004
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 18647 22936 21036 22964
rect 18647 22933 18659 22936
rect 18601 22927 18659 22933
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24581 22967 24639 22973
rect 24581 22964 24593 22967
rect 23532 22936 24593 22964
rect 23532 22924 23538 22936
rect 24581 22933 24593 22936
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 1762 22720 1768 22772
rect 1820 22760 1826 22772
rect 2041 22763 2099 22769
rect 2041 22760 2053 22763
rect 1820 22732 2053 22760
rect 1820 22720 1826 22732
rect 2041 22729 2053 22732
rect 2087 22729 2099 22763
rect 2041 22723 2099 22729
rect 5629 22763 5687 22769
rect 5629 22729 5641 22763
rect 5675 22760 5687 22763
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 5675 22732 6837 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 7193 22763 7251 22769
rect 7193 22729 7205 22763
rect 7239 22760 7251 22763
rect 8754 22760 8760 22772
rect 7239 22732 8760 22760
rect 7239 22729 7251 22732
rect 7193 22723 7251 22729
rect 8754 22720 8760 22732
rect 8812 22720 8818 22772
rect 9309 22763 9367 22769
rect 9309 22729 9321 22763
rect 9355 22760 9367 22763
rect 9950 22760 9956 22772
rect 9355 22732 9956 22760
rect 9355 22729 9367 22732
rect 9309 22723 9367 22729
rect 5902 22652 5908 22704
rect 5960 22692 5966 22704
rect 8021 22695 8079 22701
rect 5960 22664 7972 22692
rect 5960 22652 5966 22664
rect 2225 22627 2283 22633
rect 2225 22593 2237 22627
rect 2271 22624 2283 22627
rect 2866 22624 2872 22636
rect 2271 22596 2872 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22624 5779 22627
rect 6914 22624 6920 22636
rect 5767 22596 6920 22624
rect 5767 22593 5779 22596
rect 5721 22587 5779 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7558 22624 7564 22636
rect 7484 22596 7564 22624
rect 5905 22559 5963 22565
rect 5905 22525 5917 22559
rect 5951 22556 5963 22559
rect 5994 22556 6000 22568
rect 5951 22528 6000 22556
rect 5951 22525 5963 22528
rect 5905 22519 5963 22525
rect 5994 22516 6000 22528
rect 6052 22516 6058 22568
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 7484 22565 7512 22596
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 7944 22624 7972 22664
rect 8021 22661 8033 22695
rect 8067 22692 8079 22695
rect 9324 22692 9352 22723
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 10781 22763 10839 22769
rect 10781 22729 10793 22763
rect 10827 22760 10839 22763
rect 10827 22732 13308 22760
rect 10827 22729 10839 22732
rect 10781 22723 10839 22729
rect 8067 22664 9352 22692
rect 8067 22661 8079 22664
rect 8021 22655 8079 22661
rect 10042 22652 10048 22704
rect 10100 22692 10106 22704
rect 10137 22695 10195 22701
rect 10137 22692 10149 22695
rect 10100 22664 10149 22692
rect 10100 22652 10106 22664
rect 10137 22661 10149 22664
rect 10183 22692 10195 22695
rect 10873 22695 10931 22701
rect 10873 22692 10885 22695
rect 10183 22664 10885 22692
rect 10183 22661 10195 22664
rect 10137 22655 10195 22661
rect 10873 22661 10885 22664
rect 10919 22692 10931 22695
rect 12066 22692 12072 22704
rect 10919 22664 12072 22692
rect 10919 22661 10931 22664
rect 10873 22655 10931 22661
rect 12066 22652 12072 22664
rect 12124 22652 12130 22704
rect 13280 22701 13308 22732
rect 15194 22720 15200 22772
rect 15252 22720 15258 22772
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 15562 22760 15568 22772
rect 15344 22732 15568 22760
rect 15344 22720 15350 22732
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 16206 22720 16212 22772
rect 16264 22760 16270 22772
rect 16482 22760 16488 22772
rect 16264 22732 16488 22760
rect 16264 22720 16270 22732
rect 16482 22720 16488 22732
rect 16540 22720 16546 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 17494 22760 17500 22772
rect 16632 22732 17500 22760
rect 16632 22720 16638 22732
rect 17494 22720 17500 22732
rect 17552 22760 17558 22772
rect 20346 22760 20352 22772
rect 17552 22732 20352 22760
rect 17552 22720 17558 22732
rect 13265 22695 13323 22701
rect 13265 22661 13277 22695
rect 13311 22692 13323 22695
rect 15838 22692 15844 22704
rect 13311 22664 15844 22692
rect 13311 22661 13323 22664
rect 13265 22655 13323 22661
rect 15212 22636 15240 22664
rect 15838 22652 15844 22664
rect 15896 22652 15902 22704
rect 16390 22652 16396 22704
rect 16448 22652 16454 22704
rect 17880 22701 17908 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 23566 22720 23572 22772
rect 23624 22760 23630 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23624 22732 23765 22760
rect 23624 22720 23630 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 23753 22723 23811 22729
rect 24213 22763 24271 22769
rect 24213 22729 24225 22763
rect 24259 22760 24271 22763
rect 24305 22763 24363 22769
rect 24305 22760 24317 22763
rect 24259 22732 24317 22760
rect 24259 22729 24271 22732
rect 24213 22723 24271 22729
rect 24305 22729 24317 22732
rect 24351 22760 24363 22763
rect 24486 22760 24492 22772
rect 24351 22732 24492 22760
rect 24351 22729 24363 22732
rect 24305 22723 24363 22729
rect 17865 22695 17923 22701
rect 17865 22661 17877 22695
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 18598 22652 18604 22704
rect 18656 22652 18662 22704
rect 19702 22652 19708 22704
rect 19760 22652 19766 22704
rect 20364 22692 20392 22720
rect 20533 22695 20591 22701
rect 20533 22692 20545 22695
rect 20364 22664 20545 22692
rect 20533 22661 20545 22664
rect 20579 22661 20591 22695
rect 20533 22655 20591 22661
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 7944 22596 11621 22624
rect 11609 22593 11621 22596
rect 11655 22593 11667 22627
rect 11609 22587 11667 22593
rect 7469 22559 7527 22565
rect 7469 22525 7481 22559
rect 7515 22525 7527 22559
rect 7469 22519 7527 22525
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22556 11023 22559
rect 11146 22556 11152 22568
rect 11011 22528 11152 22556
rect 11011 22525 11023 22528
rect 10965 22519 11023 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 11624 22556 11652 22587
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 13078 22584 13084 22636
rect 13136 22584 13142 22636
rect 13814 22584 13820 22636
rect 13872 22624 13878 22636
rect 15105 22627 15163 22633
rect 15105 22624 15117 22627
rect 13872 22596 15117 22624
rect 13872 22584 13878 22596
rect 15105 22593 15117 22596
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 15194 22584 15200 22636
rect 15252 22584 15258 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19392 22596 19625 22624
rect 19392 22584 19398 22596
rect 19613 22593 19625 22596
rect 19659 22593 19671 22627
rect 19613 22587 19671 22593
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 22002 22624 22008 22636
rect 21407 22596 22008 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 23382 22584 23388 22636
rect 23440 22584 23446 22636
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 11624 22528 12449 22556
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13096 22556 13124 22584
rect 12667 22528 13124 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 6638 22488 6644 22500
rect 4488 22460 6644 22488
rect 4488 22448 4494 22460
rect 6638 22448 6644 22460
rect 6696 22448 6702 22500
rect 9398 22448 9404 22500
rect 9456 22488 9462 22500
rect 10413 22491 10471 22497
rect 10413 22488 10425 22491
rect 9456 22460 10425 22488
rect 9456 22448 9462 22460
rect 10413 22457 10425 22460
rect 10459 22457 10471 22491
rect 12452 22488 12480 22519
rect 13906 22516 13912 22568
rect 13964 22516 13970 22568
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 15930 22556 15936 22568
rect 15427 22528 15936 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 15930 22516 15936 22528
rect 15988 22516 15994 22568
rect 19794 22516 19800 22568
rect 19852 22516 19858 22568
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 21692 22528 22293 22556
rect 21692 22516 21698 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 23400 22556 23428 22584
rect 24228 22556 24256 22723
rect 24486 22720 24492 22732
rect 24544 22760 24550 22772
rect 24765 22763 24823 22769
rect 24765 22760 24777 22763
rect 24544 22732 24777 22760
rect 24544 22720 24550 22732
rect 24765 22729 24777 22732
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 25314 22720 25320 22772
rect 25372 22760 25378 22772
rect 25409 22763 25467 22769
rect 25409 22760 25421 22763
rect 25372 22732 25421 22760
rect 25372 22720 25378 22732
rect 25409 22729 25421 22732
rect 25455 22729 25467 22763
rect 25409 22723 25467 22729
rect 23400 22528 24256 22556
rect 22281 22519 22339 22525
rect 17862 22488 17868 22500
rect 12452 22460 17868 22488
rect 10413 22451 10471 22457
rect 17862 22448 17868 22460
rect 17920 22448 17926 22500
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 5261 22423 5319 22429
rect 5261 22420 5273 22423
rect 4304 22392 5273 22420
rect 4304 22380 4310 22392
rect 5261 22389 5273 22392
rect 5307 22389 5319 22423
rect 5261 22383 5319 22389
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 10502 22420 10508 22432
rect 7524 22392 10508 22420
rect 7524 22380 7530 22392
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 11977 22423 12035 22429
rect 11977 22389 11989 22423
rect 12023 22420 12035 22423
rect 12802 22420 12808 22432
rect 12023 22392 12808 22420
rect 12023 22389 12035 22392
rect 11977 22383 12035 22389
rect 12802 22380 12808 22392
rect 12860 22380 12866 22432
rect 14734 22380 14740 22432
rect 14792 22380 14798 22432
rect 19242 22380 19248 22432
rect 19300 22380 19306 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 13262 22176 13268 22228
rect 13320 22216 13326 22228
rect 13538 22216 13544 22228
rect 13320 22188 13544 22216
rect 13320 22176 13326 22188
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 16390 22176 16396 22228
rect 16448 22176 16454 22228
rect 19686 22219 19744 22225
rect 19686 22216 19698 22219
rect 18708 22188 19698 22216
rect 11422 22108 11428 22160
rect 11480 22108 11486 22160
rect 11790 22108 11796 22160
rect 11848 22148 11854 22160
rect 11848 22120 11928 22148
rect 11848 22108 11854 22120
rect 11900 22080 11928 22120
rect 12250 22108 12256 22160
rect 12308 22148 12314 22160
rect 18049 22151 18107 22157
rect 12308 22120 14412 22148
rect 12308 22108 12314 22120
rect 11977 22083 12035 22089
rect 11977 22080 11989 22083
rect 11900 22052 11989 22080
rect 11977 22049 11989 22052
rect 12023 22049 12035 22083
rect 11977 22043 12035 22049
rect 14274 22040 14280 22092
rect 14332 22040 14338 22092
rect 14384 22080 14412 22120
rect 18049 22117 18061 22151
rect 18095 22117 18107 22151
rect 18049 22111 18107 22117
rect 14550 22080 14556 22092
rect 14384 22052 14556 22080
rect 14550 22040 14556 22052
rect 14608 22080 14614 22092
rect 14918 22080 14924 22092
rect 14608 22052 14924 22080
rect 14608 22040 14614 22052
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 16022 22040 16028 22092
rect 16080 22040 16086 22092
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17497 22083 17555 22089
rect 16908 22052 17356 22080
rect 16908 22040 16914 22052
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 13265 22015 13323 22021
rect 11839 21984 12572 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 12544 21953 12572 21984
rect 13265 21981 13277 22015
rect 13311 22012 13323 22015
rect 13354 22012 13360 22024
rect 13311 21984 13360 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 16577 22015 16635 22021
rect 16577 21981 16589 22015
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 10888 21916 11897 21944
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 4522 21876 4528 21888
rect 4479 21848 4528 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 4522 21836 4528 21848
rect 4580 21836 4586 21888
rect 10594 21836 10600 21888
rect 10652 21876 10658 21888
rect 10888 21885 10916 21916
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 12529 21947 12587 21953
rect 12529 21913 12541 21947
rect 12575 21944 12587 21947
rect 12575 21916 14136 21944
rect 12575 21913 12587 21916
rect 12529 21907 12587 21913
rect 10873 21879 10931 21885
rect 10873 21876 10885 21879
rect 10652 21848 10885 21876
rect 10652 21836 10658 21848
rect 10873 21845 10885 21848
rect 10919 21845 10931 21879
rect 10873 21839 10931 21845
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11514 21876 11520 21888
rect 11204 21848 11520 21876
rect 11204 21836 11210 21848
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 12894 21836 12900 21888
rect 12952 21876 12958 21888
rect 13081 21879 13139 21885
rect 13081 21876 13093 21879
rect 12952 21848 13093 21876
rect 12952 21836 12958 21848
rect 13081 21845 13093 21848
rect 13127 21845 13139 21879
rect 14108 21876 14136 21916
rect 14182 21904 14188 21956
rect 14240 21944 14246 21956
rect 14553 21947 14611 21953
rect 14553 21944 14565 21947
rect 14240 21916 14565 21944
rect 14240 21904 14246 21916
rect 14553 21913 14565 21916
rect 14599 21944 14611 21947
rect 14642 21944 14648 21956
rect 14599 21916 14648 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 16390 21944 16396 21956
rect 15778 21916 16396 21944
rect 16390 21904 16396 21916
rect 16448 21904 16454 21956
rect 16592 21944 16620 21975
rect 17034 21972 17040 22024
rect 17092 22012 17098 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 17092 21984 17233 22012
rect 17092 21972 17098 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17328 21944 17356 22052
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17770 22080 17776 22092
rect 17543 22052 17776 22080
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 17770 22040 17776 22052
rect 17828 22040 17834 22092
rect 18064 22012 18092 22111
rect 18506 22040 18512 22092
rect 18564 22040 18570 22092
rect 18708 22089 18736 22188
rect 19686 22185 19698 22188
rect 19732 22216 19744 22219
rect 20254 22216 20260 22228
rect 19732 22188 20260 22216
rect 19732 22185 19744 22188
rect 19686 22179 19744 22185
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 21358 22176 21364 22228
rect 21416 22216 21422 22228
rect 21453 22219 21511 22225
rect 21453 22216 21465 22219
rect 21416 22188 21465 22216
rect 21416 22176 21422 22188
rect 21453 22185 21465 22188
rect 21499 22185 21511 22219
rect 21453 22179 21511 22185
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22049 18751 22083
rect 18693 22043 18751 22049
rect 19334 22040 19340 22092
rect 19392 22040 19398 22092
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 22002 22080 22008 22092
rect 19852 22052 22008 22080
rect 19852 22040 19858 22052
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 24029 22083 24087 22089
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 24302 22080 24308 22092
rect 24075 22052 24308 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 19352 22012 19380 22040
rect 18064 21984 19380 22012
rect 19429 22015 19487 22021
rect 19429 21981 19441 22015
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 18417 21947 18475 21953
rect 18417 21944 18429 21947
rect 16592 21916 16988 21944
rect 17328 21916 18429 21944
rect 15470 21876 15476 21888
rect 14108 21848 15476 21876
rect 13081 21839 13139 21845
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 16960 21876 16988 21916
rect 18417 21913 18429 21916
rect 18463 21913 18475 21947
rect 19444 21944 19472 21975
rect 23382 21972 23388 22024
rect 23440 21972 23446 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24176 21984 24869 22012
rect 24176 21972 24182 21984
rect 24857 21981 24869 21984
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 19794 21944 19800 21956
rect 19444 21916 19800 21944
rect 18417 21907 18475 21913
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 21450 21944 21456 21956
rect 20930 21916 21456 21944
rect 21450 21904 21456 21916
rect 21508 21904 21514 21956
rect 22278 21904 22284 21956
rect 22336 21904 22342 21956
rect 24673 21947 24731 21953
rect 24673 21913 24685 21947
rect 24719 21913 24731 21947
rect 24673 21907 24731 21913
rect 17313 21879 17371 21885
rect 17313 21876 17325 21879
rect 16960 21848 17325 21876
rect 17313 21845 17325 21848
rect 17359 21876 17371 21879
rect 19518 21876 19524 21888
rect 17359 21848 19524 21876
rect 17359 21845 17371 21848
rect 17313 21839 17371 21845
rect 19518 21836 19524 21848
rect 19576 21836 19582 21888
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 21177 21879 21235 21885
rect 21177 21876 21189 21879
rect 19944 21848 21189 21876
rect 19944 21836 19950 21848
rect 21177 21845 21189 21848
rect 21223 21845 21235 21879
rect 21177 21839 21235 21845
rect 21266 21836 21272 21888
rect 21324 21876 21330 21888
rect 24688 21876 24716 21907
rect 21324 21848 24716 21876
rect 21324 21836 21330 21848
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 7098 21632 7104 21684
rect 7156 21632 7162 21684
rect 7469 21675 7527 21681
rect 7469 21641 7481 21675
rect 7515 21672 7527 21675
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 7515 21644 8309 21672
rect 7515 21641 7527 21644
rect 7469 21635 7527 21641
rect 8297 21641 8309 21644
rect 8343 21641 8355 21675
rect 8297 21635 8355 21641
rect 8665 21675 8723 21681
rect 8665 21641 8677 21675
rect 8711 21672 8723 21675
rect 9766 21672 9772 21684
rect 8711 21644 9772 21672
rect 8711 21641 8723 21644
rect 8665 21635 8723 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 9907 21644 11713 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12069 21675 12127 21681
rect 12069 21672 12081 21675
rect 12032 21644 12081 21672
rect 12032 21632 12038 21644
rect 12069 21641 12081 21644
rect 12115 21641 12127 21675
rect 12069 21635 12127 21641
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13814 21672 13820 21684
rect 13587 21644 13820 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 17218 21672 17224 21684
rect 15436 21644 17224 21672
rect 15436 21632 15442 21644
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 18509 21675 18567 21681
rect 18509 21641 18521 21675
rect 18555 21641 18567 21675
rect 18509 21635 18567 21641
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 7708 21576 10088 21604
rect 7708 21564 7714 21576
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 1854 21536 1860 21548
rect 1811 21508 1860 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 1854 21496 1860 21508
rect 1912 21496 1918 21548
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21536 3479 21539
rect 4154 21536 4160 21548
rect 3467 21508 4160 21536
rect 3467 21505 3479 21508
rect 3421 21499 3479 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4522 21496 4528 21548
rect 4580 21496 4586 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 8938 21536 8944 21548
rect 7607 21508 8944 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 1302 21428 1308 21480
rect 1360 21468 1366 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 1360 21440 2053 21468
rect 1360 21428 1366 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 4062 21468 4068 21480
rect 3660 21440 4068 21468
rect 3660 21428 3666 21440
rect 4062 21428 4068 21440
rect 4120 21468 4126 21480
rect 4985 21471 5043 21477
rect 4985 21468 4997 21471
rect 4120 21440 4997 21468
rect 4120 21428 4126 21440
rect 4985 21437 4997 21440
rect 5031 21437 5043 21471
rect 4985 21431 5043 21437
rect 7650 21428 7656 21480
rect 7708 21428 7714 21480
rect 8754 21428 8760 21480
rect 8812 21428 8818 21480
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21468 8907 21471
rect 9030 21468 9036 21480
rect 8895 21440 9036 21468
rect 8895 21437 8907 21440
rect 8849 21431 8907 21437
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 10060 21477 10088 21576
rect 12802 21564 12808 21616
rect 12860 21604 12866 21616
rect 14001 21607 14059 21613
rect 14001 21604 14013 21607
rect 12860 21576 14013 21604
rect 12860 21564 12866 21576
rect 14001 21573 14013 21576
rect 14047 21573 14059 21607
rect 18524 21604 18552 21635
rect 18690 21632 18696 21684
rect 18748 21672 18754 21684
rect 21266 21672 21272 21684
rect 18748 21644 21272 21672
rect 18748 21632 18754 21644
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 22554 21632 22560 21684
rect 22612 21632 22618 21684
rect 23382 21632 23388 21684
rect 23440 21672 23446 21684
rect 23566 21672 23572 21684
rect 23440 21644 23572 21672
rect 23440 21632 23446 21644
rect 23566 21632 23572 21644
rect 23624 21672 23630 21684
rect 25409 21675 25467 21681
rect 25409 21672 25421 21675
rect 23624 21644 23796 21672
rect 23624 21632 23630 21644
rect 21082 21604 21088 21616
rect 14001 21567 14059 21573
rect 14108 21576 17080 21604
rect 18524 21576 21088 21604
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21536 12219 21539
rect 13906 21536 13912 21548
rect 12207 21508 13912 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 10045 21471 10103 21477
rect 10045 21437 10057 21471
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 3786 21360 3792 21412
rect 3844 21360 3850 21412
rect 6914 21360 6920 21412
rect 6972 21400 6978 21412
rect 9493 21403 9551 21409
rect 9493 21400 9505 21403
rect 6972 21372 9505 21400
rect 6972 21360 6978 21372
rect 9493 21369 9505 21372
rect 9539 21369 9551 21403
rect 9968 21400 9996 21431
rect 11054 21428 11060 21480
rect 11112 21468 11118 21480
rect 12342 21468 12348 21480
rect 11112 21440 12348 21468
rect 11112 21428 11118 21440
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 14108 21468 14136 21576
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21536 15255 21539
rect 16114 21536 16120 21548
rect 15243 21508 16120 21536
rect 15243 21505 15255 21508
rect 15197 21499 15255 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 17052 21545 17080 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 22002 21564 22008 21616
rect 22060 21604 22066 21616
rect 22060 21576 23428 21604
rect 22060 21564 22066 21576
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21505 16267 21539
rect 16209 21499 16267 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 13780 21440 14136 21468
rect 13780 21428 13786 21440
rect 14182 21428 14188 21480
rect 14240 21428 14246 21480
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 15289 21471 15347 21477
rect 15289 21468 15301 21471
rect 14700 21440 15301 21468
rect 14700 21428 14706 21440
rect 15289 21437 15301 21440
rect 15335 21437 15347 21471
rect 15289 21431 15347 21437
rect 15378 21428 15384 21480
rect 15436 21428 15442 21480
rect 10778 21400 10784 21412
rect 9968 21372 10784 21400
rect 9493 21363 9551 21369
rect 10778 21360 10784 21372
rect 10836 21360 10842 21412
rect 4801 21335 4859 21341
rect 4801 21301 4813 21335
rect 4847 21332 4859 21335
rect 5810 21332 5816 21344
rect 4847 21304 5816 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 7558 21292 7564 21344
rect 7616 21332 7622 21344
rect 8202 21332 8208 21344
rect 7616 21304 8208 21332
rect 7616 21292 7622 21304
rect 8202 21292 8208 21304
rect 8260 21332 8266 21344
rect 11072 21332 11100 21428
rect 11330 21360 11336 21412
rect 11388 21400 11394 21412
rect 16224 21400 16252 21499
rect 17402 21496 17408 21548
rect 17460 21536 17466 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 17460 21508 18705 21536
rect 17460 21496 17466 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 23290 21536 23296 21548
rect 22511 21508 23296 21536
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 23400 21545 23428 21576
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 23768 21604 23796 21644
rect 24044 21644 25421 21672
rect 24044 21604 24072 21644
rect 25409 21641 25421 21644
rect 25455 21641 25467 21675
rect 25409 21635 25467 21641
rect 23768 21576 24150 21604
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 17681 21471 17739 21477
rect 17681 21468 17693 21471
rect 17644 21440 17693 21468
rect 17644 21428 17650 21440
rect 17681 21437 17693 21440
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 20622 21468 20628 21480
rect 19576 21440 20628 21468
rect 19576 21428 19582 21440
rect 20622 21428 20628 21440
rect 20680 21468 20686 21480
rect 20990 21468 20996 21480
rect 20680 21440 20996 21468
rect 20680 21428 20686 21440
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 22278 21428 22284 21480
rect 22336 21468 22342 21480
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22336 21440 22753 21468
rect 22336 21428 22342 21440
rect 22741 21437 22753 21440
rect 22787 21468 22799 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 22787 21440 25145 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 11388 21372 16252 21400
rect 16853 21403 16911 21409
rect 11388 21360 11394 21372
rect 16853 21369 16865 21403
rect 16899 21400 16911 21403
rect 22462 21400 22468 21412
rect 16899 21372 22468 21400
rect 16899 21369 16911 21372
rect 16853 21363 16911 21369
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 8260 21304 11100 21332
rect 8260 21292 8266 21304
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 13872 21304 14841 21332
rect 13872 21292 13878 21304
rect 14829 21301 14841 21304
rect 14875 21301 14887 21335
rect 14829 21295 14887 21301
rect 16022 21292 16028 21344
rect 16080 21292 16086 21344
rect 16390 21292 16396 21344
rect 16448 21332 16454 21344
rect 19518 21332 19524 21344
rect 16448 21304 19524 21332
rect 16448 21292 16454 21304
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 20438 21292 20444 21344
rect 20496 21292 20502 21344
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 20864 21304 22109 21332
rect 20864 21292 20870 21304
rect 22097 21301 22109 21304
rect 22143 21301 22155 21335
rect 22097 21295 22155 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 2866 21088 2872 21140
rect 2924 21128 2930 21140
rect 3145 21131 3203 21137
rect 3145 21128 3157 21131
rect 2924 21100 3157 21128
rect 2924 21088 2930 21100
rect 3145 21097 3157 21100
rect 3191 21097 3203 21131
rect 3145 21091 3203 21097
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7837 21131 7895 21137
rect 7837 21128 7849 21131
rect 7340 21100 7849 21128
rect 7340 21088 7346 21100
rect 7837 21097 7849 21100
rect 7883 21097 7895 21131
rect 7837 21091 7895 21097
rect 9122 21088 9128 21140
rect 9180 21128 9186 21140
rect 10042 21128 10048 21140
rect 9180 21100 10048 21128
rect 9180 21088 9186 21100
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 16040 21100 16313 21128
rect 4065 21063 4123 21069
rect 4065 21029 4077 21063
rect 4111 21029 4123 21063
rect 4065 21023 4123 21029
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 4080 20992 4108 21023
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 14369 21063 14427 21069
rect 14369 21060 14381 21063
rect 12308 21032 14381 21060
rect 12308 21020 12314 21032
rect 14369 21029 14381 21032
rect 14415 21029 14427 21063
rect 14369 21023 14427 21029
rect 2823 20964 4108 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 8389 20995 8447 21001
rect 8389 20992 8401 20995
rect 8260 20964 8401 20992
rect 8260 20952 8266 20964
rect 8389 20961 8401 20964
rect 8435 20961 8447 20995
rect 8389 20955 8447 20961
rect 9769 20995 9827 21001
rect 9769 20961 9781 20995
rect 9815 20992 9827 20995
rect 10686 20992 10692 21004
rect 9815 20964 10692 20992
rect 9815 20961 9827 20964
rect 9769 20955 9827 20961
rect 10686 20952 10692 20964
rect 10744 20952 10750 21004
rect 11238 20952 11244 21004
rect 11296 20952 11302 21004
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 11974 20992 11980 21004
rect 11572 20964 11980 20992
rect 11572 20952 11578 20964
rect 11974 20952 11980 20964
rect 12032 20992 12038 21004
rect 13817 20995 13875 21001
rect 13817 20992 13829 20995
rect 12032 20964 13829 20992
rect 12032 20952 12038 20964
rect 13817 20961 13829 20964
rect 13863 20992 13875 20995
rect 14921 20995 14979 21001
rect 14921 20992 14933 20995
rect 13863 20964 14933 20992
rect 13863 20961 13875 20964
rect 13817 20955 13875 20961
rect 14921 20961 14933 20964
rect 14967 20961 14979 20995
rect 14921 20955 14979 20961
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20893 2283 20927
rect 2225 20887 2283 20893
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 4062 20924 4068 20936
rect 3007 20896 4068 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 2240 20856 2268 20887
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 11256 20924 11284 20952
rect 11885 20927 11943 20933
rect 11885 20924 11897 20927
rect 11178 20896 11897 20924
rect 11885 20893 11897 20896
rect 11931 20893 11943 20927
rect 13725 20927 13783 20933
rect 13725 20924 13737 20927
rect 11885 20887 11943 20893
rect 12406 20896 13737 20924
rect 8478 20856 8484 20868
rect 2240 20828 2774 20856
rect 2746 20800 2774 20828
rect 8220 20828 8484 20856
rect 1762 20748 1768 20800
rect 1820 20788 1826 20800
rect 2041 20791 2099 20797
rect 2041 20788 2053 20791
rect 1820 20760 2053 20788
rect 1820 20748 1826 20760
rect 2041 20757 2053 20760
rect 2087 20757 2099 20791
rect 2746 20760 2780 20800
rect 2041 20751 2099 20757
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 4706 20748 4712 20800
rect 4764 20788 4770 20800
rect 8220 20797 8248 20828
rect 8478 20816 8484 20828
rect 8536 20816 8542 20868
rect 10042 20816 10048 20868
rect 10100 20816 10106 20868
rect 12406 20856 12434 20896
rect 13725 20893 13737 20896
rect 13771 20924 13783 20927
rect 14829 20927 14887 20933
rect 14829 20924 14841 20927
rect 13771 20896 14841 20924
rect 13771 20893 13783 20896
rect 13725 20887 13783 20893
rect 14829 20893 14841 20896
rect 14875 20924 14887 20927
rect 15010 20924 15016 20936
rect 14875 20896 15016 20924
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 15010 20884 15016 20896
rect 15068 20884 15074 20936
rect 15746 20884 15752 20936
rect 15804 20884 15810 20936
rect 11348 20828 12434 20856
rect 14737 20859 14795 20865
rect 7469 20791 7527 20797
rect 7469 20788 7481 20791
rect 4764 20760 7481 20788
rect 4764 20748 4770 20760
rect 7469 20757 7481 20760
rect 7515 20788 7527 20791
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7515 20760 8217 20788
rect 7515 20757 7527 20760
rect 7469 20751 7527 20757
rect 8205 20757 8217 20760
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8297 20791 8355 20797
rect 8297 20757 8309 20791
rect 8343 20788 8355 20791
rect 10410 20788 10416 20800
rect 8343 20760 10416 20788
rect 8343 20757 8355 20760
rect 8297 20751 8355 20757
rect 10410 20748 10416 20760
rect 10468 20748 10474 20800
rect 10686 20748 10692 20800
rect 10744 20788 10750 20800
rect 11348 20788 11376 20828
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 16040 20856 16068 21100
rect 16301 21097 16313 21100
rect 16347 21128 16359 21131
rect 16390 21128 16396 21140
rect 16347 21100 16396 21128
rect 16347 21097 16359 21100
rect 16301 21091 16359 21097
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 17126 21128 17132 21140
rect 16991 21100 17132 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 20162 21128 20168 21140
rect 17788 21100 20168 21128
rect 16114 21020 16120 21072
rect 16172 21060 16178 21072
rect 17788 21060 17816 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 21450 21088 21456 21140
rect 21508 21128 21514 21140
rect 21913 21131 21971 21137
rect 21913 21128 21925 21131
rect 21508 21100 21925 21128
rect 21508 21088 21514 21100
rect 21913 21097 21925 21100
rect 21959 21097 21971 21131
rect 21913 21091 21971 21097
rect 16172 21032 17816 21060
rect 17880 21032 20024 21060
rect 16172 21020 16178 21032
rect 17126 20952 17132 21004
rect 17184 20992 17190 21004
rect 17880 21001 17908 21032
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 17184 20964 17693 20992
rect 17184 20952 17190 20964
rect 17681 20961 17693 20964
rect 17727 20961 17739 20995
rect 17681 20955 17739 20961
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20961 17923 20995
rect 17865 20955 17923 20961
rect 19794 20952 19800 21004
rect 19852 20992 19858 21004
rect 19889 20995 19947 21001
rect 19889 20992 19901 20995
rect 19852 20964 19901 20992
rect 19852 20952 19858 20964
rect 19889 20961 19901 20964
rect 19935 20961 19947 20995
rect 19996 20992 20024 21032
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 19996 20964 20177 20992
rect 19889 20955 19947 20961
rect 20165 20961 20177 20964
rect 20211 20992 20223 20995
rect 20530 20992 20536 21004
rect 20211 20964 20536 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 20530 20952 20536 20964
rect 20588 20952 20594 21004
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 17586 20884 17592 20936
rect 17644 20884 17650 20936
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 21450 20924 21456 20936
rect 21298 20896 21456 20924
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 25406 20924 25412 20936
rect 22879 20896 25412 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 19426 20856 19432 20868
rect 14783 20828 16068 20856
rect 17236 20828 19432 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 10744 20760 11376 20788
rect 11517 20791 11575 20797
rect 10744 20748 10750 20760
rect 11517 20757 11529 20791
rect 11563 20788 11575 20791
rect 12342 20788 12348 20800
rect 11563 20760 12348 20788
rect 11563 20757 11575 20760
rect 11517 20751 11575 20757
rect 12342 20748 12348 20760
rect 12400 20748 12406 20800
rect 15562 20748 15568 20800
rect 15620 20748 15626 20800
rect 17236 20797 17264 20828
rect 19426 20816 19432 20828
rect 19484 20816 19490 20868
rect 24854 20856 24860 20868
rect 21468 20828 24860 20856
rect 17221 20791 17279 20797
rect 17221 20757 17233 20791
rect 17267 20757 17279 20791
rect 17221 20751 17279 20757
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 21468 20788 21496 20828
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 18739 20760 21496 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 8846 20584 8852 20596
rect 6604 20556 8852 20584
rect 6604 20544 6610 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 8996 20556 9965 20584
rect 8996 20544 9002 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 9953 20547 10011 20553
rect 17310 20544 17316 20596
rect 17368 20584 17374 20596
rect 17368 20556 17724 20584
rect 17368 20544 17374 20556
rect 4249 20519 4307 20525
rect 4249 20485 4261 20519
rect 4295 20516 4307 20519
rect 4338 20516 4344 20528
rect 4295 20488 4344 20516
rect 4295 20485 4307 20488
rect 4249 20479 4307 20485
rect 4338 20476 4344 20488
rect 4396 20476 4402 20528
rect 5997 20519 6055 20525
rect 5997 20516 6009 20519
rect 5474 20488 6009 20516
rect 5997 20485 6009 20488
rect 6043 20516 6055 20519
rect 7098 20516 7104 20528
rect 6043 20488 7104 20516
rect 6043 20485 6055 20488
rect 5997 20479 6055 20485
rect 7098 20476 7104 20488
rect 7156 20516 7162 20528
rect 7156 20488 7314 20516
rect 7156 20476 7162 20488
rect 9030 20476 9036 20528
rect 9088 20516 9094 20528
rect 10413 20519 10471 20525
rect 9088 20488 9444 20516
rect 9088 20476 9094 20488
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 3988 20380 4016 20411
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 9125 20451 9183 20457
rect 9125 20448 9137 20451
rect 8720 20420 9137 20448
rect 8720 20408 8726 20420
rect 9125 20417 9137 20420
rect 9171 20417 9183 20451
rect 9125 20411 9183 20417
rect 5718 20380 5724 20392
rect 3988 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6871 20352 9168 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 8754 20272 8760 20324
rect 8812 20272 8818 20324
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 5810 20244 5816 20256
rect 5767 20216 5816 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9030 20244 9036 20256
rect 8352 20216 9036 20244
rect 8352 20204 8358 20216
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 9140 20244 9168 20352
rect 9214 20340 9220 20392
rect 9272 20340 9278 20392
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20349 9367 20383
rect 9416 20380 9444 20488
rect 10413 20485 10425 20519
rect 10459 20516 10471 20519
rect 11514 20516 11520 20528
rect 10459 20488 11520 20516
rect 10459 20485 10471 20488
rect 10413 20479 10471 20485
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 12526 20516 12532 20528
rect 11848 20488 12532 20516
rect 11848 20476 11854 20488
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 14274 20516 14280 20528
rect 13964 20488 14280 20516
rect 13964 20476 13970 20488
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 17696 20525 17724 20556
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 19392 20556 19441 20584
rect 19392 20544 19398 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 23293 20519 23351 20525
rect 23293 20485 23305 20519
rect 23339 20516 23351 20519
rect 23382 20516 23388 20528
rect 23339 20488 23388 20516
rect 23339 20485 23351 20488
rect 23293 20479 23351 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 11698 20448 11704 20460
rect 10367 20420 11704 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20448 12495 20451
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12483 20420 13277 20448
rect 12483 20417 12495 20420
rect 12437 20411 12495 20417
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 13688 20420 15669 20448
rect 13688 20408 13694 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20448 19395 20451
rect 19426 20448 19432 20460
rect 19383 20420 19432 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 24026 20448 24032 20460
rect 22327 20420 24032 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 24026 20408 24032 20420
rect 24084 20408 24090 20460
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24210 20448 24216 20460
rect 24167 20420 24216 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 10505 20383 10563 20389
rect 10505 20380 10517 20383
rect 9416 20352 10517 20380
rect 9309 20343 9367 20349
rect 10505 20349 10517 20352
rect 10551 20349 10563 20383
rect 10505 20343 10563 20349
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 9324 20244 9352 20343
rect 12158 20312 12164 20324
rect 11716 20284 12164 20312
rect 11716 20244 11744 20284
rect 12158 20272 12164 20284
rect 12216 20272 12222 20324
rect 9140 20216 11744 20244
rect 12066 20204 12072 20256
rect 12124 20204 12130 20256
rect 12544 20244 12572 20343
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 19613 20383 19671 20389
rect 19613 20349 19625 20383
rect 19659 20380 19671 20383
rect 21634 20380 21640 20392
rect 19659 20352 21640 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23348 20352 24409 20380
rect 23348 20340 23354 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 13906 20272 13912 20324
rect 13964 20312 13970 20324
rect 14642 20312 14648 20324
rect 13964 20284 14648 20312
rect 13964 20272 13970 20284
rect 14642 20272 14648 20284
rect 14700 20272 14706 20324
rect 15473 20315 15531 20321
rect 15473 20281 15485 20315
rect 15519 20312 15531 20315
rect 20990 20312 20996 20324
rect 15519 20284 20996 20312
rect 15519 20281 15531 20284
rect 15473 20275 15531 20281
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 13630 20244 13636 20256
rect 12544 20216 13636 20244
rect 13630 20204 13636 20216
rect 13688 20244 13694 20256
rect 13725 20247 13783 20253
rect 13725 20244 13737 20247
rect 13688 20216 13737 20244
rect 13688 20204 13694 20216
rect 13725 20213 13737 20216
rect 13771 20244 13783 20247
rect 13998 20244 14004 20256
rect 13771 20216 14004 20244
rect 13771 20213 13783 20216
rect 13725 20207 13783 20213
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 17770 20204 17776 20256
rect 17828 20204 17834 20256
rect 18325 20247 18383 20253
rect 18325 20213 18337 20247
rect 18371 20244 18383 20247
rect 18782 20244 18788 20256
rect 18371 20216 18788 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 18969 20247 19027 20253
rect 18969 20213 18981 20247
rect 19015 20244 19027 20247
rect 19794 20244 19800 20256
rect 19015 20216 19800 20244
rect 19015 20213 19027 20216
rect 18969 20207 19027 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 5074 20000 5080 20052
rect 5132 20000 5138 20052
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 6546 20040 6552 20052
rect 5776 20012 6552 20040
rect 5776 20000 5782 20012
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 11698 20000 11704 20052
rect 11756 20000 11762 20052
rect 14274 20000 14280 20052
rect 14332 20000 14338 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19150 20040 19156 20052
rect 18932 20012 19156 20040
rect 18932 20000 18938 20012
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 20254 20000 20260 20052
rect 20312 20000 20318 20052
rect 5736 19913 5764 20000
rect 15381 19975 15439 19981
rect 15381 19941 15393 19975
rect 15427 19972 15439 19975
rect 18322 19972 18328 19984
rect 15427 19944 18328 19972
rect 15427 19941 15439 19944
rect 15381 19935 15439 19941
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19904 6055 19907
rect 8294 19904 8300 19916
rect 6043 19876 8300 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8846 19864 8852 19916
rect 8904 19904 8910 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 8904 19876 9137 19904
rect 8904 19864 8910 19876
rect 9125 19873 9137 19876
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 11149 19907 11207 19913
rect 11149 19873 11161 19907
rect 11195 19904 11207 19907
rect 11790 19904 11796 19916
rect 11195 19876 11796 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 12158 19904 12164 19916
rect 11900 19876 12164 19904
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5276 19700 5304 19799
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7745 19839 7803 19845
rect 7745 19836 7757 19839
rect 7156 19808 7757 19836
rect 7156 19796 7162 19808
rect 7745 19805 7757 19808
rect 7791 19836 7803 19839
rect 7834 19836 7840 19848
rect 7791 19808 7840 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 7834 19796 7840 19808
rect 7892 19836 7898 19848
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 7892 19808 8401 19836
rect 7892 19796 7898 19808
rect 8389 19805 8401 19808
rect 8435 19836 8447 19839
rect 8938 19836 8944 19848
rect 8435 19808 8944 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11900 19836 11928 19876
rect 12158 19864 12164 19876
rect 12216 19904 12222 19916
rect 12253 19907 12311 19913
rect 12253 19904 12265 19907
rect 12216 19876 12265 19904
rect 12216 19864 12222 19876
rect 12253 19873 12265 19876
rect 12299 19873 12311 19907
rect 12253 19867 12311 19873
rect 13906 19864 13912 19916
rect 13964 19904 13970 19916
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13964 19876 14841 19904
rect 13964 19864 13970 19876
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 11756 19808 11928 19836
rect 12069 19839 12127 19845
rect 11756 19796 11762 19808
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12434 19836 12440 19848
rect 12115 19808 12440 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 15396 19836 15424 19935
rect 18322 19932 18328 19944
rect 18380 19972 18386 19984
rect 19978 19972 19984 19984
rect 18380 19944 19984 19972
rect 18380 19932 18386 19944
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 19150 19904 19156 19916
rect 16080 19876 19156 19904
rect 16080 19864 16086 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19904 23903 19907
rect 24946 19904 24952 19916
rect 23891 19876 24952 19904
rect 23891 19873 23903 19876
rect 23845 19867 23903 19873
rect 24946 19864 24952 19876
rect 25004 19864 25010 19916
rect 14691 19808 15424 19836
rect 17221 19839 17279 19845
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17267 19808 17785 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17773 19805 17785 19808
rect 17819 19836 17831 19839
rect 17862 19836 17868 19848
rect 17819 19808 17868 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18966 19836 18972 19848
rect 18739 19808 18972 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 22005 19839 22063 19845
rect 22005 19836 22017 19839
rect 20772 19808 22017 19836
rect 20772 19796 20778 19808
rect 22005 19805 22017 19808
rect 22051 19805 22063 19839
rect 22005 19799 22063 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 25038 19836 25044 19848
rect 22879 19808 25044 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 25038 19796 25044 19808
rect 25096 19796 25102 19848
rect 7650 19768 7656 19780
rect 7484 19740 7656 19768
rect 7374 19700 7380 19712
rect 5276 19672 7380 19700
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 7484 19709 7512 19740
rect 7650 19728 7656 19740
rect 7708 19768 7714 19780
rect 9401 19771 9459 19777
rect 9401 19768 9413 19771
rect 7708 19740 9413 19768
rect 7708 19728 7714 19740
rect 9401 19737 9413 19740
rect 9447 19737 9459 19771
rect 9401 19731 9459 19737
rect 9508 19740 9890 19768
rect 7469 19703 7527 19709
rect 7469 19669 7481 19703
rect 7515 19669 7527 19703
rect 7469 19663 7527 19669
rect 8662 19660 8668 19712
rect 8720 19660 8726 19712
rect 8938 19660 8944 19712
rect 8996 19700 9002 19712
rect 9508 19700 9536 19740
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 11974 19768 11980 19780
rect 11848 19740 11980 19768
rect 11848 19728 11854 19740
rect 11974 19728 11980 19740
rect 12032 19728 12038 19780
rect 12161 19771 12219 19777
rect 12161 19737 12173 19771
rect 12207 19768 12219 19771
rect 14182 19768 14188 19780
rect 12207 19740 14188 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 14568 19740 17325 19768
rect 8996 19672 9536 19700
rect 8996 19660 9002 19672
rect 10962 19660 10968 19712
rect 11020 19700 11026 19712
rect 13722 19700 13728 19712
rect 11020 19672 13728 19700
rect 11020 19660 11026 19672
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 14568 19700 14596 19740
rect 14752 19709 14780 19740
rect 17313 19737 17325 19740
rect 17359 19768 17371 19771
rect 17586 19768 17592 19780
rect 17359 19740 17592 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17957 19771 18015 19777
rect 17957 19737 17969 19771
rect 18003 19768 18015 19771
rect 18598 19768 18604 19780
rect 18003 19740 18604 19768
rect 18003 19737 18015 19740
rect 17957 19731 18015 19737
rect 18598 19728 18604 19740
rect 18656 19728 18662 19780
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19768 22247 19771
rect 23658 19768 23664 19780
rect 22235 19740 23664 19768
rect 22235 19737 22247 19740
rect 22189 19731 22247 19737
rect 23658 19728 23664 19740
rect 23716 19728 23722 19780
rect 13955 19672 14596 19700
rect 14737 19703 14795 19709
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 14737 19669 14749 19703
rect 14783 19700 14795 19703
rect 14826 19700 14832 19712
rect 14783 19672 14832 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 18966 19700 18972 19712
rect 18555 19672 18972 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 19337 19703 19395 19709
rect 19337 19669 19349 19703
rect 19383 19700 19395 19703
rect 19518 19700 19524 19712
rect 19383 19672 19524 19700
rect 19383 19669 19395 19672
rect 19337 19663 19395 19669
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 1544 19468 2053 19496
rect 1544 19456 1550 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2041 19459 2099 19465
rect 4154 19456 4160 19508
rect 4212 19496 4218 19508
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 4212 19468 4261 19496
rect 4212 19456 4218 19468
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8757 19499 8815 19505
rect 8757 19496 8769 19499
rect 7892 19468 8769 19496
rect 7892 19456 7898 19468
rect 8757 19465 8769 19468
rect 8803 19465 8815 19499
rect 8757 19459 8815 19465
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19496 9275 19499
rect 9398 19496 9404 19508
rect 9263 19468 9404 19496
rect 9263 19465 9275 19468
rect 9217 19459 9275 19465
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 11701 19499 11759 19505
rect 11701 19465 11713 19499
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 12069 19499 12127 19505
rect 12069 19465 12081 19499
rect 12115 19496 12127 19499
rect 12802 19496 12808 19508
rect 12115 19468 12808 19496
rect 12115 19465 12127 19468
rect 12069 19459 12127 19465
rect 7098 19388 7104 19440
rect 7156 19428 7162 19440
rect 7156 19400 7314 19428
rect 7156 19388 7162 19400
rect 9306 19388 9312 19440
rect 9364 19428 9370 19440
rect 11716 19428 11744 19459
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19496 13323 19499
rect 14001 19499 14059 19505
rect 14001 19496 14013 19499
rect 13311 19468 14013 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 14001 19465 14013 19468
rect 14047 19496 14059 19499
rect 14090 19496 14096 19508
rect 14047 19468 14096 19496
rect 14047 19465 14059 19468
rect 14001 19459 14059 19465
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 17310 19496 17316 19508
rect 16899 19468 17316 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 19889 19499 19947 19505
rect 17543 19468 19840 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 9364 19400 11744 19428
rect 9364 19388 9370 19400
rect 13722 19388 13728 19440
rect 13780 19428 13786 19440
rect 13780 19400 17080 19428
rect 13780 19388 13786 19400
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 3602 19360 3608 19372
rect 2271 19332 3608 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19360 4491 19363
rect 6270 19360 6276 19372
rect 4479 19332 6276 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8386 19320 8392 19372
rect 8444 19360 8450 19372
rect 8846 19360 8852 19372
rect 8444 19332 8852 19360
rect 8444 19320 8450 19332
rect 8846 19320 8852 19332
rect 8904 19360 8910 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 8904 19332 9137 19360
rect 8904 19320 8910 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 11974 19360 11980 19372
rect 9125 19323 9183 19329
rect 11072 19332 11980 19360
rect 6822 19252 6828 19304
rect 6880 19252 6886 19304
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 9309 19295 9367 19301
rect 9309 19292 9321 19295
rect 9272 19264 9321 19292
rect 9272 19252 9278 19264
rect 9309 19261 9321 19264
rect 9355 19261 9367 19295
rect 11072 19292 11100 19332
rect 11974 19320 11980 19332
rect 12032 19360 12038 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 12032 19332 12173 19360
rect 12032 19320 12038 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 14642 19360 14648 19372
rect 13955 19332 14648 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 17052 19369 17080 19400
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 17865 19431 17923 19437
rect 17865 19428 17877 19431
rect 17644 19400 17877 19428
rect 17644 19388 17650 19400
rect 17865 19397 17877 19400
rect 17911 19397 17923 19431
rect 17865 19391 17923 19397
rect 18785 19431 18843 19437
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 19242 19428 19248 19440
rect 18831 19400 19248 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 19242 19388 19248 19400
rect 19300 19388 19306 19440
rect 19812 19428 19840 19468
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20254 19496 20260 19508
rect 19935 19468 20260 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20717 19499 20775 19505
rect 20717 19465 20729 19499
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 20530 19428 20536 19440
rect 19812 19400 20536 19428
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 20732 19428 20760 19459
rect 21174 19456 21180 19508
rect 21232 19456 21238 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 21968 19468 23765 19496
rect 21968 19456 21974 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 21450 19428 21456 19440
rect 20732 19400 21456 19428
rect 21450 19388 21456 19400
rect 21508 19388 21514 19440
rect 23566 19428 23572 19440
rect 23506 19400 23572 19428
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 19576 19332 19809 19360
rect 19576 19320 19582 19332
rect 19797 19329 19809 19332
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 19944 19332 21097 19360
rect 19944 19320 19950 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 9309 19255 9367 19261
rect 10888 19264 11100 19292
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 7616 19128 8309 19156
rect 7616 19116 7622 19128
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10888 19165 10916 19264
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 12268 19224 12296 19255
rect 13354 19224 13360 19236
rect 11072 19196 13360 19224
rect 11072 19168 11100 19196
rect 13354 19184 13360 19196
rect 13412 19224 13418 19236
rect 13412 19196 13860 19224
rect 13412 19184 13418 19196
rect 10873 19159 10931 19165
rect 10873 19156 10885 19159
rect 10284 19128 10885 19156
rect 10284 19116 10290 19128
rect 10873 19125 10885 19128
rect 10919 19125 10931 19159
rect 10873 19119 10931 19125
rect 11054 19116 11060 19168
rect 11112 19116 11118 19168
rect 13538 19116 13544 19168
rect 13596 19116 13602 19168
rect 13832 19156 13860 19196
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 14108 19224 14136 19255
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17736 19264 17969 19292
rect 17736 19252 17742 19264
rect 17957 19261 17969 19264
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 19334 19292 19340 19304
rect 18187 19264 19340 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 20073 19295 20131 19301
rect 20073 19261 20085 19295
rect 20119 19292 20131 19295
rect 21266 19292 21272 19304
rect 20119 19264 21272 19292
rect 20119 19261 20131 19264
rect 20073 19255 20131 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21910 19292 21916 19304
rect 21407 19264 21916 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 22002 19252 22008 19304
rect 22060 19252 22066 19304
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 14737 19227 14795 19233
rect 14737 19224 14749 19227
rect 13964 19196 14136 19224
rect 14200 19196 14749 19224
rect 13964 19184 13970 19196
rect 14200 19156 14228 19196
rect 14737 19193 14749 19196
rect 14783 19224 14795 19227
rect 14826 19224 14832 19236
rect 14783 19196 14832 19224
rect 14783 19193 14795 19196
rect 14737 19187 14795 19193
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 18969 19227 19027 19233
rect 18969 19193 18981 19227
rect 19015 19224 19027 19227
rect 19242 19224 19248 19236
rect 19015 19196 19248 19224
rect 19015 19193 19027 19196
rect 18969 19187 19027 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 13832 19128 14228 19156
rect 14642 19116 14648 19168
rect 14700 19116 14706 19168
rect 19429 19159 19487 19165
rect 19429 19125 19441 19159
rect 19475 19156 19487 19159
rect 20714 19156 20720 19168
rect 19475 19128 20720 19156
rect 19475 19125 19487 19128
rect 19429 19119 19487 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 24121 19159 24179 19165
rect 24121 19125 24133 19159
rect 24167 19156 24179 19159
rect 24394 19156 24400 19168
rect 24167 19128 24400 19156
rect 24167 19125 24179 19128
rect 24121 19119 24179 19125
rect 24394 19116 24400 19128
rect 24452 19116 24458 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 10594 18952 10600 18964
rect 5224 18924 10600 18952
rect 5224 18912 5230 18924
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11296 18924 11897 18952
rect 11296 18912 11302 18924
rect 11885 18921 11897 18924
rect 11931 18921 11943 18955
rect 11885 18915 11943 18921
rect 12158 18912 12164 18964
rect 12216 18912 12222 18964
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 14240 18924 14289 18952
rect 14240 18912 14246 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 16040 18924 17540 18952
rect 8938 18844 8944 18896
rect 8996 18844 9002 18896
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1360 18788 2053 18816
rect 1360 18776 1366 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 9401 18819 9459 18825
rect 9401 18816 9413 18819
rect 6236 18788 9413 18816
rect 6236 18776 6242 18788
rect 9401 18785 9413 18788
rect 9447 18816 9459 18819
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9447 18788 10057 18816
rect 9447 18785 9459 18788
rect 9401 18779 9459 18785
rect 10045 18785 10057 18788
rect 10091 18816 10103 18819
rect 11054 18816 11060 18828
rect 10091 18788 11060 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9232 18720 9781 18748
rect 9232 18689 9260 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 11256 18748 11284 18912
rect 11330 18844 11336 18896
rect 11388 18884 11394 18896
rect 13906 18884 13912 18896
rect 11388 18856 13912 18884
rect 11388 18844 11394 18856
rect 13906 18844 13912 18856
rect 13964 18844 13970 18896
rect 12710 18776 12716 18828
rect 12768 18816 12774 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12768 18788 13553 18816
rect 12768 18776 12774 18788
rect 13541 18785 13553 18788
rect 13587 18816 13599 18819
rect 14366 18816 14372 18828
rect 13587 18788 14372 18816
rect 13587 18785 13599 18788
rect 13541 18779 13599 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 11178 18720 11284 18748
rect 13449 18751 13507 18757
rect 9769 18711 9827 18717
rect 13449 18717 13461 18751
rect 13495 18748 13507 18751
rect 13814 18748 13820 18760
rect 13495 18720 13820 18748
rect 13495 18717 13507 18720
rect 13449 18711 13507 18717
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 16040 18748 16068 18924
rect 17512 18884 17540 18924
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18325 18955 18383 18961
rect 18325 18952 18337 18955
rect 17736 18924 18337 18952
rect 17736 18912 17742 18924
rect 18325 18921 18337 18924
rect 18371 18921 18383 18955
rect 18325 18915 18383 18921
rect 19058 18912 19064 18964
rect 19116 18912 19122 18964
rect 22278 18912 22284 18964
rect 22336 18952 22342 18964
rect 24029 18955 24087 18961
rect 24029 18952 24041 18955
rect 22336 18924 24041 18952
rect 22336 18912 22342 18924
rect 24029 18921 24041 18924
rect 24075 18921 24087 18955
rect 24029 18915 24087 18921
rect 24394 18912 24400 18964
rect 24452 18912 24458 18964
rect 18966 18884 18972 18896
rect 17512 18856 18972 18884
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 16482 18776 16488 18828
rect 16540 18816 16546 18828
rect 17957 18819 18015 18825
rect 17957 18816 17969 18819
rect 16540 18788 17969 18816
rect 16540 18776 16546 18788
rect 17957 18785 17969 18788
rect 18003 18785 18015 18819
rect 17957 18779 18015 18785
rect 14691 18720 16068 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 16206 18708 16212 18760
rect 16264 18708 16270 18760
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19116 18720 19625 18748
rect 19116 18708 19122 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20349 18751 20407 18757
rect 20349 18717 20361 18751
rect 20395 18748 20407 18751
rect 20438 18748 20444 18760
rect 20395 18720 20444 18748
rect 20395 18717 20407 18720
rect 20349 18711 20407 18717
rect 20438 18708 20444 18720
rect 20496 18748 20502 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 20496 18720 21557 18748
rect 20496 18708 20502 18720
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 22060 18720 22293 18748
rect 22060 18708 22066 18720
rect 9217 18683 9275 18689
rect 9217 18680 9229 18683
rect 8496 18652 9229 18680
rect 8496 18624 8524 18652
rect 9217 18649 9229 18652
rect 9263 18649 9275 18683
rect 16485 18683 16543 18689
rect 9217 18643 9275 18649
rect 11348 18652 12434 18680
rect 8478 18572 8484 18624
rect 8536 18572 8542 18624
rect 8665 18615 8723 18621
rect 8665 18581 8677 18615
rect 8711 18612 8723 18615
rect 8846 18612 8852 18624
rect 8711 18584 8852 18612
rect 8711 18581 8723 18584
rect 8665 18575 8723 18581
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11348 18612 11376 18652
rect 10928 18584 11376 18612
rect 11517 18615 11575 18621
rect 10928 18572 10934 18584
rect 11517 18581 11529 18615
rect 11563 18612 11575 18615
rect 11606 18612 11612 18624
rect 11563 18584 11612 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 12406 18612 12434 18652
rect 16485 18649 16497 18683
rect 16531 18649 16543 18683
rect 18414 18680 18420 18692
rect 17710 18652 18420 18680
rect 16485 18643 16543 18649
rect 12989 18615 13047 18621
rect 12989 18612 13001 18615
rect 12406 18584 13001 18612
rect 12989 18581 13001 18584
rect 13035 18581 13047 18615
rect 12989 18575 13047 18581
rect 13354 18572 13360 18624
rect 13412 18572 13418 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 14737 18615 14795 18621
rect 14737 18612 14749 18615
rect 13780 18584 14749 18612
rect 13780 18572 13786 18584
rect 14737 18581 14749 18584
rect 14783 18581 14795 18615
rect 16500 18612 16528 18643
rect 18414 18640 18420 18652
rect 18472 18680 18478 18692
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 18472 18652 18521 18680
rect 18472 18640 18478 18652
rect 18509 18649 18521 18652
rect 18555 18680 18567 18683
rect 19426 18680 19432 18692
rect 18555 18652 19432 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 21085 18683 21143 18689
rect 21085 18680 21097 18683
rect 20956 18652 21097 18680
rect 20956 18640 20962 18652
rect 21085 18649 21097 18652
rect 21131 18680 21143 18683
rect 22112 18680 22140 18720
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 21131 18652 22140 18680
rect 21131 18649 21143 18652
rect 21085 18643 21143 18649
rect 22554 18640 22560 18692
rect 22612 18640 22618 18692
rect 24394 18680 24400 18692
rect 23782 18652 24400 18680
rect 24394 18640 24400 18652
rect 24452 18640 24458 18692
rect 18322 18612 18328 18624
rect 16500 18584 18328 18612
rect 14737 18575 14795 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 7742 18368 7748 18420
rect 7800 18368 7806 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 8496 18380 9781 18408
rect 8496 18349 8524 18380
rect 9769 18377 9781 18380
rect 9815 18408 9827 18411
rect 9950 18408 9956 18420
rect 9815 18380 9956 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10410 18368 10416 18420
rect 10468 18368 10474 18420
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 12158 18408 12164 18420
rect 10827 18380 12164 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13412 18380 14289 18408
rect 13412 18368 13418 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 14691 18380 15393 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 15381 18377 15393 18380
rect 15427 18408 15439 18411
rect 18690 18408 18696 18420
rect 15427 18380 18696 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 18690 18368 18696 18380
rect 18748 18408 18754 18420
rect 18874 18408 18880 18420
rect 18748 18380 18880 18408
rect 18748 18368 18754 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 19334 18368 19340 18420
rect 19392 18368 19398 18420
rect 8481 18343 8539 18349
rect 8481 18309 8493 18343
rect 8527 18309 8539 18343
rect 8481 18303 8539 18309
rect 11146 18300 11152 18352
rect 11204 18340 11210 18352
rect 11606 18340 11612 18352
rect 11204 18312 11612 18340
rect 11204 18300 11210 18312
rect 11606 18300 11612 18312
rect 11664 18300 11670 18352
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 13538 18340 13544 18352
rect 12115 18312 13544 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 13633 18343 13691 18349
rect 13633 18309 13645 18343
rect 13679 18340 13691 18343
rect 14090 18340 14096 18352
rect 13679 18312 14096 18340
rect 13679 18309 13691 18312
rect 13633 18303 13691 18309
rect 7653 18275 7711 18281
rect 7653 18272 7665 18275
rect 6932 18244 7665 18272
rect 4890 18028 4896 18080
rect 4948 18068 4954 18080
rect 6932 18077 6960 18244
rect 7653 18241 7665 18244
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 9858 18232 9864 18284
rect 9916 18272 9922 18284
rect 10042 18272 10048 18284
rect 9916 18244 10048 18272
rect 9916 18232 9922 18244
rect 10042 18232 10048 18244
rect 10100 18272 10106 18284
rect 11330 18272 11336 18284
rect 10100 18244 11336 18272
rect 10100 18232 10106 18244
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7616 18176 7849 18204
rect 7616 18164 7622 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8536 18176 9229 18204
rect 8536 18164 8542 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10686 18204 10692 18216
rect 10183 18176 10692 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10686 18164 10692 18176
rect 10744 18204 10750 18216
rect 10980 18213 11008 18244
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10744 18176 10885 18204
rect 10744 18164 10750 18176
rect 10873 18173 10885 18176
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 12158 18164 12164 18216
rect 12216 18164 12222 18216
rect 12342 18164 12348 18216
rect 12400 18164 12406 18216
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 11701 18139 11759 18145
rect 11701 18136 11713 18139
rect 10836 18108 11713 18136
rect 10836 18096 10842 18108
rect 11701 18105 11713 18108
rect 11747 18105 11759 18139
rect 13648 18136 13676 18303
rect 14090 18300 14096 18312
rect 14148 18300 14154 18352
rect 17221 18343 17279 18349
rect 17221 18309 17233 18343
rect 17267 18340 17279 18343
rect 17494 18340 17500 18352
rect 17267 18312 17500 18340
rect 17267 18309 17279 18312
rect 17221 18303 17279 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 19153 18343 19211 18349
rect 19153 18309 19165 18343
rect 19199 18340 19211 18343
rect 19352 18340 19380 18368
rect 19199 18312 19380 18340
rect 19199 18309 19211 18312
rect 19153 18303 19211 18309
rect 19426 18300 19432 18352
rect 19484 18340 19490 18352
rect 19484 18312 19642 18340
rect 19484 18300 19490 18312
rect 21082 18300 21088 18352
rect 21140 18340 21146 18352
rect 21269 18343 21327 18349
rect 21269 18340 21281 18343
rect 21140 18312 21281 18340
rect 21140 18300 21146 18312
rect 21269 18309 21281 18312
rect 21315 18309 21327 18343
rect 21269 18303 21327 18309
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13780 18244 13921 18272
rect 13780 18232 13786 18244
rect 13909 18241 13921 18244
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14737 18207 14795 18213
rect 14737 18204 14749 18207
rect 13872 18176 14749 18204
rect 13872 18164 13878 18176
rect 14737 18173 14749 18176
rect 14783 18173 14795 18207
rect 14737 18167 14795 18173
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18204 14979 18207
rect 15378 18204 15384 18216
rect 14967 18176 15384 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 14936 18136 14964 18167
rect 15378 18164 15384 18176
rect 15436 18204 15442 18216
rect 16022 18204 16028 18216
rect 15436 18176 16028 18204
rect 15436 18164 15442 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 16482 18204 16488 18216
rect 16264 18176 16488 18204
rect 16264 18164 16270 18176
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 16540 18176 18337 18204
rect 16540 18164 16546 18176
rect 18325 18173 18337 18176
rect 18371 18204 18383 18207
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18371 18176 18889 18204
rect 18371 18173 18383 18176
rect 18325 18167 18383 18173
rect 18877 18173 18889 18176
rect 18923 18173 18935 18207
rect 18877 18167 18935 18173
rect 20162 18164 20168 18216
rect 20220 18204 20226 18216
rect 21082 18204 21088 18216
rect 20220 18176 21088 18204
rect 20220 18164 20226 18176
rect 21082 18164 21088 18176
rect 21140 18164 21146 18216
rect 23293 18207 23351 18213
rect 23293 18173 23305 18207
rect 23339 18204 23351 18207
rect 23382 18204 23388 18216
rect 23339 18176 23388 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 23382 18164 23388 18176
rect 23440 18164 23446 18216
rect 24762 18164 24768 18216
rect 24820 18164 24826 18216
rect 11701 18099 11759 18105
rect 12406 18108 13676 18136
rect 13740 18108 14964 18136
rect 21453 18139 21511 18145
rect 6917 18071 6975 18077
rect 6917 18068 6929 18071
rect 4948 18040 6929 18068
rect 4948 18028 4954 18040
rect 6917 18037 6929 18040
rect 6963 18037 6975 18071
rect 6917 18031 6975 18037
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 8662 18068 8668 18080
rect 7331 18040 8668 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 12406 18068 12434 18108
rect 13740 18080 13768 18108
rect 21453 18105 21465 18139
rect 21499 18136 21511 18139
rect 22738 18136 22744 18148
rect 21499 18108 22744 18136
rect 21499 18105 21511 18108
rect 21453 18099 21511 18105
rect 22738 18096 22744 18108
rect 22796 18096 22802 18148
rect 11296 18040 12434 18068
rect 11296 18028 11302 18040
rect 13722 18028 13728 18080
rect 13780 18028 13786 18080
rect 13814 18028 13820 18080
rect 13872 18028 13878 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20220 18040 20637 18068
rect 20220 18028 20226 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 6270 17824 6276 17876
rect 6328 17824 6334 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 7432 17836 9137 17864
rect 7432 17824 7438 17836
rect 9125 17833 9137 17836
rect 9171 17833 9183 17867
rect 9125 17827 9183 17833
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 12529 17867 12587 17873
rect 12529 17864 12541 17867
rect 12032 17836 12541 17864
rect 12032 17824 12038 17836
rect 12529 17833 12541 17836
rect 12575 17864 12587 17867
rect 12618 17864 12624 17876
rect 12575 17836 12624 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 19518 17864 19524 17876
rect 15896 17836 19524 17864
rect 15896 17824 15902 17836
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 21266 17824 21272 17876
rect 21324 17864 21330 17876
rect 21637 17867 21695 17873
rect 21637 17864 21649 17867
rect 21324 17836 21649 17864
rect 21324 17824 21330 17836
rect 21637 17833 21649 17836
rect 21683 17864 21695 17867
rect 21683 17836 22232 17864
rect 21683 17833 21695 17836
rect 21637 17827 21695 17833
rect 15562 17796 15568 17808
rect 14660 17768 15568 17796
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 6914 17728 6920 17740
rect 6871 17700 6920 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 6914 17688 6920 17700
rect 6972 17688 6978 17740
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7892 17700 7941 17728
rect 7892 17688 7898 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 8386 17728 8392 17740
rect 8159 17700 8392 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9456 17700 9689 17728
rect 9456 17688 9462 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 11885 17731 11943 17737
rect 11885 17728 11897 17731
rect 9677 17691 9735 17697
rect 9784 17700 11897 17728
rect 4522 17620 4528 17672
rect 4580 17660 4586 17672
rect 4580 17632 8800 17660
rect 4580 17620 4586 17632
rect 6641 17595 6699 17601
rect 6641 17561 6653 17595
rect 6687 17592 6699 17595
rect 6687 17564 7512 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 7282 17524 7288 17536
rect 6779 17496 7288 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 7484 17533 7512 17564
rect 8772 17536 8800 17632
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 9784 17660 9812 17700
rect 11885 17697 11897 17700
rect 11931 17697 11943 17731
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 11885 17691 11943 17697
rect 12406 17700 12725 17728
rect 9640 17632 9812 17660
rect 9640 17620 9646 17632
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10502 17660 10508 17672
rect 10008 17632 10508 17660
rect 10008 17620 10014 17632
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 12406 17660 12434 17700
rect 12713 17697 12725 17700
rect 12759 17728 12771 17731
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 12759 17700 13553 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 11756 17632 12434 17660
rect 11756 17620 11762 17632
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 12676 17632 13461 17660
rect 12676 17620 12682 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 14660 17660 14688 17768
rect 15562 17756 15568 17768
rect 15620 17796 15626 17808
rect 16114 17796 16120 17808
rect 15620 17768 16120 17796
rect 15620 17756 15626 17768
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16209 17799 16267 17805
rect 16209 17765 16221 17799
rect 16255 17796 16267 17799
rect 18874 17796 18880 17808
rect 16255 17768 18880 17796
rect 16255 17765 16267 17768
rect 16209 17759 16267 17765
rect 18874 17756 18880 17768
rect 18932 17756 18938 17808
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16356 17700 16681 17728
rect 16356 17688 16362 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16853 17731 16911 17737
rect 16853 17697 16865 17731
rect 16899 17728 16911 17731
rect 17126 17728 17132 17740
rect 16899 17700 17132 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 13449 17623 13507 17629
rect 14016 17632 14688 17660
rect 11330 17552 11336 17604
rect 11388 17552 11394 17604
rect 13357 17595 13415 17601
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 14016 17592 14044 17632
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 14792 17632 15577 17660
rect 14792 17620 14798 17632
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 16684 17660 16712 17691
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 19889 17731 19947 17737
rect 19889 17697 19901 17731
rect 19935 17728 19947 17731
rect 20898 17728 20904 17740
rect 19935 17700 20904 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 20898 17688 20904 17700
rect 20956 17728 20962 17740
rect 22097 17731 22155 17737
rect 22097 17728 22109 17731
rect 20956 17700 22109 17728
rect 20956 17688 20962 17700
rect 22097 17697 22109 17700
rect 22143 17697 22155 17731
rect 22204 17728 22232 17836
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 23845 17867 23903 17873
rect 23845 17864 23857 17867
rect 22612 17836 23857 17864
rect 22612 17824 22618 17836
rect 23845 17833 23857 17836
rect 23891 17833 23903 17867
rect 23845 17827 23903 17833
rect 24213 17867 24271 17873
rect 24213 17833 24225 17867
rect 24259 17864 24271 17867
rect 24394 17864 24400 17876
rect 24259 17836 24400 17864
rect 24259 17833 24271 17836
rect 24213 17827 24271 17833
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 22204 17700 22385 17728
rect 22097 17691 22155 17697
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 17221 17663 17279 17669
rect 17221 17660 17233 17663
rect 16684 17632 17233 17660
rect 15565 17623 15623 17629
rect 17221 17629 17233 17632
rect 17267 17629 17279 17663
rect 23842 17660 23848 17672
rect 23506 17632 23848 17660
rect 17221 17623 17279 17629
rect 23842 17620 23848 17632
rect 23900 17660 23906 17672
rect 24228 17660 24256 17827
rect 24394 17824 24400 17836
rect 24452 17824 24458 17876
rect 23900 17632 24256 17660
rect 23900 17620 23906 17632
rect 24854 17620 24860 17672
rect 24912 17620 24918 17672
rect 13403 17564 14044 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 14090 17552 14096 17604
rect 14148 17592 14154 17604
rect 14148 17564 14780 17592
rect 14148 17552 14154 17564
rect 7469 17527 7527 17533
rect 7469 17493 7481 17527
rect 7515 17493 7527 17527
rect 7469 17487 7527 17493
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8570 17524 8576 17536
rect 7883 17496 8576 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8754 17484 8760 17536
rect 8812 17484 8818 17536
rect 9490 17484 9496 17536
rect 9548 17484 9554 17536
rect 9585 17527 9643 17533
rect 9585 17493 9597 17527
rect 9631 17524 9643 17527
rect 10134 17524 10140 17536
rect 9631 17496 10140 17524
rect 9631 17493 9643 17496
rect 9585 17487 9643 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12989 17527 13047 17533
rect 12989 17524 13001 17527
rect 12768 17496 13001 17524
rect 12768 17484 12774 17496
rect 12989 17493 13001 17496
rect 13035 17493 13047 17527
rect 12989 17487 13047 17493
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 13596 17496 14289 17524
rect 13596 17484 13602 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 14277 17487 14335 17493
rect 14642 17484 14648 17536
rect 14700 17484 14706 17536
rect 14752 17533 14780 17564
rect 20162 17552 20168 17604
rect 20220 17552 20226 17604
rect 20272 17564 20654 17592
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17493 14795 17527
rect 14737 17487 14795 17493
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15620 17496 15669 17524
rect 15620 17484 15626 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 16574 17484 16580 17536
rect 16632 17484 16638 17536
rect 19426 17484 19432 17536
rect 19484 17524 19490 17536
rect 20272 17524 20300 17564
rect 19484 17496 20300 17524
rect 19484 17484 19490 17496
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24268 17496 24685 17524
rect 24268 17484 24274 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4120 17292 8156 17320
rect 4120 17280 4126 17292
rect 7958 17156 8064 17184
rect 6546 17076 6552 17128
rect 6604 17076 6610 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 8036 17048 8064 17156
rect 8128 17116 8156 17292
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9548 17292 10057 17320
rect 9548 17280 9554 17292
rect 10045 17289 10057 17292
rect 10091 17289 10103 17323
rect 10045 17283 10103 17289
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 10560 17292 11529 17320
rect 10560 17280 10566 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 13722 17320 13728 17332
rect 12584 17292 13728 17320
rect 12584 17280 12590 17292
rect 8573 17255 8631 17261
rect 8573 17221 8585 17255
rect 8619 17252 8631 17255
rect 9858 17252 9864 17264
rect 8619 17224 9864 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 10413 17255 10471 17261
rect 10413 17221 10425 17255
rect 10459 17252 10471 17255
rect 12066 17252 12072 17264
rect 10459 17224 12072 17252
rect 10459 17221 10471 17224
rect 10413 17215 10471 17221
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 12912 17261 12940 17292
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 13872 17292 16037 17320
rect 13872 17280 13878 17292
rect 16025 17289 16037 17292
rect 16071 17320 16083 17323
rect 16574 17320 16580 17332
rect 16071 17292 16580 17320
rect 16071 17289 16083 17292
rect 16025 17283 16083 17289
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 20898 17320 20904 17332
rect 17696 17292 20904 17320
rect 12897 17255 12955 17261
rect 12897 17221 12909 17255
rect 12943 17221 12955 17255
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 14122 17238 14933 17252
rect 12897 17215 12955 17221
rect 14108 17224 14933 17238
rect 8754 17144 8760 17196
rect 8812 17184 8818 17196
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8812 17156 9045 17184
rect 8812 17144 8818 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 12526 17184 12532 17196
rect 9272 17156 12532 17184
rect 9272 17144 9278 17156
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 8128 17088 9505 17116
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 10502 17076 10508 17128
rect 10560 17076 10566 17128
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10962 17116 10968 17128
rect 10735 17088 10968 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11388 17088 12633 17116
rect 11388 17076 11394 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 14108 17116 14136 17224
rect 14921 17221 14933 17224
rect 14967 17221 14979 17255
rect 14921 17215 14979 17221
rect 14826 17144 14832 17196
rect 14884 17144 14890 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 17696 17193 17724 17292
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 23842 17320 23848 17332
rect 21560 17292 23848 17320
rect 18414 17212 18420 17264
rect 18472 17212 18478 17264
rect 19426 17212 19432 17264
rect 19484 17252 19490 17264
rect 21560 17261 21588 17292
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 19705 17255 19763 17261
rect 19705 17252 19717 17255
rect 19484 17224 19717 17252
rect 19484 17212 19490 17224
rect 19705 17221 19717 17224
rect 19751 17252 19763 17255
rect 20993 17255 21051 17261
rect 20993 17252 21005 17255
rect 19751 17224 21005 17252
rect 19751 17221 19763 17224
rect 19705 17215 19763 17221
rect 20993 17221 21005 17224
rect 21039 17252 21051 17255
rect 21545 17255 21603 17261
rect 21545 17252 21557 17255
rect 21039 17224 21557 17252
rect 21039 17221 21051 17224
rect 20993 17215 21051 17221
rect 21545 17221 21557 17224
rect 21591 17221 21603 17255
rect 21545 17215 21603 17221
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 22833 17255 22891 17261
rect 22833 17252 22845 17255
rect 22520 17224 22845 17252
rect 22520 17212 22526 17224
rect 22833 17221 22845 17224
rect 22879 17221 22891 17255
rect 22833 17215 22891 17221
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16724 17156 17049 17184
rect 16724 17144 16730 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 17681 17147 17739 17153
rect 19168 17156 22109 17184
rect 19168 17128 19196 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 23750 17144 23756 17196
rect 23808 17184 23814 17196
rect 23937 17187 23995 17193
rect 23937 17184 23949 17187
rect 23808 17156 23949 17184
rect 23808 17144 23814 17156
rect 23937 17153 23949 17156
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 13412 17088 14136 17116
rect 13412 17076 13418 17088
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 17957 17119 18015 17125
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18598 17116 18604 17128
rect 18003 17088 18604 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19150 17076 19156 17128
rect 19208 17076 19214 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19429 17119 19487 17125
rect 19429 17116 19441 17119
rect 19392 17088 19441 17116
rect 19392 17076 19398 17088
rect 19429 17085 19441 17088
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 20438 17076 20444 17128
rect 20496 17076 20502 17128
rect 24670 17076 24676 17128
rect 24728 17076 24734 17128
rect 8294 17048 8300 17060
rect 8036 17020 8300 17048
rect 8294 17008 8300 17020
rect 8352 17048 8358 17060
rect 8938 17048 8944 17060
rect 8352 17020 8944 17048
rect 8352 17008 8358 17020
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 14642 17008 14648 17060
rect 14700 17048 14706 17060
rect 15197 17051 15255 17057
rect 15197 17048 15209 17051
rect 14700 17020 15209 17048
rect 14700 17008 14706 17020
rect 15197 17017 15209 17020
rect 15243 17048 15255 17051
rect 22281 17051 22339 17057
rect 15243 17020 16988 17048
rect 15243 17017 15255 17020
rect 15197 17011 15255 17017
rect 7006 16940 7012 16992
rect 7064 16980 7070 16992
rect 7466 16980 7472 16992
rect 7064 16952 7472 16980
rect 7064 16940 7070 16952
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 9306 16940 9312 16992
rect 9364 16940 9370 16992
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 16960 16980 16988 17020
rect 22281 17017 22293 17051
rect 22327 17048 22339 17051
rect 22646 17048 22652 17060
rect 22327 17020 22652 17048
rect 22327 17017 22339 17020
rect 22281 17011 22339 17017
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 23017 17051 23075 17057
rect 23017 17017 23029 17051
rect 23063 17048 23075 17051
rect 23290 17048 23296 17060
rect 23063 17020 23296 17048
rect 23063 17017 23075 17020
rect 23017 17011 23075 17017
rect 23290 17008 23296 17020
rect 23348 17008 23354 17060
rect 19058 16980 19064 16992
rect 16960 16952 19064 16980
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 5616 16779 5674 16785
rect 5616 16745 5628 16779
rect 5662 16776 5674 16779
rect 5662 16748 6868 16776
rect 5662 16745 5674 16748
rect 5616 16739 5674 16745
rect 6840 16708 6868 16748
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7101 16779 7159 16785
rect 7101 16776 7113 16779
rect 6972 16748 7113 16776
rect 6972 16736 6978 16748
rect 7101 16745 7113 16748
rect 7147 16745 7159 16779
rect 7101 16739 7159 16745
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 8294 16776 8300 16788
rect 7524 16748 8300 16776
rect 7524 16736 7530 16748
rect 8294 16736 8300 16748
rect 8352 16776 8358 16788
rect 8352 16748 8524 16776
rect 8352 16736 8358 16748
rect 8386 16708 8392 16720
rect 6840 16680 8392 16708
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 8496 16708 8524 16748
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 8628 16748 9137 16776
rect 8628 16736 8634 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10505 16779 10563 16785
rect 10505 16776 10517 16779
rect 10192 16748 10517 16776
rect 10192 16736 10198 16748
rect 10505 16745 10517 16748
rect 10551 16745 10563 16779
rect 11606 16776 11612 16788
rect 10505 16739 10563 16745
rect 10888 16748 11612 16776
rect 8665 16711 8723 16717
rect 8665 16708 8677 16711
rect 8496 16680 8677 16708
rect 8665 16677 8677 16680
rect 8711 16708 8723 16711
rect 8754 16708 8760 16720
rect 8711 16680 8760 16708
rect 8711 16677 8723 16680
rect 8665 16671 8723 16677
rect 8754 16668 8760 16680
rect 8812 16668 8818 16720
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 9364 16680 10241 16708
rect 9364 16668 9370 16680
rect 10229 16677 10241 16680
rect 10275 16708 10287 16711
rect 10888 16708 10916 16748
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 23842 16736 23848 16788
rect 23900 16736 23906 16788
rect 14274 16708 14280 16720
rect 10275 16680 10916 16708
rect 10980 16680 14280 16708
rect 10275 16677 10287 16680
rect 10229 16671 10287 16677
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 6638 16640 6644 16652
rect 5399 16612 6644 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 6638 16600 6644 16612
rect 6696 16640 6702 16652
rect 7653 16643 7711 16649
rect 7653 16640 7665 16643
rect 6696 16612 7665 16640
rect 6696 16600 6702 16612
rect 7653 16609 7665 16612
rect 7699 16640 7711 16643
rect 8478 16640 8484 16652
rect 7699 16612 8484 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 10980 16649 11008 16680
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 19334 16708 19340 16720
rect 15764 16680 19340 16708
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9416 16612 9689 16640
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 1544 16544 1593 16572
rect 1544 16532 1550 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 7466 16572 7472 16584
rect 6762 16544 7472 16572
rect 1581 16535 1639 16541
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 9214 16572 9220 16584
rect 8352 16544 9220 16572
rect 8352 16532 8358 16544
rect 9214 16532 9220 16544
rect 9272 16572 9278 16584
rect 9416 16572 9444 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11054 16600 11060 16652
rect 11112 16600 11118 16652
rect 12250 16600 12256 16652
rect 12308 16600 12314 16652
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16640 12403 16643
rect 12618 16640 12624 16652
rect 12391 16612 12624 16640
rect 12391 16609 12403 16612
rect 12345 16603 12403 16609
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16640 15071 16643
rect 15102 16640 15108 16652
rect 15059 16612 15108 16640
rect 15059 16609 15071 16612
rect 15013 16603 15071 16609
rect 15102 16600 15108 16612
rect 15160 16640 15166 16652
rect 15764 16649 15792 16680
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15160 16612 15761 16640
rect 15160 16600 15166 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16022 16640 16028 16652
rect 15979 16612 16028 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16022 16600 16028 16612
rect 16080 16600 16086 16652
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20625 16643 20683 16649
rect 20625 16640 20637 16643
rect 20220 16612 20637 16640
rect 20220 16600 20226 16612
rect 20625 16609 20637 16612
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21729 16643 21787 16649
rect 21729 16640 21741 16643
rect 20956 16612 21741 16640
rect 20956 16600 20962 16612
rect 21729 16609 21741 16612
rect 21775 16609 21787 16643
rect 21729 16603 21787 16609
rect 22002 16600 22008 16652
rect 22060 16600 22066 16652
rect 23382 16640 23388 16652
rect 23124 16612 23388 16640
rect 9272 16544 9444 16572
rect 9493 16575 9551 16581
rect 9272 16532 9278 16544
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 9582 16572 9588 16584
rect 9539 16544 9588 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10870 16532 10876 16584
rect 10928 16532 10934 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12710 16572 12716 16584
rect 12207 16544 12716 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 23124 16558 23152 16612
rect 23382 16600 23388 16612
rect 23440 16640 23446 16652
rect 23860 16640 23888 16736
rect 23440 16612 23888 16640
rect 23440 16600 23446 16612
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 10318 16504 10324 16516
rect 2501 16467 2559 16473
rect 9968 16476 10324 16504
rect 9968 16448 9996 16476
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 12066 16464 12072 16516
rect 12124 16504 12130 16516
rect 22094 16504 22100 16516
rect 12124 16476 12434 16504
rect 12124 16464 12130 16476
rect 8478 16396 8484 16448
rect 8536 16396 8542 16448
rect 9585 16439 9643 16445
rect 9585 16405 9597 16439
rect 9631 16436 9643 16439
rect 9950 16436 9956 16448
rect 9631 16408 9956 16436
rect 9631 16405 9643 16408
rect 9585 16399 9643 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 12406 16436 12434 16476
rect 20088 16476 22100 16504
rect 13814 16436 13820 16448
rect 12406 16408 13820 16436
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 15286 16396 15292 16448
rect 15344 16396 15350 16448
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16436 15715 16439
rect 15746 16436 15752 16448
rect 15703 16408 15752 16436
rect 15703 16405 15715 16408
rect 15657 16399 15715 16405
rect 15746 16396 15752 16408
rect 15804 16436 15810 16448
rect 16393 16439 16451 16445
rect 16393 16436 16405 16439
rect 15804 16408 16405 16436
rect 15804 16396 15810 16408
rect 16393 16405 16405 16408
rect 16439 16436 16451 16439
rect 16942 16436 16948 16448
rect 16439 16408 16948 16436
rect 16439 16405 16451 16408
rect 16393 16399 16451 16405
rect 16942 16396 16948 16408
rect 17000 16396 17006 16448
rect 20088 16445 20116 16476
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 23477 16439 23535 16445
rect 23477 16436 23489 16439
rect 21232 16408 23489 16436
rect 21232 16396 21238 16408
rect 23477 16405 23489 16408
rect 23523 16405 23535 16439
rect 23477 16399 23535 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 7340 16204 8953 16232
rect 7340 16192 7346 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 10502 16232 10508 16244
rect 10183 16204 10508 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 11422 16232 11428 16244
rect 10643 16204 11428 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11701 16235 11759 16241
rect 11701 16232 11713 16235
rect 11572 16204 11713 16232
rect 11572 16192 11578 16204
rect 11701 16201 11713 16204
rect 11747 16201 11759 16235
rect 11701 16195 11759 16201
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 12584 16204 13093 16232
rect 12584 16192 12590 16204
rect 13081 16201 13093 16204
rect 13127 16232 13139 16235
rect 13354 16232 13360 16244
rect 13127 16204 13360 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13504 16204 13737 16232
rect 13504 16192 13510 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 14734 16192 14740 16244
rect 14792 16192 14798 16244
rect 18598 16192 18604 16244
rect 18656 16192 18662 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16232 19303 16235
rect 19886 16232 19892 16244
rect 19291 16204 19892 16232
rect 19291 16201 19303 16204
rect 19245 16195 19303 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 22465 16235 22523 16241
rect 22465 16232 22477 16235
rect 20772 16204 22477 16232
rect 20772 16192 20778 16204
rect 22465 16201 22477 16204
rect 22511 16201 22523 16235
rect 22465 16195 22523 16201
rect 23201 16235 23259 16241
rect 23201 16201 23213 16235
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 2501 16167 2559 16173
rect 2501 16133 2513 16167
rect 2547 16164 2559 16167
rect 4062 16164 4068 16176
rect 2547 16136 4068 16164
rect 2547 16133 2559 16136
rect 2501 16127 2559 16133
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 7466 16124 7472 16176
rect 7524 16124 7530 16176
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 11790 16164 11796 16176
rect 9355 16136 11796 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 12069 16167 12127 16173
rect 12069 16133 12081 16167
rect 12115 16164 12127 16167
rect 13538 16164 13544 16176
rect 12115 16136 13544 16164
rect 12115 16133 12127 16136
rect 12069 16127 12127 16133
rect 13538 16124 13544 16136
rect 13596 16124 13602 16176
rect 14185 16167 14243 16173
rect 14185 16133 14197 16167
rect 14231 16164 14243 16167
rect 14752 16164 14780 16192
rect 14231 16136 14780 16164
rect 14231 16133 14243 16136
rect 14185 16127 14243 16133
rect 15930 16124 15936 16176
rect 15988 16164 15994 16176
rect 16393 16167 16451 16173
rect 16393 16164 16405 16167
rect 15988 16136 16405 16164
rect 15988 16124 15994 16136
rect 16393 16133 16405 16136
rect 16439 16133 16451 16167
rect 16393 16127 16451 16133
rect 17126 16124 17132 16176
rect 17184 16124 17190 16176
rect 18414 16164 18420 16176
rect 18354 16136 18420 16164
rect 18414 16124 18420 16136
rect 18472 16164 18478 16176
rect 18877 16167 18935 16173
rect 18877 16164 18889 16167
rect 18472 16136 18889 16164
rect 18472 16124 18478 16136
rect 18877 16133 18889 16136
rect 18923 16133 18935 16167
rect 18877 16127 18935 16133
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19705 16167 19763 16173
rect 19705 16164 19717 16167
rect 19392 16136 19717 16164
rect 19392 16124 19398 16136
rect 19705 16133 19717 16136
rect 19751 16133 19763 16167
rect 19705 16127 19763 16133
rect 20990 16124 20996 16176
rect 21048 16164 21054 16176
rect 21269 16167 21327 16173
rect 21269 16164 21281 16167
rect 21048 16136 21281 16164
rect 21048 16124 21054 16136
rect 21269 16133 21281 16136
rect 21315 16133 21327 16167
rect 21269 16127 21327 16133
rect 21634 16124 21640 16176
rect 21692 16164 21698 16176
rect 23216 16164 23244 16195
rect 21692 16136 23244 16164
rect 21692 16124 21698 16136
rect 6638 16056 6644 16108
rect 6696 16056 6702 16108
rect 8404 16068 9536 16096
rect 8404 16040 8432 16068
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 8294 16028 8300 16040
rect 6963 16000 8300 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 8386 15988 8392 16040
rect 8444 15988 8450 16040
rect 9508 16037 9536 16068
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 10468 16068 10517 16096
rect 10468 16056 10474 16068
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12802 16096 12808 16108
rect 12207 16068 12808 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20441 16099 20499 16105
rect 20441 16096 20453 16099
rect 19659 16068 20453 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 20441 16065 20453 16068
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 22370 16056 22376 16108
rect 22428 16056 22434 16108
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22520 16068 23397 16096
rect 22520 16056 22526 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 24118 16056 24124 16108
rect 24176 16056 24182 16108
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9493 16031 9551 16037
rect 9493 15997 9505 16031
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 15997 10747 16031
rect 10689 15991 10747 15997
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2593 15895 2651 15901
rect 2593 15892 2605 15895
rect 1820 15864 2605 15892
rect 1820 15852 1826 15864
rect 2593 15861 2605 15864
rect 2639 15861 2651 15895
rect 9416 15892 9444 15991
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 10704 15960 10732 15991
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 11204 16000 12265 16028
rect 11204 15988 11210 16000
rect 12253 15997 12265 16000
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 15997 19947 16031
rect 22278 16028 22284 16040
rect 19889 15991 19947 15997
rect 20548 16000 22284 16028
rect 10284 15932 10732 15960
rect 19904 15960 19932 15991
rect 20548 15960 20576 16000
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 22554 15988 22560 16040
rect 22612 15988 22618 16040
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 19904 15932 20576 15960
rect 21453 15963 21511 15969
rect 10284 15920 10290 15932
rect 21453 15929 21465 15963
rect 21499 15960 21511 15963
rect 23842 15960 23848 15972
rect 21499 15932 23848 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 23842 15920 23848 15932
rect 23900 15920 23906 15972
rect 12342 15892 12348 15904
rect 9416 15864 12348 15892
rect 2593 15855 2651 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 14090 15852 14096 15904
rect 14148 15892 14154 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 14148 15864 14289 15892
rect 14148 15852 14154 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15804 15864 16037 15892
rect 15804 15852 15810 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 21818 15892 21824 15904
rect 17368 15864 21824 15892
rect 17368 15852 17374 15864
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22005 15895 22063 15901
rect 22005 15892 22017 15895
rect 21968 15864 22017 15892
rect 21968 15852 21974 15864
rect 22005 15861 22017 15864
rect 22051 15861 22063 15895
rect 22005 15855 22063 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 9950 15648 9956 15700
rect 10008 15648 10014 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10284 15660 12388 15688
rect 10284 15648 10290 15660
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11330 15552 11336 15564
rect 11103 15524 11336 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 12360 15552 12388 15660
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 12492 15660 13553 15688
rect 12492 15648 12498 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 14274 15648 14280 15700
rect 14332 15648 14338 15700
rect 17313 15623 17371 15629
rect 17313 15589 17325 15623
rect 17359 15620 17371 15623
rect 19334 15620 19340 15632
rect 17359 15592 19340 15620
rect 17359 15589 17371 15592
rect 17313 15583 17371 15589
rect 19334 15580 19340 15592
rect 19392 15580 19398 15632
rect 14366 15552 14372 15564
rect 12360 15524 14372 15552
rect 14366 15512 14372 15524
rect 14424 15552 14430 15564
rect 14829 15555 14887 15561
rect 14829 15552 14841 15555
rect 14424 15524 14841 15552
rect 14424 15512 14430 15524
rect 14829 15521 14841 15524
rect 14875 15521 14887 15555
rect 14829 15515 14887 15521
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17460 15524 17877 15552
rect 17460 15512 17466 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 20073 15555 20131 15561
rect 20073 15521 20085 15555
rect 20119 15552 20131 15555
rect 21174 15552 21180 15564
rect 20119 15524 21180 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 13446 15444 13452 15496
rect 13504 15444 13510 15496
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15484 14703 15487
rect 15286 15484 15292 15496
rect 14691 15456 15292 15484
rect 14691 15453 14703 15456
rect 14645 15447 14703 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 16390 15444 16396 15496
rect 16448 15484 16454 15496
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 16448 15456 17785 15484
rect 16448 15444 16454 15456
rect 17773 15453 17785 15456
rect 17819 15484 17831 15487
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 17819 15456 18337 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 19242 15484 19248 15496
rect 18748 15456 19248 15484
rect 18748 15444 18754 15456
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 19886 15484 19892 15496
rect 19843 15456 19892 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 19886 15444 19892 15456
rect 19944 15444 19950 15496
rect 20806 15444 20812 15496
rect 20864 15444 20870 15496
rect 22833 15487 22891 15493
rect 22833 15453 22845 15487
rect 22879 15484 22891 15487
rect 24210 15484 24216 15496
rect 22879 15456 24216 15484
rect 22879 15453 22891 15456
rect 22833 15447 22891 15453
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 11333 15419 11391 15425
rect 11333 15385 11345 15419
rect 11379 15385 11391 15419
rect 11333 15379 11391 15385
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 10229 15351 10287 15357
rect 10229 15317 10241 15351
rect 10275 15348 10287 15351
rect 10410 15348 10416 15360
rect 10275 15320 10416 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 10410 15308 10416 15320
rect 10468 15308 10474 15360
rect 10781 15351 10839 15357
rect 10781 15317 10793 15351
rect 10827 15348 10839 15351
rect 10870 15348 10876 15360
rect 10827 15320 10876 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 10870 15308 10876 15320
rect 10928 15348 10934 15360
rect 11348 15348 11376 15379
rect 11790 15376 11796 15428
rect 11848 15376 11854 15428
rect 16758 15376 16764 15428
rect 16816 15416 16822 15428
rect 21085 15419 21143 15425
rect 21085 15416 21097 15419
rect 16816 15388 19932 15416
rect 16816 15376 16822 15388
rect 11698 15348 11704 15360
rect 10928 15320 11704 15348
rect 10928 15308 10934 15320
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12676 15320 12817 15348
rect 12676 15308 12682 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 15654 15348 15660 15360
rect 14783 15320 15660 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 17034 15308 17040 15360
rect 17092 15348 17098 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17092 15320 17693 15348
rect 17092 15308 17098 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 18690 15308 18696 15360
rect 18748 15308 18754 15360
rect 19429 15351 19487 15357
rect 19429 15317 19441 15351
rect 19475 15348 19487 15351
rect 19610 15348 19616 15360
rect 19475 15320 19616 15348
rect 19475 15317 19487 15320
rect 19429 15311 19487 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 19904 15357 19932 15388
rect 20088 15388 21097 15416
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20088 15348 20116 15388
rect 21085 15385 21097 15388
rect 21131 15385 21143 15419
rect 21085 15379 21143 15385
rect 21818 15376 21824 15428
rect 21876 15376 21882 15428
rect 23845 15419 23903 15425
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 26050 15416 26056 15428
rect 23891 15388 26056 15416
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 26050 15376 26056 15388
rect 26108 15376 26114 15428
rect 19935 15320 20116 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 21542 15308 21548 15360
rect 21600 15348 21606 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 21600 15320 21925 15348
rect 21600 15308 21606 15320
rect 21913 15317 21925 15320
rect 21959 15317 21971 15351
rect 21913 15311 21971 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 8812 15116 9536 15144
rect 8812 15104 8818 15116
rect 9398 15036 9404 15088
rect 9456 15036 9462 15088
rect 9508 15076 9536 15116
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12216 15116 13001 15144
rect 12216 15104 12222 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 17310 15144 17316 15156
rect 14231 15116 17316 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18748 15116 18797 15144
rect 18748 15104 18754 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 18874 15104 18880 15156
rect 18932 15104 18938 15156
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22370 15144 22376 15156
rect 22327 15116 22376 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 12526 15076 12532 15088
rect 9508 15048 9890 15076
rect 12406 15048 12532 15076
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9125 14903 9183 14909
rect 9140 14804 9168 14903
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10928 14912 11161 14940
rect 10928 14900 10934 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 9950 14804 9956 14816
rect 9140 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 10560 14776 11529 14804
rect 10560 14764 10566 14776
rect 11517 14773 11529 14776
rect 11563 14804 11575 14807
rect 11790 14804 11796 14816
rect 11563 14776 11796 14804
rect 11563 14773 11575 14776
rect 11517 14767 11575 14773
rect 11790 14764 11796 14776
rect 11848 14804 11854 14816
rect 12406 14804 12434 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 12713 15079 12771 15085
rect 12713 15045 12725 15079
rect 12759 15076 12771 15079
rect 13446 15076 13452 15088
rect 12759 15048 13452 15076
rect 12759 15045 12771 15048
rect 12713 15039 12771 15045
rect 13446 15036 13452 15048
rect 13504 15076 13510 15088
rect 17034 15076 17040 15088
rect 13504 15048 17040 15076
rect 13504 15036 13510 15048
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 17276 15048 17693 15076
rect 17276 15036 17282 15048
rect 17681 15045 17693 15048
rect 17727 15045 17739 15079
rect 17681 15039 17739 15045
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 14645 15011 14703 15017
rect 14645 14977 14657 15011
rect 14691 15008 14703 15011
rect 14691 14980 15332 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13906 14940 13912 14952
rect 13679 14912 13912 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 15304 14949 15332 14980
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 15528 14980 15669 15008
rect 15528 14968 15534 14980
rect 15657 14977 15669 14980
rect 15703 15008 15715 15011
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15703 14980 16129 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 16117 14977 16129 14980
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18656 14980 19012 15008
rect 18656 14968 18662 14980
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 16390 14940 16396 14952
rect 15335 14912 16396 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 18984 14949 19012 14980
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 23937 15011 23995 15017
rect 23937 15008 23949 15011
rect 23716 14980 23949 15008
rect 23716 14968 23722 14980
rect 23937 14977 23949 14980
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14909 19027 14943
rect 18969 14903 19027 14909
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 15841 14875 15899 14881
rect 15841 14841 15853 14875
rect 15887 14872 15899 14875
rect 16666 14872 16672 14884
rect 15887 14844 16672 14872
rect 15887 14841 15899 14844
rect 15841 14835 15899 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 17405 14875 17463 14881
rect 17405 14841 17417 14875
rect 17451 14872 17463 14875
rect 19518 14872 19524 14884
rect 17451 14844 19524 14872
rect 17451 14841 17463 14844
rect 17405 14835 17463 14841
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 11848 14776 12434 14804
rect 18417 14807 18475 14813
rect 11848 14764 11854 14776
rect 18417 14773 18429 14807
rect 18463 14804 18475 14807
rect 19150 14804 19156 14816
rect 18463 14776 19156 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 19794 14804 19800 14816
rect 19659 14776 19800 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 19886 14764 19892 14816
rect 19944 14804 19950 14816
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 19944 14776 20085 14804
rect 19944 14764 19950 14776
rect 20073 14773 20085 14776
rect 20119 14773 20131 14807
rect 20073 14767 20131 14773
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 10836 14572 12434 14600
rect 10836 14560 10842 14572
rect 11330 14492 11336 14544
rect 11388 14492 11394 14544
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 11977 14535 12035 14541
rect 11977 14532 11989 14535
rect 11848 14504 11989 14532
rect 11848 14492 11854 14504
rect 11977 14501 11989 14504
rect 12023 14501 12035 14535
rect 12406 14532 12434 14572
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12860 14572 13001 14600
rect 12860 14560 12866 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 17126 14560 17132 14612
rect 17184 14560 17190 14612
rect 23017 14603 23075 14609
rect 23017 14569 23029 14603
rect 23063 14600 23075 14603
rect 23382 14600 23388 14612
rect 23063 14572 23388 14600
rect 23063 14569 23075 14572
rect 23017 14563 23075 14569
rect 14093 14535 14151 14541
rect 14093 14532 14105 14535
rect 12406 14504 14105 14532
rect 11977 14495 12035 14501
rect 14093 14501 14105 14504
rect 14139 14532 14151 14535
rect 14550 14532 14556 14544
rect 14139 14504 14556 14532
rect 14139 14501 14151 14504
rect 14093 14495 14151 14501
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 16942 14492 16948 14544
rect 17000 14532 17006 14544
rect 20806 14532 20812 14544
rect 17000 14504 20812 14532
rect 17000 14492 17006 14504
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11348 14464 11376 14492
rect 10008 14436 11376 14464
rect 10008 14424 10014 14436
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 13446 14464 13452 14476
rect 12584 14436 13452 14464
rect 12584 14424 12590 14436
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 14734 14464 14740 14476
rect 13679 14436 14740 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 13648 14396 13676 14427
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16390 14464 16396 14476
rect 15436 14436 16396 14464
rect 15436 14424 15442 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 12759 14368 13676 14396
rect 18233 14399 18291 14405
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18506 14396 18512 14408
rect 18279 14368 18512 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18564 14368 18613 14396
rect 18564 14356 18570 14368
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14396 19487 14399
rect 20070 14396 20076 14408
rect 19475 14368 20076 14396
rect 19475 14365 19487 14368
rect 19429 14359 19487 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20898 14356 20904 14408
rect 20956 14356 20962 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 23032 14396 23060 14563
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 22336 14368 23060 14396
rect 22336 14356 22342 14368
rect 10226 14288 10232 14340
rect 10284 14288 10290 14340
rect 10502 14288 10508 14340
rect 10560 14328 10566 14340
rect 10560 14300 10718 14328
rect 10560 14288 10566 14300
rect 13354 14288 13360 14340
rect 13412 14288 13418 14340
rect 15657 14331 15715 14337
rect 15657 14297 15669 14331
rect 15703 14328 15715 14331
rect 15930 14328 15936 14340
rect 15703 14300 15936 14328
rect 15703 14297 15715 14300
rect 15657 14291 15715 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 18785 14331 18843 14337
rect 16882 14300 17540 14328
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10962 14260 10968 14272
rect 9916 14232 10968 14260
rect 9916 14220 9922 14232
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 11020 14232 11713 14260
rect 11020 14220 11026 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 13372 14260 13400 14288
rect 14369 14263 14427 14269
rect 14369 14260 14381 14263
rect 13372 14232 14381 14260
rect 11701 14223 11759 14229
rect 14369 14229 14381 14232
rect 14415 14260 14427 14263
rect 14553 14263 14611 14269
rect 14553 14260 14565 14263
rect 14415 14232 14565 14260
rect 14415 14229 14427 14232
rect 14369 14223 14427 14229
rect 14553 14229 14565 14232
rect 14599 14260 14611 14263
rect 15562 14260 15568 14272
rect 14599 14232 15568 14260
rect 14599 14229 14611 14232
rect 14553 14223 14611 14229
rect 15562 14220 15568 14232
rect 15620 14260 15626 14272
rect 16390 14260 16396 14272
rect 15620 14232 16396 14260
rect 15620 14220 15626 14232
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16960 14260 16988 14300
rect 17512 14269 17540 14300
rect 18785 14297 18797 14331
rect 18831 14328 18843 14331
rect 21174 14328 21180 14340
rect 18831 14300 21180 14328
rect 18831 14297 18843 14300
rect 18785 14291 18843 14297
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 16540 14232 16988 14260
rect 17497 14263 17555 14269
rect 16540 14220 16546 14232
rect 17497 14229 17509 14263
rect 17543 14260 17555 14263
rect 18414 14260 18420 14272
rect 17543 14232 18420 14260
rect 17543 14229 17555 14232
rect 17497 14223 17555 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 18966 14260 18972 14272
rect 18564 14232 18972 14260
rect 18564 14220 18570 14232
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19978 14220 19984 14272
rect 20036 14220 20042 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22649 14263 22707 14269
rect 22649 14260 22661 14263
rect 21876 14232 22661 14260
rect 21876 14220 21882 14232
rect 22649 14229 22661 14232
rect 22695 14229 22707 14263
rect 22649 14223 22707 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 9950 14056 9956 14068
rect 8128 14028 9956 14056
rect 8128 13988 8156 14028
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12299 14028 13124 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 8036 13960 8156 13988
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 8036 13929 8064 13960
rect 8754 13948 8760 14000
rect 8812 13948 8818 14000
rect 11882 13948 11888 14000
rect 11940 13948 11946 14000
rect 13096 13988 13124 14028
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13596 14028 13645 14056
rect 13596 14016 13602 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 18322 14016 18328 14068
rect 18380 14056 18386 14068
rect 18874 14056 18880 14068
rect 18380 14028 18880 14056
rect 18380 14016 18386 14028
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21140 14028 21833 14056
rect 21140 14016 21146 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 21821 14019 21879 14025
rect 23017 14059 23075 14065
rect 23017 14025 23029 14059
rect 23063 14056 23075 14059
rect 23382 14056 23388 14068
rect 23063 14028 23388 14056
rect 23063 14025 23075 14028
rect 23017 14019 23075 14025
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 15286 13988 15292 14000
rect 12544 13960 12848 13988
rect 13096 13960 15292 13988
rect 8021 13923 8079 13929
rect 8021 13889 8033 13923
rect 8067 13889 8079 13923
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 8021 13883 8079 13889
rect 9324 13892 10057 13920
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9324 13852 9352 13892
rect 10045 13889 10057 13892
rect 10091 13920 10103 13923
rect 10226 13920 10232 13932
rect 10091 13892 10232 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10502 13920 10508 13932
rect 10284 13892 10508 13920
rect 10284 13880 10290 13892
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 11900 13920 11928 13948
rect 12544 13920 12572 13960
rect 11900 13892 12572 13920
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 12820 13920 12848 13960
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 17402 13948 17408 14000
rect 17460 13948 17466 14000
rect 19889 13991 19947 13997
rect 18432 13932 18460 13974
rect 19889 13957 19901 13991
rect 19935 13988 19947 13991
rect 21361 13991 21419 13997
rect 19935 13960 21312 13988
rect 19935 13957 19947 13960
rect 19889 13951 19947 13957
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12820 13892 13553 13920
rect 12621 13883 12679 13889
rect 13541 13889 13553 13892
rect 13587 13920 13599 13923
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13587 13892 14013 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 8812 13824 9352 13852
rect 8812 13812 8818 13824
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 9548 13824 9781 13852
rect 9548 13812 9554 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 10468 13824 11897 13852
rect 10468 13812 10474 13824
rect 11885 13821 11897 13824
rect 11931 13852 11943 13855
rect 12636 13852 12664 13883
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 17126 13920 17132 13932
rect 16632 13892 17132 13920
rect 16632 13880 16638 13892
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 18414 13880 18420 13932
rect 18472 13880 18478 13932
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13920 19763 13923
rect 19978 13920 19984 13932
rect 19751 13892 19984 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 20438 13880 20444 13932
rect 20496 13880 20502 13932
rect 21082 13880 21088 13932
rect 21140 13920 21146 13932
rect 21177 13923 21235 13929
rect 21177 13920 21189 13923
rect 21140 13892 21189 13920
rect 21140 13880 21146 13892
rect 21177 13889 21189 13892
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 11931 13824 12664 13852
rect 12713 13855 12771 13861
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 12802 13852 12808 13864
rect 12759 13824 12808 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 18432 13852 18460 13880
rect 18966 13852 18972 13864
rect 18432 13824 18972 13852
rect 12897 13815 12955 13821
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 11848 13756 12434 13784
rect 11848 13744 11854 13756
rect 8284 13719 8342 13725
rect 8284 13685 8296 13719
rect 8330 13716 8342 13719
rect 9858 13716 9864 13728
rect 8330 13688 9864 13716
rect 8330 13685 8342 13688
rect 8284 13679 8342 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 12406 13716 12434 13756
rect 12912 13716 12940 13815
rect 18966 13812 18972 13824
rect 19024 13852 19030 13864
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 19024 13824 19257 13852
rect 19024 13812 19030 13824
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20404 13824 20637 13852
rect 20404 13812 20410 13824
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 21284 13784 21312 13960
rect 21361 13957 21373 13991
rect 21407 13988 21419 13991
rect 21726 13988 21732 14000
rect 21407 13960 21732 13988
rect 21407 13957 21419 13960
rect 21361 13951 21419 13957
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 22738 13948 22744 14000
rect 22796 13988 22802 14000
rect 22796 13960 23980 13988
rect 22796 13948 22802 13960
rect 21450 13880 21456 13932
rect 21508 13920 21514 13932
rect 23952 13929 23980 13960
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 21508 13892 23213 13920
rect 21508 13880 21514 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 23750 13852 23756 13864
rect 21416 13824 23756 13852
rect 21416 13812 21422 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 22186 13784 22192 13796
rect 21284 13756 22192 13784
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 12406 13688 12940 13716
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 7098 13521 7104 13524
rect 7088 13515 7104 13521
rect 7088 13481 7100 13515
rect 7156 13512 7162 13524
rect 7558 13512 7564 13524
rect 7156 13484 7564 13512
rect 7088 13475 7104 13481
rect 7098 13472 7104 13475
rect 7156 13472 7162 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8812 13484 8953 13512
rect 8812 13472 8818 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 11606 13472 11612 13524
rect 11664 13472 11670 13524
rect 12342 13472 12348 13524
rect 12400 13472 12406 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 12860 13484 13369 13512
rect 12860 13472 12866 13484
rect 13357 13481 13369 13484
rect 13403 13512 13415 13515
rect 13403 13484 15884 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 13262 13444 13268 13456
rect 12406 13416 13268 13444
rect 8478 13376 8484 13388
rect 6840 13348 8484 13376
rect 6840 13320 6868 13348
rect 8478 13336 8484 13348
rect 8536 13376 8542 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 8536 13348 9137 13376
rect 8536 13336 8542 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 8386 13308 8392 13320
rect 8234 13280 8392 13308
rect 8386 13268 8392 13280
rect 8444 13308 8450 13320
rect 8754 13308 8760 13320
rect 8444 13280 8760 13308
rect 8444 13268 8450 13280
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 10137 13243 10195 13249
rect 10137 13240 10149 13243
rect 8404 13212 10149 13240
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 8404 13172 8432 13212
rect 10137 13209 10149 13212
rect 10183 13209 10195 13243
rect 10137 13203 10195 13209
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 10594 13240 10600 13252
rect 10284 13212 10600 13240
rect 10284 13200 10290 13212
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 5868 13144 8432 13172
rect 8573 13175 8631 13181
rect 5868 13132 5874 13144
rect 8573 13141 8585 13175
rect 8619 13172 8631 13175
rect 8754 13172 8760 13184
rect 8619 13144 8760 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11977 13175 12035 13181
rect 11977 13172 11989 13175
rect 11572 13144 11989 13172
rect 11572 13132 11578 13144
rect 11977 13141 11989 13144
rect 12023 13172 12035 13175
rect 12406 13172 12434 13416
rect 13262 13404 13268 13416
rect 13320 13404 13326 13456
rect 12618 13336 12624 13388
rect 12676 13376 12682 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12676 13348 12909 13376
rect 12676 13336 12682 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15378 13376 15384 13388
rect 14599 13348 15384 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15856 13376 15884 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15988 13484 16313 13512
rect 15988 13472 15994 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 18874 13472 18880 13524
rect 18932 13512 18938 13524
rect 18932 13484 20116 13512
rect 18932 13472 18938 13484
rect 18785 13447 18843 13453
rect 18785 13444 18797 13447
rect 18248 13416 18797 13444
rect 18248 13385 18276 13416
rect 18785 13413 18797 13416
rect 18831 13413 18843 13447
rect 18785 13407 18843 13413
rect 19426 13404 19432 13456
rect 19484 13404 19490 13456
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 15856 13348 18245 13376
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18417 13379 18475 13385
rect 18417 13345 18429 13379
rect 18463 13376 18475 13379
rect 18506 13376 18512 13388
rect 18463 13348 18512 13376
rect 18463 13345 18475 13348
rect 18417 13339 18475 13345
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 20088 13385 20116 13484
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20717 13515 20775 13521
rect 20717 13512 20729 13515
rect 20496 13484 20729 13512
rect 20496 13472 20502 13484
rect 20717 13481 20729 13484
rect 20763 13481 20775 13515
rect 20717 13475 20775 13481
rect 20073 13379 20131 13385
rect 18564 13348 19932 13376
rect 18564 13336 18570 13348
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 14458 13308 14464 13320
rect 12759 13280 14464 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 16172 13280 17509 13308
rect 16172 13268 16178 13280
rect 17497 13277 17509 13280
rect 17543 13308 17555 13311
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 17543 13280 18153 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19904 13308 19932 13348
rect 20073 13345 20085 13379
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 21450 13308 21456 13320
rect 19904 13280 21456 13308
rect 19797 13271 19855 13277
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 14366 13240 14372 13252
rect 12851 13212 14372 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 14550 13200 14556 13252
rect 14608 13240 14614 13252
rect 14826 13240 14832 13252
rect 14608 13212 14832 13240
rect 14608 13200 14614 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 16206 13240 16212 13252
rect 16054 13212 16212 13240
rect 16206 13200 16212 13212
rect 16264 13240 16270 13252
rect 16482 13240 16488 13252
rect 16264 13212 16488 13240
rect 16264 13200 16270 13212
rect 16482 13200 16488 13212
rect 16540 13200 16546 13252
rect 19812 13240 19840 13271
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 20070 13240 20076 13252
rect 19812 13212 20076 13240
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 25130 13240 25136 13252
rect 23891 13212 25136 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 12023 13144 12434 13172
rect 16853 13175 16911 13181
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 16853 13141 16865 13175
rect 16899 13172 16911 13175
rect 17218 13172 17224 13184
rect 16899 13144 17224 13172
rect 16899 13141 16911 13144
rect 16853 13135 16911 13141
rect 17218 13132 17224 13144
rect 17276 13132 17282 13184
rect 17773 13175 17831 13181
rect 17773 13141 17785 13175
rect 17819 13172 17831 13175
rect 18874 13172 18880 13184
rect 17819 13144 18880 13172
rect 17819 13141 17831 13144
rect 17773 13135 17831 13141
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19889 13175 19947 13181
rect 19889 13172 19901 13175
rect 19392 13144 19901 13172
rect 19392 13132 19398 13144
rect 19889 13141 19901 13144
rect 19935 13141 19947 13175
rect 19889 13135 19947 13141
rect 21637 13175 21695 13181
rect 21637 13141 21649 13175
rect 21683 13172 21695 13175
rect 22278 13172 22284 13184
rect 21683 13144 22284 13172
rect 21683 13141 21695 13144
rect 21637 13135 21695 13141
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 8386 12968 8392 12980
rect 6696 12940 8392 12968
rect 6696 12928 6702 12940
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8662 12928 8668 12980
rect 8720 12928 8726 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 11149 12971 11207 12977
rect 10652 12940 11008 12968
rect 10652 12928 10658 12940
rect 9674 12900 9680 12912
rect 9416 12872 9680 12900
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 6604 12804 8585 12832
rect 6604 12792 6610 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 8662 12792 8668 12844
rect 8720 12832 8726 12844
rect 8846 12832 8852 12844
rect 8720 12804 8852 12832
rect 8720 12792 8726 12804
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9416 12841 9444 12872
rect 9674 12860 9680 12872
rect 9732 12900 9738 12912
rect 9950 12900 9956 12912
rect 9732 12872 9956 12900
rect 9732 12860 9738 12872
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 10226 12860 10232 12912
rect 10284 12860 10290 12912
rect 10980 12900 11008 12940
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11790 12968 11796 12980
rect 11195 12940 11796 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13262 12928 13268 12980
rect 13320 12928 13326 12980
rect 14918 12928 14924 12980
rect 14976 12928 14982 12980
rect 16114 12928 16120 12980
rect 16172 12928 16178 12980
rect 16482 12928 16488 12980
rect 16540 12928 16546 12980
rect 17218 12928 17224 12980
rect 17276 12928 17282 12980
rect 17310 12928 17316 12980
rect 17368 12928 17374 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 18524 12940 19073 12968
rect 11514 12900 11520 12912
rect 10980 12872 11520 12900
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 14461 12903 14519 12909
rect 14461 12869 14473 12903
rect 14507 12900 14519 12903
rect 14936 12900 14964 12928
rect 14507 12872 14964 12900
rect 14507 12869 14519 12872
rect 14461 12863 14519 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 18524 12909 18552 12940
rect 19061 12937 19073 12940
rect 19107 12968 19119 12971
rect 19242 12968 19248 12980
rect 19107 12940 19248 12968
rect 19107 12937 19119 12940
rect 19061 12931 19119 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 20898 12968 20904 12980
rect 19720 12940 20904 12968
rect 15381 12903 15439 12909
rect 15381 12900 15393 12903
rect 15252 12872 15393 12900
rect 15252 12860 15258 12872
rect 15381 12869 15393 12872
rect 15427 12900 15439 12903
rect 15841 12903 15899 12909
rect 15841 12900 15853 12903
rect 15427 12872 15853 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15841 12869 15853 12872
rect 15887 12869 15899 12903
rect 15841 12863 15899 12869
rect 18509 12903 18567 12909
rect 18509 12869 18521 12903
rect 18555 12869 18567 12903
rect 18509 12863 18567 12869
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13688 12804 13737 12832
rect 13688 12792 13694 12804
rect 13725 12801 13737 12804
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 15988 12804 17448 12832
rect 15988 12792 15994 12804
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 8812 12736 9689 12764
rect 8812 12724 8818 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 14826 12764 14832 12776
rect 9677 12727 9735 12733
rect 10704 12736 14832 12764
rect 8205 12631 8263 12637
rect 8205 12597 8217 12631
rect 8251 12628 8263 12631
rect 10704 12628 10732 12736
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 17420 12773 17448 12804
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 19518 12832 19524 12844
rect 18932 12804 19524 12832
rect 18932 12792 18938 12804
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 19720 12773 19748 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21450 12928 21456 12980
rect 21508 12928 21514 12980
rect 22278 12900 22284 12912
rect 21206 12872 22284 12900
rect 22278 12860 22284 12872
rect 22336 12900 22342 12912
rect 22646 12900 22652 12912
rect 22336 12872 22652 12900
rect 22336 12860 22342 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22833 12835 22891 12841
rect 22833 12832 22845 12835
rect 22152 12804 22845 12832
rect 22152 12792 22158 12804
rect 22833 12801 22845 12804
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23348 12804 23949 12832
rect 23348 12792 23354 12804
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 19705 12767 19763 12773
rect 19705 12764 19717 12767
rect 18380 12736 19717 12764
rect 18380 12724 18386 12736
rect 19705 12733 19717 12736
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 21818 12764 21824 12776
rect 20027 12736 21824 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 21818 12724 21824 12736
rect 21876 12724 21882 12776
rect 22002 12724 22008 12776
rect 22060 12724 22066 12776
rect 24762 12724 24768 12776
rect 24820 12724 24826 12776
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 14274 12696 14280 12708
rect 13955 12668 14280 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14642 12656 14648 12708
rect 14700 12656 14706 12708
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 16899 12668 19840 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 8251 12600 10732 12628
rect 15473 12631 15531 12637
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 15473 12597 15485 12631
rect 15519 12628 15531 12631
rect 16298 12628 16304 12640
rect 15519 12600 16304 12628
rect 15519 12597 15531 12600
rect 15473 12591 15531 12597
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 18598 12588 18604 12640
rect 18656 12588 18662 12640
rect 19812 12628 19840 12668
rect 20530 12628 20536 12640
rect 19812 12600 20536 12628
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22612 12600 22661 12628
rect 22612 12588 22618 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 8662 12424 8668 12436
rect 2740 12396 8668 12424
rect 2740 12384 2746 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 10928 12396 12848 12424
rect 10928 12384 10934 12396
rect 12820 12356 12848 12396
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13872 12396 14105 12424
rect 13872 12384 13878 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 14093 12387 14151 12393
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 17402 12424 17408 12436
rect 16040 12396 17408 12424
rect 12820 12328 13952 12356
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10962 12288 10968 12300
rect 9732 12260 10968 12288
rect 9732 12248 9738 12260
rect 10962 12248 10968 12260
rect 11020 12288 11026 12300
rect 11517 12291 11575 12297
rect 11517 12288 11529 12291
rect 11020 12260 11529 12288
rect 11020 12248 11026 12260
rect 11517 12257 11529 12260
rect 11563 12257 11575 12291
rect 11517 12251 11575 12257
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 13924 12297 13952 12328
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 13955 12260 15117 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 15105 12257 15117 12260
rect 15151 12288 15163 12291
rect 15930 12288 15936 12300
rect 15151 12260 15936 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 13688 12192 13737 12220
rect 13688 12180 13694 12192
rect 13725 12189 13737 12192
rect 13771 12220 13783 12223
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 13771 12192 14933 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14921 12189 14933 12192
rect 14967 12220 14979 12223
rect 15838 12220 15844 12232
rect 14967 12192 15844 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 16040 12229 16068 12396
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 17552 12396 18889 12424
rect 17552 12384 17558 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 19610 12316 19616 12368
rect 19668 12356 19674 12368
rect 21085 12359 21143 12365
rect 19668 12328 20576 12356
rect 19668 12316 19674 12328
rect 16206 12248 16212 12300
rect 16264 12248 16270 12300
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 17405 12291 17463 12297
rect 17405 12257 17417 12291
rect 17451 12288 17463 12291
rect 19978 12288 19984 12300
rect 17451 12260 19984 12288
rect 17451 12257 17463 12260
rect 17405 12251 17463 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 20548 12288 20576 12328
rect 21085 12325 21097 12359
rect 21131 12356 21143 12359
rect 22830 12356 22836 12368
rect 21131 12328 22836 12356
rect 21131 12325 21143 12328
rect 21085 12319 21143 12325
rect 22830 12316 22836 12328
rect 22888 12316 22894 12368
rect 21545 12291 21603 12297
rect 21545 12288 21557 12291
rect 20548 12260 21557 12288
rect 21545 12257 21557 12260
rect 21591 12257 21603 12291
rect 21545 12251 21603 12257
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12288 21787 12291
rect 21818 12288 21824 12300
rect 21775 12260 21824 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 21968 12260 23428 12288
rect 21968 12248 21974 12260
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 18966 12220 18972 12232
rect 18538 12192 18972 12220
rect 16025 12183 16083 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 19208 12192 20637 12220
rect 19208 12180 19214 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12220 21511 12223
rect 22002 12220 22008 12232
rect 21499 12192 22008 12220
rect 21499 12189 21511 12192
rect 21453 12183 21511 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 23400 12229 23428 12260
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 13446 12152 13452 12164
rect 13018 12124 13452 12152
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 14829 12155 14887 12161
rect 14829 12121 14841 12155
rect 14875 12152 14887 12155
rect 16850 12152 16856 12164
rect 14875 12124 16856 12152
rect 14875 12121 14887 12124
rect 14829 12115 14887 12121
rect 16850 12112 16856 12124
rect 16908 12152 16914 12164
rect 17310 12152 17316 12164
rect 16908 12124 17316 12152
rect 16908 12112 16914 12124
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 19794 12152 19800 12164
rect 18708 12124 19800 12152
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13265 12087 13323 12093
rect 13265 12084 13277 12087
rect 13228 12056 13277 12084
rect 13228 12044 13234 12056
rect 13265 12053 13277 12056
rect 13311 12053 13323 12087
rect 13265 12047 13323 12053
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 16022 12084 16028 12096
rect 15436 12056 16028 12084
rect 15436 12044 15442 12056
rect 16022 12044 16028 12056
rect 16080 12084 16086 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 16080 12056 16129 12084
rect 16080 12044 16086 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 18708 12084 18736 12124
rect 19794 12112 19800 12124
rect 19852 12112 19858 12164
rect 22738 12152 22744 12164
rect 20456 12124 22744 12152
rect 17460 12056 18736 12084
rect 17460 12044 17466 12056
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19242 12084 19248 12096
rect 19024 12056 19248 12084
rect 19024 12044 19030 12056
rect 19242 12044 19248 12056
rect 19300 12084 19306 12096
rect 20456 12093 20484 12124
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 19337 12087 19395 12093
rect 19337 12084 19349 12087
rect 19300 12056 19349 12084
rect 19300 12044 19306 12056
rect 19337 12053 19349 12056
rect 19383 12053 19395 12087
rect 19337 12047 19395 12053
rect 20441 12087 20499 12093
rect 20441 12053 20453 12087
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 24118 12084 24124 12096
rect 23247 12056 24124 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13504 11852 14412 11880
rect 13504 11840 13510 11852
rect 14384 11812 14412 11852
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15473 11883 15531 11889
rect 15473 11880 15485 11883
rect 15252 11852 15485 11880
rect 15252 11840 15258 11852
rect 15473 11849 15485 11852
rect 15519 11849 15531 11883
rect 15473 11843 15531 11849
rect 16114 11840 16120 11892
rect 16172 11840 16178 11892
rect 17494 11840 17500 11892
rect 17552 11840 17558 11892
rect 18322 11880 18328 11892
rect 18248 11852 18328 11880
rect 16132 11812 16160 11840
rect 14306 11784 16160 11812
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 17512 11812 17540 11840
rect 16991 11784 17540 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 10962 11704 10968 11756
rect 11020 11744 11026 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 11020 11716 12817 11744
rect 11020 11704 11026 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 18248 11753 18276 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19300 11852 19840 11880
rect 19300 11840 19306 11852
rect 18506 11772 18512 11824
rect 18564 11772 18570 11824
rect 19812 11812 19840 11852
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 22646 11880 22652 11892
rect 20395 11852 22652 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 20364 11812 20392 11843
rect 22646 11840 22652 11852
rect 22704 11880 22710 11892
rect 24213 11883 24271 11889
rect 24213 11880 24225 11883
rect 22704 11852 24225 11880
rect 22704 11840 22710 11852
rect 24213 11849 24225 11852
rect 24259 11849 24271 11883
rect 24213 11843 24271 11849
rect 19734 11784 20392 11812
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 20901 11815 20959 11821
rect 20901 11812 20913 11815
rect 20864 11784 20913 11812
rect 20864 11772 20870 11784
rect 20901 11781 20913 11784
rect 20947 11812 20959 11815
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 20947 11784 21373 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14792 11716 15393 11744
rect 14792 11704 14798 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 18233 11747 18291 11753
rect 18233 11713 18245 11747
rect 18279 11713 18291 11747
rect 18233 11707 18291 11713
rect 22370 11704 22376 11756
rect 22428 11744 22434 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22428 11716 22937 11744
rect 22428 11704 22434 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13170 11676 13176 11688
rect 13127 11648 13176 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13170 11636 13176 11648
rect 13228 11676 13234 11688
rect 15565 11679 15623 11685
rect 13228 11648 14136 11676
rect 13228 11636 13234 11648
rect 14108 11608 14136 11648
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15565 11639 15623 11645
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21358 11676 21364 11688
rect 21131 11648 21364 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 15580 11608 15608 11639
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 14108 11580 15608 11608
rect 15013 11543 15071 11549
rect 15013 11509 15025 11543
rect 15059 11540 15071 11543
rect 15746 11540 15752 11552
rect 15059 11512 15752 11540
rect 15059 11509 15071 11512
rect 15013 11503 15071 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 17037 11543 17095 11549
rect 17037 11540 17049 11543
rect 16908 11512 17049 11540
rect 16908 11500 16914 11512
rect 17037 11509 17049 11512
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 14366 11296 14372 11348
rect 14424 11336 14430 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14424 11308 15485 11336
rect 14424 11296 14430 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 14734 11160 14740 11212
rect 14792 11160 14798 11212
rect 16022 11160 16028 11212
rect 16080 11160 16086 11212
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 19886 11132 19892 11144
rect 15988 11104 19892 11132
rect 15988 11092 15994 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 5902 11024 5908 11076
rect 5960 11064 5966 11076
rect 10134 11064 10140 11076
rect 5960 11036 10140 11064
rect 5960 11024 5966 11036
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 15841 11067 15899 11073
rect 15841 11033 15853 11067
rect 15887 11064 15899 11067
rect 20622 11064 20628 11076
rect 15887 11036 20628 11064
rect 15887 11033 15899 11036
rect 15841 11027 15899 11033
rect 20622 11024 20628 11036
rect 20680 11024 20686 11076
rect 20806 11024 20812 11076
rect 20864 11024 20870 11076
rect 20993 11067 21051 11073
rect 20993 11033 21005 11067
rect 21039 11064 21051 11067
rect 23934 11064 23940 11076
rect 21039 11036 23940 11064
rect 21039 11033 21051 11036
rect 20993 11027 21051 11033
rect 23934 11024 23940 11036
rect 23992 11024 23998 11076
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 19610 10956 19616 11008
rect 19668 10956 19674 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 14645 10795 14703 10801
rect 14645 10761 14657 10795
rect 14691 10792 14703 10795
rect 19521 10795 19579 10801
rect 14691 10764 16574 10792
rect 14691 10761 14703 10764
rect 14645 10755 14703 10761
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 12069 10727 12127 10733
rect 12069 10724 12081 10727
rect 10100 10696 12081 10724
rect 10100 10684 10106 10696
rect 12069 10693 12081 10696
rect 12115 10724 12127 10727
rect 12529 10727 12587 10733
rect 12529 10724 12541 10727
rect 12115 10696 12541 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 12529 10693 12541 10696
rect 12575 10693 12587 10727
rect 12529 10687 12587 10693
rect 15381 10727 15439 10733
rect 15381 10693 15393 10727
rect 15427 10724 15439 10727
rect 16022 10724 16028 10736
rect 15427 10696 16028 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 16022 10684 16028 10696
rect 16080 10684 16086 10736
rect 16546 10724 16574 10764
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19610 10792 19616 10804
rect 19567 10764 19616 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20349 10795 20407 10801
rect 20349 10761 20361 10795
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 20364 10724 20392 10755
rect 16546 10696 19840 10724
rect 20364 10696 23428 10724
rect 14826 10616 14832 10668
rect 14884 10616 14890 10668
rect 15746 10616 15752 10668
rect 15804 10656 15810 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 15804 10628 18429 10656
rect 15804 10616 15810 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 19518 10616 19524 10668
rect 19576 10656 19582 10668
rect 19613 10659 19671 10665
rect 19613 10656 19625 10659
rect 19576 10628 19625 10656
rect 19576 10616 19582 10628
rect 19613 10625 19625 10628
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10557 19763 10591
rect 19812 10588 19840 10696
rect 20530 10616 20536 10668
rect 20588 10616 20594 10668
rect 23400 10665 23428 10696
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23900 10628 23949 10656
rect 23900 10616 23906 10628
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 20806 10588 20812 10600
rect 19812 10560 20812 10588
rect 19705 10551 19763 10557
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12802 10520 12808 10532
rect 12299 10492 12808 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 15197 10523 15255 10529
rect 15197 10489 15209 10523
rect 15243 10520 15255 10523
rect 15930 10520 15936 10532
rect 15243 10492 15936 10520
rect 15243 10489 15255 10492
rect 15197 10483 15255 10489
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 19720 10520 19748 10551
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 24762 10548 24768 10600
rect 24820 10548 24826 10600
rect 19978 10520 19984 10532
rect 19720 10492 19984 10520
rect 19978 10480 19984 10492
rect 20036 10480 20042 10532
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 20622 10452 20628 10464
rect 19199 10424 20628 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 23290 10452 23296 10464
rect 23247 10424 23296 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 23290 10412 23296 10424
rect 23348 10412 23354 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 21269 10183 21327 10189
rect 21269 10149 21281 10183
rect 21315 10180 21327 10183
rect 22462 10180 22468 10192
rect 21315 10152 22468 10180
rect 21315 10149 21327 10152
rect 21269 10143 21327 10149
rect 22462 10140 22468 10152
rect 22520 10140 22526 10192
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18288 10084 22232 10112
rect 18288 10072 18294 10084
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13412 10016 14657 10044
rect 13412 10004 13418 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10044 14887 10047
rect 19426 10044 19432 10056
rect 14875 10016 19432 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 22204 10053 22232 10084
rect 21453 10047 21511 10053
rect 21453 10044 21465 10047
rect 21324 10016 21465 10044
rect 21324 10004 21330 10016
rect 21453 10013 21465 10016
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24946 10044 24952 10056
rect 23891 10016 24952 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 16761 9979 16819 9985
rect 16761 9945 16773 9979
rect 16807 9945 16819 9979
rect 16761 9939 16819 9945
rect 16776 9908 16804 9939
rect 16942 9936 16948 9988
rect 17000 9936 17006 9988
rect 22664 9976 22692 10007
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 22020 9948 22692 9976
rect 18782 9908 18788 9920
rect 16776 9880 18788 9908
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 22020 9917 22048 9948
rect 22738 9936 22744 9988
rect 22796 9976 22802 9988
rect 24673 9979 24731 9985
rect 24673 9976 24685 9979
rect 22796 9948 24685 9976
rect 22796 9936 22802 9948
rect 24673 9945 24685 9948
rect 24719 9945 24731 9979
rect 24673 9939 24731 9945
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 24084 9880 24777 9908
rect 24084 9868 24090 9880
rect 24765 9877 24777 9880
rect 24811 9877 24823 9911
rect 24765 9871 24823 9877
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16448 9608 16957 9636
rect 16448 9596 16454 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 17770 9596 17776 9648
rect 17828 9636 17834 9648
rect 18690 9636 18696 9648
rect 17828 9608 18696 9636
rect 17828 9596 17834 9608
rect 18690 9596 18696 9608
rect 18748 9596 18754 9648
rect 21542 9596 21548 9648
rect 21600 9636 21606 9648
rect 21600 9608 23980 9636
rect 21600 9596 21606 9608
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 5859 9540 6929 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 18472 9540 19257 9568
rect 18472 9528 18478 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 22830 9528 22836 9580
rect 22888 9568 22894 9580
rect 23952 9577 23980 9608
rect 22925 9571 22983 9577
rect 22925 9568 22937 9571
rect 22888 9540 22937 9568
rect 22888 9528 22894 9540
rect 22925 9537 22937 9540
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 4304 9472 7021 9500
rect 4304 9460 4310 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 24670 9460 24676 9512
rect 24728 9460 24734 9512
rect 6546 9392 6552 9444
rect 6604 9392 6610 9444
rect 17129 9435 17187 9441
rect 17129 9401 17141 9435
rect 17175 9432 17187 9435
rect 17586 9432 17592 9444
rect 17175 9404 17592 9432
rect 17175 9401 17187 9404
rect 17129 9395 17187 9401
rect 17586 9392 17592 9404
rect 17644 9392 17650 9444
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 19061 9367 19119 9373
rect 19061 9364 19073 9367
rect 17736 9336 19073 9364
rect 17736 9324 17742 9336
rect 19061 9333 19073 9336
rect 19107 9333 19119 9367
rect 19061 9327 19119 9333
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 22741 9367 22799 9373
rect 22741 9364 22753 9367
rect 22336 9336 22753 9364
rect 22336 9324 22342 9336
rect 22741 9333 22753 9336
rect 22787 9333 22799 9367
rect 22741 9327 22799 9333
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 5534 9160 5540 9172
rect 4120 9132 5540 9160
rect 4120 9120 4126 9132
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 22646 9052 22652 9104
rect 22704 9092 22710 9104
rect 24673 9095 24731 9101
rect 24673 9092 24685 9095
rect 22704 9064 24685 9092
rect 22704 9052 22710 9064
rect 24673 9061 24685 9064
rect 24719 9061 24731 9095
rect 24673 9055 24731 9061
rect 22554 8984 22560 9036
rect 22612 9024 22618 9036
rect 22612 8996 24900 9024
rect 22612 8984 22618 8996
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 20680 8928 21741 8956
rect 20680 8916 20686 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 23382 8916 23388 8968
rect 23440 8956 23446 8968
rect 24872 8965 24900 8996
rect 23937 8959 23995 8965
rect 23937 8956 23949 8959
rect 23440 8928 23949 8956
rect 23440 8916 23446 8928
rect 23937 8925 23949 8928
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8925 24915 8959
rect 24857 8919 24915 8925
rect 21545 8823 21603 8829
rect 21545 8789 21557 8823
rect 21591 8820 21603 8823
rect 22830 8820 22836 8832
rect 21591 8792 22836 8820
rect 21591 8789 21603 8792
rect 21545 8783 21603 8789
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 23474 8780 23480 8832
rect 23532 8820 23538 8832
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23532 8792 23765 8820
rect 23532 8780 23538 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19058 8508 19064 8560
rect 19116 8548 19122 8560
rect 19153 8551 19211 8557
rect 19153 8548 19165 8551
rect 19116 8520 19165 8548
rect 19116 8508 19122 8520
rect 19153 8517 19165 8520
rect 19199 8548 19211 8551
rect 19613 8551 19671 8557
rect 19613 8548 19625 8551
rect 19199 8520 19625 8548
rect 19199 8517 19211 8520
rect 19153 8511 19211 8517
rect 19613 8517 19625 8520
rect 19659 8517 19671 8551
rect 19613 8511 19671 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 21634 8548 21640 8560
rect 20763 8520 21640 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 13906 8412 13912 8424
rect 10100 8384 13912 8412
rect 10100 8372 10106 8384
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 22002 8412 22008 8424
rect 19383 8384 22008 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 20901 8347 20959 8353
rect 20901 8313 20913 8347
rect 20947 8344 20959 8347
rect 21266 8344 21272 8356
rect 20947 8316 21272 8344
rect 20947 8313 20959 8316
rect 20901 8307 20959 8313
rect 21266 8304 21272 8316
rect 21324 8304 21330 8356
rect 22296 8344 22324 8443
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 22554 8372 22560 8424
rect 22612 8372 22618 8424
rect 24578 8372 24584 8424
rect 24636 8372 24642 8424
rect 24854 8344 24860 8356
rect 22296 8316 24860 8344
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 4080 8044 6653 8072
rect 4080 7945 4108 8044
rect 6641 8041 6653 8044
rect 6687 8072 6699 8075
rect 6822 8072 6828 8084
rect 6687 8044 6828 8072
rect 6687 8041 6699 8044
rect 6641 8035 6699 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 22370 8032 22376 8084
rect 22428 8072 22434 8084
rect 25225 8075 25283 8081
rect 25225 8072 25237 8075
rect 22428 8044 25237 8072
rect 22428 8032 22434 8044
rect 25225 8041 25237 8044
rect 25271 8041 25283 8075
rect 25225 8035 25283 8041
rect 4065 7939 4123 7945
rect 4065 7905 4077 7939
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7936 6147 7939
rect 6178 7936 6184 7948
rect 6135 7908 6184 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6638 7936 6644 7948
rect 6503 7908 6644 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6472 7868 6500 7899
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 5474 7840 6500 7868
rect 19794 7828 19800 7880
rect 19852 7868 19858 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19852 7840 20453 7868
rect 19852 7828 19858 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 20588 7840 21281 7868
rect 20588 7828 20594 7840
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7868 22891 7871
rect 23474 7868 23480 7880
rect 22879 7840 23480 7868
rect 22879 7837 22891 7840
rect 22833 7831 22891 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7868 24639 7871
rect 25038 7868 25044 7880
rect 24627 7840 25044 7868
rect 24627 7837 24639 7840
rect 24581 7831 24639 7837
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 20257 7735 20315 7741
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 20806 7732 20812 7744
rect 20303 7704 20812 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 17368 7432 18797 7460
rect 17368 7420 17374 7432
rect 18785 7429 18797 7432
rect 18831 7429 18843 7463
rect 18785 7423 18843 7429
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20898 7392 20904 7404
rect 20303 7364 20904 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 22060 7364 22109 7392
rect 22060 7352 22066 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 23290 7352 23296 7404
rect 23348 7392 23354 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23348 7364 23949 7392
rect 23348 7352 23354 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21634 7324 21640 7336
rect 21315 7296 21640 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22557 7327 22615 7333
rect 22557 7324 22569 7327
rect 22336 7296 22569 7324
rect 22336 7284 22342 7296
rect 22557 7293 22569 7296
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 24670 7284 24676 7336
rect 24728 7284 24734 7336
rect 18969 7259 19027 7265
rect 18969 7225 18981 7259
rect 19015 7256 19027 7259
rect 20622 7256 20628 7268
rect 19015 7228 20628 7256
rect 19015 7225 19027 7228
rect 18969 7219 19027 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 22370 6876 22376 6928
rect 22428 6916 22434 6928
rect 22738 6916 22744 6928
rect 22428 6888 22744 6916
rect 22428 6876 22434 6888
rect 22738 6876 22744 6888
rect 22796 6876 22802 6928
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 10686 6848 10692 6860
rect 5868 6820 10692 6848
rect 5868 6808 5874 6820
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 6362 6780 6368 6792
rect 4120 6752 6368 6780
rect 4120 6740 4126 6752
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 16448 6752 19717 6780
rect 16448 6740 16454 6752
rect 19705 6749 19717 6752
rect 19751 6780 19763 6783
rect 19981 6783 20039 6789
rect 19981 6780 19993 6783
rect 19751 6752 19993 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 19981 6749 19993 6752
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 22830 6740 22836 6792
rect 22888 6740 22894 6792
rect 24118 6740 24124 6792
rect 24176 6780 24182 6792
rect 24857 6783 24915 6789
rect 24857 6780 24869 6783
rect 24176 6752 24869 6780
rect 24176 6740 24182 6752
rect 24857 6749 24869 6752
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 22002 6672 22008 6724
rect 22060 6672 22066 6724
rect 23845 6715 23903 6721
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 24946 6712 24952 6724
rect 23891 6684 24952 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 24946 6672 24952 6684
rect 25004 6672 25010 6724
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 18564 6616 19533 6644
rect 18564 6604 18570 6616
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 24670 6604 24676 6656
rect 24728 6604 24734 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 4338 6440 4344 6452
rect 3743 6412 4344 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 11664 6412 17969 6440
rect 11664 6400 11670 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 17972 6304 18000 6403
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17972 6276 18245 6304
rect 3053 6267 3111 6273
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 21082 6304 21088 6316
rect 20303 6276 21088 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21416 6276 22017 6304
rect 21416 6264 21422 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 22244 6276 23949 6304
rect 22244 6264 22250 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6236 19303 6239
rect 20806 6236 20812 6248
rect 19291 6208 20812 6236
rect 19291 6205 19303 6208
rect 19245 6199 19303 6205
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21726 6236 21732 6248
rect 21315 6208 21732 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 21968 6208 22477 6236
rect 21968 6196 21974 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 24578 6196 24584 6248
rect 24636 6196 24642 6248
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 20956 5868 24777 5896
rect 20956 5856 20962 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20993 5763 21051 5769
rect 20993 5760 21005 5763
rect 20496 5732 21005 5760
rect 20496 5720 20502 5732
rect 20993 5729 21005 5732
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21542 5720 21548 5772
rect 21600 5760 21606 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 21600 5732 22845 5760
rect 21600 5720 21606 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 11974 5692 11980 5704
rect 7156 5664 11980 5692
rect 7156 5652 7162 5664
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 17678 5652 17684 5704
rect 17736 5652 17742 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 20404 5664 20545 5692
rect 20404 5652 20410 5664
rect 20533 5661 20545 5664
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 20680 5664 22385 5692
rect 20680 5652 20686 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 22462 5652 22468 5704
rect 22520 5692 22526 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 22520 5664 24685 5692
rect 22520 5652 22526 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 18693 5627 18751 5633
rect 18693 5593 18705 5627
rect 18739 5624 18751 5627
rect 21082 5624 21088 5636
rect 18739 5596 21088 5624
rect 18739 5593 18751 5596
rect 18693 5587 18751 5593
rect 21082 5584 21088 5596
rect 21140 5584 21146 5636
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 4706 5556 4712 5568
rect 3476 5528 4712 5556
rect 3476 5516 3482 5528
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2866 5352 2872 5364
rect 1627 5324 2872 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19702 5284 19708 5296
rect 18831 5256 19708 5284
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19702 5244 19708 5256
rect 19760 5244 19766 5296
rect 1762 5176 1768 5228
rect 1820 5176 1826 5228
rect 17770 5176 17776 5228
rect 17828 5176 17834 5228
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 21818 5176 21824 5228
rect 21876 5216 21882 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21876 5188 22017 5216
rect 21876 5176 21882 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 24026 5176 24032 5228
rect 24084 5176 24090 5228
rect 19610 5108 19616 5160
rect 19668 5148 19674 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19668 5120 19901 5148
rect 19668 5108 19674 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 22462 5108 22468 5160
rect 22520 5108 22526 5160
rect 24762 5108 24768 5160
rect 24820 5108 24826 5160
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 23845 4811 23903 4817
rect 23845 4808 23857 4811
rect 17828 4780 23857 4808
rect 17828 4768 17834 4780
rect 23845 4777 23857 4780
rect 23891 4777 23903 4811
rect 23845 4771 23903 4777
rect 2041 4743 2099 4749
rect 2041 4709 2053 4743
rect 2087 4740 2099 4743
rect 4890 4740 4896 4752
rect 2087 4712 4896 4740
rect 2087 4709 2099 4712
rect 2041 4703 2099 4709
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 24854 4700 24860 4752
rect 24912 4700 24918 4752
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 12618 4672 12624 4684
rect 11848 4644 12624 4672
rect 11848 4632 11854 4644
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 19886 4632 19892 4684
rect 19944 4632 19950 4684
rect 20714 4632 20720 4684
rect 20772 4672 20778 4684
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 20772 4644 21741 4672
rect 20772 4632 20778 4644
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18506 4604 18512 4616
rect 17727 4576 18512 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 18656 4576 19441 4604
rect 18656 4564 18662 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 22738 4564 22744 4616
rect 22796 4604 22802 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 22796 4576 24041 4604
rect 22796 4564 22802 4576
rect 24029 4573 24041 4576
rect 24075 4573 24087 4607
rect 24029 4567 24087 4573
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4536 1915 4539
rect 2038 4536 2044 4548
rect 1903 4508 2044 4536
rect 1903 4505 1915 4508
rect 1857 4499 1915 4505
rect 2038 4496 2044 4508
rect 2096 4536 2102 4548
rect 2317 4539 2375 4545
rect 2317 4536 2329 4539
rect 2096 4508 2329 4536
rect 2096 4496 2102 4508
rect 2317 4505 2329 4508
rect 2363 4505 2375 4539
rect 2317 4499 2375 4505
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 20622 4536 20628 4548
rect 18739 4508 20628 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 23290 4496 23296 4548
rect 23348 4536 23354 4548
rect 24673 4539 24731 4545
rect 24673 4536 24685 4539
rect 23348 4508 24685 4536
rect 23348 4496 23354 4508
rect 24673 4505 24685 4508
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 14182 4468 14188 4480
rect 12676 4440 14188 4468
rect 12676 4428 12682 4440
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 2409 4267 2467 4273
rect 2409 4264 2421 4267
rect 1820 4236 2421 4264
rect 1820 4224 1826 4236
rect 2409 4233 2421 4236
rect 2455 4233 2467 4267
rect 2409 4227 2467 4233
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 10318 4264 10324 4276
rect 9364 4236 10324 4264
rect 9364 4224 9370 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13596 4236 13676 4264
rect 13596 4224 13602 4236
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2222 4128 2228 4140
rect 1811 4100 2228 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 13648 4137 13676 4236
rect 25130 4156 25136 4208
rect 25188 4156 25194 4208
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2464 4100 2881 4128
rect 2464 4088 2470 4100
rect 2869 4097 2881 4100
rect 2915 4128 2927 4131
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 2915 4100 3433 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 5994 4060 6000 4072
rect 4120 4032 6000 4060
rect 4120 4020 4126 4032
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 11606 4060 11612 4072
rect 11379 4032 11612 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11606 4020 11612 4032
rect 11664 4060 11670 4072
rect 11701 4063 11759 4069
rect 11701 4060 11713 4063
rect 11664 4032 11713 4060
rect 11664 4020 11670 4032
rect 11701 4029 11713 4032
rect 11747 4029 11759 4063
rect 11701 4023 11759 4029
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 3053 3995 3111 4001
rect 3053 3961 3065 3995
rect 3099 3992 3111 3995
rect 3418 3992 3424 4004
rect 3099 3964 3424 3992
rect 3099 3961 3111 3964
rect 3053 3955 3111 3961
rect 3418 3952 3424 3964
rect 3476 3952 3482 4004
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9953 3995 10011 4001
rect 9953 3992 9965 3995
rect 9088 3964 9965 3992
rect 9088 3952 9094 3964
rect 9953 3961 9965 3964
rect 9999 3961 10011 3995
rect 9953 3955 10011 3961
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 9490 3884 9496 3936
rect 9548 3884 9554 3936
rect 9766 3884 9772 3936
rect 9824 3884 9830 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10376 3896 11069 3924
rect 10376 3884 10382 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11992 3924 12020 4023
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13504 4032 14013 4060
rect 13504 4020 13510 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 12158 3952 12164 4004
rect 12216 3992 12222 4004
rect 16132 3992 16160 4091
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16724 4100 16865 4128
rect 16724 4088 16730 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 24121 4131 24179 4137
rect 24121 4097 24133 4131
rect 24167 4128 24179 4131
rect 24670 4128 24676 4140
rect 24167 4100 24676 4128
rect 24167 4097 24179 4100
rect 24121 4091 24179 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16448 4032 17325 4060
rect 16448 4020 16454 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 17552 4032 19165 4060
rect 17552 4020 17558 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 20070 4020 20076 4072
rect 20128 4060 20134 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 20128 4032 22477 4060
rect 20128 4020 20134 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 12216 3964 16160 3992
rect 12216 3952 12222 3964
rect 19702 3952 19708 4004
rect 19760 3992 19766 4004
rect 22094 3992 22100 4004
rect 19760 3964 22100 3992
rect 19760 3952 19766 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 15930 3924 15936 3936
rect 11992 3896 15936 3924
rect 11057 3887 11115 3893
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16209 3927 16267 3933
rect 16209 3893 16221 3927
rect 16255 3924 16267 3927
rect 22186 3924 22192 3936
rect 16255 3896 22192 3924
rect 16255 3893 16267 3896
rect 16209 3887 16267 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 1946 3680 1952 3732
rect 2004 3680 2010 3732
rect 2682 3680 2688 3732
rect 2740 3680 2746 3732
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 4246 3720 4252 3732
rect 3283 3692 4252 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 8202 3680 8208 3732
rect 8260 3680 8266 3732
rect 9306 3680 9312 3732
rect 9364 3680 9370 3732
rect 10042 3680 10048 3732
rect 10100 3680 10106 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 18782 3720 18788 3732
rect 18647 3692 18788 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 5261 3655 5319 3661
rect 5261 3621 5273 3655
rect 5307 3621 5319 3655
rect 5261 3615 5319 3621
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 12158 3652 12164 3664
rect 5951 3624 12164 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 3510 3584 3516 3596
rect 1780 3556 3516 3584
rect 1780 3525 1808 3556
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 5276 3584 5304 3615
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 15102 3652 15108 3664
rect 12406 3624 15108 3652
rect 8938 3584 8944 3596
rect 5276 3556 8944 3584
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 12406 3584 12434 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 20806 3612 20812 3664
rect 20864 3652 20870 3664
rect 24946 3652 24952 3664
rect 20864 3624 24952 3652
rect 20864 3612 20870 3624
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 11287 3556 12434 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12768 3556 12817 3584
rect 12768 3544 12774 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 14918 3544 14924 3596
rect 14976 3584 14982 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 14976 3556 15485 3584
rect 14976 3544 14982 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 16080 3556 17325 3584
rect 16080 3544 16086 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 19889 3587 19947 3593
rect 19889 3584 19901 3587
rect 17920 3556 19901 3584
rect 17920 3544 17926 3556
rect 19889 3553 19901 3556
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 1535 3488 1777 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 2866 3516 2872 3528
rect 2547 3488 2872 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3467 3488 3801 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 3789 3479 3847 3485
rect 5000 3488 5089 3516
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 3436 3448 3464 3479
rect 1728 3420 3464 3448
rect 1728 3408 1734 3420
rect 5000 3392 5028 3488
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 7834 3516 7840 3528
rect 7791 3488 7840 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 7834 3476 7840 3488
rect 7892 3516 7898 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7892 3488 8033 3516
rect 7892 3476 7898 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3516 9183 3519
rect 9490 3516 9496 3528
rect 9171 3488 9496 3516
rect 9171 3485 9183 3488
rect 9125 3479 9183 3485
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9824 3488 9873 3516
rect 9824 3476 9830 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10870 3516 10876 3528
rect 10551 3488 10876 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10928 3488 10977 3516
rect 10928 3476 10934 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15562 3516 15568 3528
rect 15151 3488 15568 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16298 3476 16304 3528
rect 16356 3516 16362 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16356 3488 16865 3516
rect 16356 3476 16362 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19392 3488 19441 3516
rect 19392 3476 19398 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 21174 3476 21180 3528
rect 21232 3516 21238 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21232 3488 21281 3516
rect 21232 3476 21238 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 7561 3451 7619 3457
rect 7561 3417 7573 3451
rect 7607 3448 7619 3451
rect 8294 3448 8300 3460
rect 7607 3420 8300 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 21744 3448 21772 3547
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3516 24087 3519
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24075 3488 24593 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 19024 3420 21772 3448
rect 23400 3448 23428 3479
rect 24118 3448 24124 3460
rect 23400 3420 24124 3448
rect 19024 3408 19030 3420
rect 24118 3408 24124 3420
rect 24176 3408 24182 3460
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4982 3380 4988 3392
rect 4847 3352 4988 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 6880 3352 7205 3380
rect 6880 3340 6886 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 11238 3380 11244 3392
rect 10735 3352 11244 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 11238 3340 11244 3352
rect 11296 3380 11302 3392
rect 11698 3380 11704 3392
rect 11296 3352 11704 3380
rect 11296 3340 11302 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22830 3380 22836 3392
rect 22060 3352 22836 3380
rect 22060 3340 22066 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 25225 3383 25283 3389
rect 25225 3380 25237 3383
rect 24636 3352 25237 3380
rect 24636 3340 24642 3352
rect 25225 3349 25237 3352
rect 25271 3349 25283 3383
rect 25225 3343 25283 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 2866 3136 2872 3188
rect 2924 3136 2930 3188
rect 5166 3136 5172 3188
rect 5224 3136 5230 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3176 6515 3179
rect 6546 3176 6552 3188
rect 6503 3148 6552 3176
rect 6503 3145 6515 3148
rect 6457 3139 6515 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 7006 3136 7012 3188
rect 7064 3136 7070 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7248 3148 7757 3176
rect 7248 3136 7254 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 8846 3176 8852 3188
rect 8527 3148 8852 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11388 3148 11897 3176
rect 11388 3136 11394 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 25038 3136 25044 3188
rect 25096 3176 25102 3188
rect 25133 3179 25191 3185
rect 25133 3176 25145 3179
rect 25096 3148 25145 3176
rect 25096 3136 25102 3148
rect 25133 3145 25145 3148
rect 25179 3145 25191 3179
rect 25133 3139 25191 3145
rect 13630 3108 13636 3120
rect 10612 3080 13636 3108
rect 1578 3000 1584 3052
rect 1636 3000 1642 3052
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4755 3012 4997 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5350 3040 5356 3052
rect 5031 3012 5356 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8202 3040 8208 3052
rect 7607 3012 8208 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8662 3040 8668 3052
rect 8343 3012 8668 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9030 3000 9036 3052
rect 9088 3000 9094 3052
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9582 3040 9588 3052
rect 9355 3012 9588 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 10612 3049 10640 3080
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 12618 3000 12624 3052
rect 12676 3000 12682 3052
rect 14274 3000 14280 3052
rect 14332 3000 14338 3052
rect 16850 3000 16856 3052
rect 16908 3000 16914 3052
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 2777 2975 2835 2981
rect 2777 2941 2789 2975
rect 2823 2972 2835 2975
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 2823 2944 3249 2972
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 3237 2941 3249 2944
rect 3283 2972 3295 2975
rect 3418 2972 3424 2984
rect 3283 2944 3424 2972
rect 3283 2941 3295 2944
rect 3237 2935 3295 2941
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 10410 2972 10416 2984
rect 3559 2944 10416 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 13354 2932 13360 2984
rect 13412 2932 13418 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14240 2944 14749 2972
rect 14240 2932 14246 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15712 2944 17325 2972
rect 15712 2932 15718 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 17126 2864 17132 2916
rect 17184 2904 17190 2916
rect 19168 2904 19196 2935
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 23382 2972 23388 2984
rect 20680 2944 23388 2972
rect 20680 2932 20686 2944
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 17184 2876 19196 2904
rect 17184 2864 17190 2876
rect 19702 2864 19708 2916
rect 19760 2904 19766 2916
rect 20714 2904 20720 2916
rect 19760 2876 20720 2904
rect 19760 2864 19766 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 20806 2864 20812 2916
rect 20864 2904 20870 2916
rect 22462 2904 22468 2916
rect 20864 2876 22468 2904
rect 20864 2864 20870 2876
rect 22462 2864 22468 2876
rect 22520 2864 22526 2916
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4341 2839 4399 2845
rect 4341 2836 4353 2839
rect 4304 2808 4353 2836
rect 4304 2796 4310 2808
rect 4341 2805 4353 2808
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17954 2836 17960 2848
rect 16816 2808 17960 2836
rect 16816 2796 16822 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 19886 2836 19892 2848
rect 18656 2808 19892 2836
rect 18656 2796 18662 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 21726 2796 21732 2848
rect 21784 2836 21790 2848
rect 22646 2836 22652 2848
rect 21784 2808 22652 2836
rect 21784 2796 21790 2808
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 24118 2796 24124 2848
rect 24176 2796 24182 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 1636 2604 2237 2632
rect 1636 2592 1642 2604
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 3326 2592 3332 2644
rect 3384 2592 3390 2644
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 7098 2592 7104 2644
rect 7156 2592 7162 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9858 2632 9864 2644
rect 9815 2604 9864 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 15378 2632 15384 2644
rect 11747 2604 15384 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 18601 2635 18659 2641
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 18690 2632 18696 2644
rect 18647 2604 18696 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 25225 2635 25283 2641
rect 25225 2601 25237 2635
rect 25271 2632 25283 2635
rect 25314 2632 25320 2644
rect 25271 2604 25320 2632
rect 25271 2601 25283 2604
rect 25225 2595 25283 2601
rect 25314 2592 25320 2604
rect 25372 2592 25378 2644
rect 11790 2564 11796 2576
rect 7944 2536 11796 2564
rect 7944 2505 7972 2536
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 17586 2524 17592 2576
rect 17644 2564 17650 2576
rect 17644 2536 22048 2564
rect 17644 2524 17650 2536
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 4724 2468 5825 2496
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2428 1639 2431
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 1627 2400 2513 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3145 2431 3203 2437
rect 3145 2428 3157 2431
rect 2915 2400 3157 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3145 2397 3157 2400
rect 3191 2428 3203 2431
rect 3878 2428 3884 2440
rect 3191 2400 3884 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4246 2428 4252 2440
rect 4019 2400 4252 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4724 2437 4752 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 11698 2496 11704 2508
rect 10643 2468 11704 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11974 2496 11980 2508
rect 11900 2468 11980 2496
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5994 2428 6000 2440
rect 5031 2400 6000 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6503 2400 6929 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 7190 2428 7196 2440
rect 6963 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9171 2400 9597 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9585 2397 9597 2400
rect 9631 2428 9643 2431
rect 10134 2428 10140 2440
rect 9631 2400 10140 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11900 2437 11928 2468
rect 11974 2456 11980 2468
rect 12032 2496 12038 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 12032 2468 14105 2496
rect 12032 2456 12038 2468
rect 14093 2465 14105 2468
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14608 2468 15209 2496
rect 14608 2456 14614 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 15344 2468 17325 2496
rect 15344 2456 15350 2468
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 18012 2468 19901 2496
rect 18012 2456 18018 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12802 2428 12808 2440
rect 12575 2400 12808 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5776 2332 6101 2360
rect 5776 2320 5782 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7576 2360 7604 2388
rect 6687 2332 7604 2360
rect 9309 2363 9367 2369
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 10336 2360 10364 2391
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 14642 2388 14648 2440
rect 14700 2388 14706 2440
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 22020 2437 22048 2536
rect 22465 2499 22523 2505
rect 22465 2465 22477 2499
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 24029 2499 24087 2505
rect 24029 2465 24041 2499
rect 24075 2496 24087 2499
rect 24854 2496 24860 2508
rect 24075 2468 24860 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 12342 2360 12348 2372
rect 9355 2332 12348 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2360 13599 2363
rect 13814 2360 13820 2372
rect 13587 2332 13820 2360
rect 13587 2329 13599 2332
rect 13541 2323 13599 2329
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 22480 2360 22508 2459
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 18380 2332 22508 2360
rect 18380 2320 18386 2332
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 3976 54315 4028 54324
rect 3976 54281 3985 54315
rect 3985 54281 4019 54315
rect 4019 54281 4028 54315
rect 3976 54272 4028 54281
rect 9956 54272 10008 54324
rect 14740 54272 14792 54324
rect 16212 54272 16264 54324
rect 7840 54204 7892 54256
rect 11428 54204 11480 54256
rect 2320 54136 2372 54188
rect 5356 54136 5408 54188
rect 5908 54068 5960 54120
rect 9956 54179 10008 54188
rect 9956 54145 9965 54179
rect 9965 54145 9999 54179
rect 9999 54145 10008 54179
rect 9956 54136 10008 54145
rect 12900 54204 12952 54256
rect 12348 54179 12400 54188
rect 12348 54145 12357 54179
rect 12357 54145 12391 54179
rect 12391 54145 12400 54179
rect 12348 54136 12400 54145
rect 15200 54136 15252 54188
rect 24492 54315 24544 54324
rect 24492 54281 24501 54315
rect 24501 54281 24535 54315
rect 24535 54281 24544 54315
rect 24492 54272 24544 54281
rect 17684 54204 17736 54256
rect 18880 54204 18932 54256
rect 16948 54136 17000 54188
rect 11244 54068 11296 54120
rect 12532 54068 12584 54120
rect 18420 54068 18472 54120
rect 19524 54136 19576 54188
rect 20720 54136 20772 54188
rect 21364 54136 21416 54188
rect 22468 54136 22520 54188
rect 24952 54179 25004 54188
rect 24952 54145 24961 54179
rect 24961 54145 24995 54179
rect 24995 54145 25004 54179
rect 24952 54136 25004 54145
rect 19708 54068 19760 54120
rect 15568 54000 15620 54052
rect 3792 53975 3844 53984
rect 3792 53941 3801 53975
rect 3801 53941 3835 53975
rect 3835 53941 3844 53975
rect 3792 53932 3844 53941
rect 12256 53932 12308 53984
rect 14924 53932 14976 53984
rect 15200 53932 15252 53984
rect 17040 53975 17092 53984
rect 17040 53941 17049 53975
rect 17049 53941 17083 53975
rect 17083 53941 17092 53975
rect 17040 53932 17092 53941
rect 18420 53932 18472 53984
rect 19340 53932 19392 53984
rect 20904 53932 20956 53984
rect 21640 53932 21692 53984
rect 22192 53975 22244 53984
rect 22192 53941 22201 53975
rect 22201 53941 22235 53975
rect 22235 53941 22244 53975
rect 22192 53932 22244 53941
rect 22284 53932 22336 53984
rect 23940 53975 23992 53984
rect 23940 53941 23949 53975
rect 23949 53941 23983 53975
rect 23983 53941 23992 53975
rect 23940 53932 23992 53941
rect 25780 53932 25832 53984
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 16580 53728 16632 53780
rect 18880 53771 18932 53780
rect 18880 53737 18889 53771
rect 18889 53737 18923 53771
rect 18923 53737 18932 53771
rect 18880 53728 18932 53737
rect 5540 53660 5592 53712
rect 21548 53660 21600 53712
rect 22376 53660 22428 53712
rect 7380 53592 7432 53644
rect 8852 53592 8904 53644
rect 11060 53635 11112 53644
rect 11060 53601 11069 53635
rect 11069 53601 11103 53635
rect 11103 53601 11112 53635
rect 11060 53592 11112 53601
rect 12164 53592 12216 53644
rect 3976 53567 4028 53576
rect 3976 53533 3985 53567
rect 3985 53533 4019 53567
rect 4019 53533 4028 53567
rect 3976 53524 4028 53533
rect 5540 53567 5592 53576
rect 5540 53533 5549 53567
rect 5549 53533 5583 53567
rect 5583 53533 5592 53567
rect 5540 53524 5592 53533
rect 9128 53524 9180 53576
rect 12072 53524 12124 53576
rect 12624 53524 12676 53576
rect 14004 53524 14056 53576
rect 15476 53524 15528 53576
rect 16580 53524 16632 53576
rect 17316 53524 17368 53576
rect 18328 53524 18380 53576
rect 19156 53524 19208 53576
rect 19892 53524 19944 53576
rect 20996 53524 21048 53576
rect 21732 53524 21784 53576
rect 22100 53524 22152 53576
rect 22836 53524 22888 53576
rect 23388 53524 23440 53576
rect 24768 53524 24820 53576
rect 7564 53456 7616 53508
rect 16396 53456 16448 53508
rect 18512 53456 18564 53508
rect 20628 53456 20680 53508
rect 24032 53499 24084 53508
rect 24032 53465 24041 53499
rect 24041 53465 24075 53499
rect 24075 53465 24084 53499
rect 24032 53456 24084 53465
rect 4620 53431 4672 53440
rect 4620 53397 4629 53431
rect 4629 53397 4663 53431
rect 4663 53397 4672 53431
rect 4620 53388 4672 53397
rect 14464 53431 14516 53440
rect 14464 53397 14473 53431
rect 14473 53397 14507 53431
rect 14507 53397 14516 53431
rect 14464 53388 14516 53397
rect 16856 53431 16908 53440
rect 16856 53397 16865 53431
rect 16865 53397 16899 53431
rect 16899 53397 16908 53431
rect 16856 53388 16908 53397
rect 17408 53431 17460 53440
rect 17408 53397 17417 53431
rect 17417 53397 17451 53431
rect 17451 53397 17460 53431
rect 17408 53388 17460 53397
rect 19616 53431 19668 53440
rect 19616 53397 19625 53431
rect 19625 53397 19659 53431
rect 19659 53397 19668 53431
rect 19616 53388 19668 53397
rect 21364 53388 21416 53440
rect 22468 53431 22520 53440
rect 22468 53397 22477 53431
rect 22477 53397 22511 53431
rect 22511 53397 22520 53431
rect 22468 53388 22520 53397
rect 25688 53388 25740 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 5172 53184 5224 53236
rect 6184 53184 6236 53236
rect 17316 53227 17368 53236
rect 17316 53193 17325 53227
rect 17325 53193 17359 53227
rect 17359 53193 17368 53227
rect 17316 53184 17368 53193
rect 19156 53184 19208 53236
rect 19708 53227 19760 53236
rect 19708 53193 19717 53227
rect 19717 53193 19751 53227
rect 19751 53193 19760 53227
rect 19708 53184 19760 53193
rect 20996 53227 21048 53236
rect 20996 53193 21005 53227
rect 21005 53193 21039 53227
rect 21039 53193 21048 53227
rect 20996 53184 21048 53193
rect 21732 53184 21784 53236
rect 22100 53184 22152 53236
rect 22560 53227 22612 53236
rect 22560 53193 22569 53227
rect 22569 53193 22603 53227
rect 22603 53193 22612 53227
rect 22560 53184 22612 53193
rect 23296 53184 23348 53236
rect 4436 53116 4488 53168
rect 6276 53116 6328 53168
rect 9220 53116 9272 53168
rect 13636 53116 13688 53168
rect 20720 53116 20772 53168
rect 1676 53091 1728 53100
rect 1676 53057 1685 53091
rect 1685 53057 1719 53091
rect 1719 53057 1728 53091
rect 1676 53048 1728 53057
rect 4160 53048 4212 53100
rect 4712 53091 4764 53100
rect 4712 53057 4721 53091
rect 4721 53057 4755 53091
rect 4755 53057 4764 53091
rect 4712 53048 4764 53057
rect 7288 53048 7340 53100
rect 9312 53048 9364 53100
rect 11888 53091 11940 53100
rect 11888 53057 11897 53091
rect 11897 53057 11931 53091
rect 11931 53057 11940 53091
rect 11888 53048 11940 53057
rect 14372 53048 14424 53100
rect 15844 53048 15896 53100
rect 18788 53048 18840 53100
rect 20260 53048 20312 53100
rect 23572 53048 23624 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 10324 53023 10376 53032
rect 10324 52989 10333 53023
rect 10333 52989 10367 53023
rect 10367 52989 10376 53023
rect 10324 52980 10376 52989
rect 11796 52980 11848 53032
rect 1860 52912 1912 52964
rect 3516 52912 3568 52964
rect 14004 52955 14056 52964
rect 14004 52921 14013 52955
rect 14013 52921 14047 52955
rect 14047 52921 14056 52955
rect 14004 52912 14056 52921
rect 1768 52844 1820 52896
rect 14740 52844 14792 52896
rect 15936 52887 15988 52896
rect 15936 52853 15945 52887
rect 15945 52853 15979 52887
rect 15979 52853 15988 52887
rect 15936 52844 15988 52853
rect 18604 52844 18656 52896
rect 20168 52844 20220 52896
rect 22192 52844 22244 52896
rect 23388 52844 23440 52896
rect 24952 52844 25004 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 2228 52640 2280 52692
rect 3424 52640 3476 52692
rect 12624 52683 12676 52692
rect 12624 52649 12633 52683
rect 12633 52649 12667 52683
rect 12667 52649 12676 52683
rect 12624 52640 12676 52649
rect 13636 52640 13688 52692
rect 24768 52640 24820 52692
rect 1308 52572 1360 52624
rect 3792 52572 3844 52624
rect 3700 52504 3752 52556
rect 25964 52572 26016 52624
rect 5172 52436 5224 52488
rect 6000 52436 6052 52488
rect 6644 52436 6696 52488
rect 7380 52479 7432 52488
rect 7380 52445 7389 52479
rect 7389 52445 7423 52479
rect 7423 52445 7432 52479
rect 7380 52436 7432 52445
rect 7748 52547 7800 52556
rect 7748 52513 7757 52547
rect 7757 52513 7791 52547
rect 7791 52513 7800 52547
rect 7748 52504 7800 52513
rect 10692 52504 10744 52556
rect 8668 52436 8720 52488
rect 9588 52436 9640 52488
rect 12808 52479 12860 52488
rect 12808 52445 12817 52479
rect 12817 52445 12851 52479
rect 12851 52445 12860 52479
rect 12808 52436 12860 52445
rect 13544 52436 13596 52488
rect 24768 52479 24820 52488
rect 24768 52445 24777 52479
rect 24777 52445 24811 52479
rect 24811 52445 24820 52479
rect 24768 52436 24820 52445
rect 13360 52368 13412 52420
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 1676 52096 1728 52148
rect 4160 52096 4212 52148
rect 11888 52096 11940 52148
rect 12348 52139 12400 52148
rect 12348 52105 12357 52139
rect 12357 52105 12391 52139
rect 12391 52105 12400 52139
rect 12348 52096 12400 52105
rect 13360 52096 13412 52148
rect 25320 52139 25372 52148
rect 25320 52105 25329 52139
rect 25329 52105 25363 52139
rect 25363 52105 25372 52139
rect 25320 52096 25372 52105
rect 4620 52028 4672 52080
rect 9036 52028 9088 52080
rect 7196 51960 7248 52012
rect 3332 51935 3384 51944
rect 3332 51901 3341 51935
rect 3341 51901 3375 51935
rect 3375 51901 3384 51935
rect 3332 51892 3384 51901
rect 4896 51892 4948 51944
rect 9680 52003 9732 52012
rect 9680 51969 9689 52003
rect 9689 51969 9723 52003
rect 9723 51969 9732 52003
rect 9680 51960 9732 51969
rect 10876 51960 10928 52012
rect 11980 51960 12032 52012
rect 8484 51935 8536 51944
rect 8484 51901 8493 51935
rect 8493 51901 8527 51935
rect 8527 51901 8536 51935
rect 8484 51892 8536 51901
rect 9772 51892 9824 51944
rect 10416 51824 10468 51876
rect 4896 51756 4948 51808
rect 25504 51799 25556 51808
rect 25504 51765 25513 51799
rect 25513 51765 25547 51799
rect 25547 51765 25556 51799
rect 25504 51756 25556 51765
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 9956 51552 10008 51604
rect 2872 51459 2924 51468
rect 2872 51425 2881 51459
rect 2881 51425 2915 51459
rect 2915 51425 2924 51459
rect 2872 51416 2924 51425
rect 6920 51416 6972 51468
rect 7012 51416 7064 51468
rect 3976 51391 4028 51400
rect 3976 51357 3985 51391
rect 3985 51357 4019 51391
rect 4019 51357 4028 51391
rect 3976 51348 4028 51357
rect 6736 51348 6788 51400
rect 7104 51391 7156 51400
rect 7104 51357 7113 51391
rect 7113 51357 7147 51391
rect 7147 51357 7156 51391
rect 7104 51348 7156 51357
rect 9220 51348 9272 51400
rect 25504 51348 25556 51400
rect 6184 51323 6236 51332
rect 6184 51289 6193 51323
rect 6193 51289 6227 51323
rect 6227 51289 6236 51323
rect 6184 51280 6236 51289
rect 7012 51280 7064 51332
rect 7196 51280 7248 51332
rect 4252 51212 4304 51264
rect 25228 51255 25280 51264
rect 25228 51221 25237 51255
rect 25237 51221 25271 51255
rect 25271 51221 25280 51255
rect 25228 51212 25280 51221
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 3976 51008 4028 51060
rect 6920 51051 6972 51060
rect 6920 51017 6929 51051
rect 6929 51017 6963 51051
rect 6963 51017 6972 51051
rect 6920 51008 6972 51017
rect 2320 50940 2372 50992
rect 1768 50915 1820 50924
rect 1768 50881 1777 50915
rect 1777 50881 1811 50915
rect 1811 50881 1820 50915
rect 1768 50872 1820 50881
rect 2780 50847 2832 50856
rect 2780 50813 2789 50847
rect 2789 50813 2823 50847
rect 2823 50813 2832 50847
rect 2780 50804 2832 50813
rect 5448 50872 5500 50924
rect 7656 50872 7708 50924
rect 9588 50983 9640 50992
rect 9588 50949 9597 50983
rect 9597 50949 9631 50983
rect 9631 50949 9640 50983
rect 9588 50940 9640 50949
rect 7840 50872 7892 50924
rect 25044 50915 25096 50924
rect 25044 50881 25053 50915
rect 25053 50881 25087 50915
rect 25087 50881 25096 50915
rect 25044 50872 25096 50881
rect 4344 50804 4396 50856
rect 7472 50847 7524 50856
rect 7472 50813 7481 50847
rect 7481 50813 7515 50847
rect 7515 50813 7524 50847
rect 7472 50804 7524 50813
rect 4160 50736 4212 50788
rect 25872 50668 25924 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 9128 50464 9180 50516
rect 1308 50328 1360 50380
rect 3424 50328 3476 50380
rect 5816 50260 5868 50312
rect 9404 50303 9456 50312
rect 9404 50269 9413 50303
rect 9413 50269 9447 50303
rect 9447 50269 9456 50303
rect 9404 50260 9456 50269
rect 8576 50192 8628 50244
rect 5080 50124 5132 50176
rect 25320 50124 25372 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 3516 49852 3568 49904
rect 1952 49827 2004 49836
rect 1952 49793 1961 49827
rect 1961 49793 1995 49827
rect 1995 49793 2004 49827
rect 1952 49784 2004 49793
rect 9864 49920 9916 49972
rect 20812 49920 20864 49972
rect 4252 49895 4304 49904
rect 4252 49861 4261 49895
rect 4261 49861 4295 49895
rect 4295 49861 4304 49895
rect 4252 49852 4304 49861
rect 8944 49852 8996 49904
rect 9312 49895 9364 49904
rect 9312 49861 9321 49895
rect 9321 49861 9355 49895
rect 9355 49861 9364 49895
rect 9312 49852 9364 49861
rect 7748 49784 7800 49836
rect 25320 49827 25372 49836
rect 25320 49793 25329 49827
rect 25329 49793 25363 49827
rect 25363 49793 25372 49827
rect 25320 49784 25372 49793
rect 8852 49716 8904 49768
rect 16028 49716 16080 49768
rect 16856 49716 16908 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 11980 49376 12032 49428
rect 1492 49240 1544 49292
rect 10692 49172 10744 49224
rect 25320 49215 25372 49224
rect 25320 49181 25329 49215
rect 25329 49181 25363 49215
rect 25363 49181 25372 49215
rect 25320 49172 25372 49181
rect 10784 49036 10836 49088
rect 19064 49036 19116 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 12808 48832 12860 48884
rect 12808 48696 12860 48748
rect 25504 48535 25556 48544
rect 25504 48501 25513 48535
rect 25513 48501 25547 48535
rect 25547 48501 25556 48535
rect 25504 48492 25556 48501
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 7288 48084 7340 48136
rect 9956 48084 10008 48136
rect 25320 48127 25372 48136
rect 25320 48093 25329 48127
rect 25329 48093 25363 48127
rect 25363 48093 25372 48127
rect 25320 48084 25372 48093
rect 1308 48016 1360 48068
rect 4068 47948 4120 48000
rect 17592 47948 17644 48000
rect 18420 47948 18472 48000
rect 20536 47948 20588 48000
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9036 47744 9088 47796
rect 15936 47744 15988 47796
rect 17408 47744 17460 47796
rect 11796 47608 11848 47660
rect 17592 47608 17644 47660
rect 18512 47651 18564 47660
rect 18512 47617 18521 47651
rect 18521 47617 18555 47651
rect 18555 47617 18564 47651
rect 18512 47608 18564 47617
rect 18696 47608 18748 47660
rect 25504 47608 25556 47660
rect 16304 47472 16356 47524
rect 18420 47472 18472 47524
rect 22744 47540 22796 47592
rect 16580 47404 16632 47456
rect 17500 47404 17552 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9864 47243 9916 47252
rect 9864 47209 9873 47243
rect 9873 47209 9907 47243
rect 9907 47209 9916 47243
rect 9864 47200 9916 47209
rect 18420 47200 18472 47252
rect 21456 47200 21508 47252
rect 18512 47132 18564 47184
rect 16672 47064 16724 47116
rect 17684 47064 17736 47116
rect 18604 47107 18656 47116
rect 18604 47073 18613 47107
rect 18613 47073 18647 47107
rect 18647 47073 18656 47107
rect 18604 47064 18656 47073
rect 19340 47064 19392 47116
rect 25596 47132 25648 47184
rect 22468 47107 22520 47116
rect 22468 47073 22477 47107
rect 22477 47073 22511 47107
rect 22511 47073 22520 47107
rect 22468 47064 22520 47073
rect 22836 47064 22888 47116
rect 8944 46928 8996 46980
rect 10508 46971 10560 46980
rect 10508 46937 10517 46971
rect 10517 46937 10551 46971
rect 10551 46937 10560 46971
rect 10508 46928 10560 46937
rect 10600 46860 10652 46912
rect 12624 46928 12676 46980
rect 16396 46928 16448 46980
rect 18328 46928 18380 46980
rect 19248 46971 19300 46980
rect 19248 46937 19257 46971
rect 19257 46937 19291 46971
rect 19291 46937 19300 46971
rect 19248 46928 19300 46937
rect 21456 46928 21508 46980
rect 24768 46928 24820 46980
rect 12164 46860 12216 46912
rect 17408 46860 17460 46912
rect 22008 46903 22060 46912
rect 22008 46869 22017 46903
rect 22017 46869 22051 46903
rect 22051 46869 22060 46903
rect 22008 46860 22060 46869
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 7472 46656 7524 46708
rect 10876 46699 10928 46708
rect 10876 46665 10885 46699
rect 10885 46665 10919 46699
rect 10919 46665 10928 46699
rect 10876 46656 10928 46665
rect 14464 46656 14516 46708
rect 18420 46656 18472 46708
rect 18972 46656 19024 46708
rect 21916 46656 21968 46708
rect 22100 46656 22152 46708
rect 23388 46656 23440 46708
rect 12716 46588 12768 46640
rect 15108 46588 15160 46640
rect 16396 46588 16448 46640
rect 17408 46588 17460 46640
rect 19248 46588 19300 46640
rect 9588 46520 9640 46572
rect 11060 46563 11112 46572
rect 11060 46529 11069 46563
rect 11069 46529 11103 46563
rect 11103 46529 11112 46563
rect 11060 46520 11112 46529
rect 11888 46316 11940 46368
rect 12716 46316 12768 46368
rect 16764 46452 16816 46504
rect 18604 46452 18656 46504
rect 13728 46316 13780 46368
rect 16304 46359 16356 46368
rect 16304 46325 16313 46359
rect 16313 46325 16347 46359
rect 16347 46325 16356 46359
rect 16304 46316 16356 46325
rect 16672 46316 16724 46368
rect 19340 46495 19392 46504
rect 19340 46461 19349 46495
rect 19349 46461 19383 46495
rect 19383 46461 19392 46495
rect 19340 46452 19392 46461
rect 22468 46452 22520 46504
rect 24492 46495 24544 46504
rect 24492 46461 24501 46495
rect 24501 46461 24535 46495
rect 24535 46461 24544 46495
rect 24492 46452 24544 46461
rect 24584 46452 24636 46504
rect 19524 46316 19576 46368
rect 21088 46359 21140 46368
rect 21088 46325 21097 46359
rect 21097 46325 21131 46359
rect 21131 46325 21140 46359
rect 21088 46316 21140 46325
rect 21916 46359 21968 46368
rect 21916 46325 21925 46359
rect 21925 46325 21959 46359
rect 21959 46325 21968 46359
rect 21916 46316 21968 46325
rect 22652 46316 22704 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 6000 46112 6052 46164
rect 9220 46112 9272 46164
rect 10692 46155 10744 46164
rect 10692 46121 10701 46155
rect 10701 46121 10735 46155
rect 10735 46121 10744 46155
rect 10692 46112 10744 46121
rect 17408 46112 17460 46164
rect 19156 46112 19208 46164
rect 24492 46112 24544 46164
rect 25504 46112 25556 46164
rect 7656 46044 7708 46096
rect 9128 45976 9180 46028
rect 11888 46019 11940 46028
rect 11888 45985 11897 46019
rect 11897 45985 11931 46019
rect 11931 45985 11940 46019
rect 11888 45976 11940 45985
rect 12164 46019 12216 46028
rect 12164 45985 12173 46019
rect 12173 45985 12207 46019
rect 12207 45985 12216 46019
rect 12164 45976 12216 45985
rect 12624 45976 12676 46028
rect 14096 46019 14148 46028
rect 14096 45985 14105 46019
rect 14105 45985 14139 46019
rect 14139 45985 14148 46019
rect 14096 45976 14148 45985
rect 20168 46019 20220 46028
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 20444 45976 20496 46028
rect 21364 46019 21416 46028
rect 21364 45985 21373 46019
rect 21373 45985 21407 46019
rect 21407 45985 21416 46019
rect 21364 45976 21416 45985
rect 21456 46019 21508 46028
rect 21456 45985 21465 46019
rect 21465 45985 21499 46019
rect 21499 45985 21508 46019
rect 21456 45976 21508 45985
rect 1308 45908 1360 45960
rect 7472 45908 7524 45960
rect 10048 45908 10100 45960
rect 6920 45840 6972 45892
rect 11704 45840 11756 45892
rect 12624 45840 12676 45892
rect 19616 45840 19668 45892
rect 11152 45815 11204 45824
rect 11152 45781 11161 45815
rect 11161 45781 11195 45815
rect 11195 45781 11204 45815
rect 11152 45772 11204 45781
rect 13452 45772 13504 45824
rect 16396 45815 16448 45824
rect 16396 45781 16405 45815
rect 16405 45781 16439 45815
rect 16439 45781 16448 45815
rect 16396 45772 16448 45781
rect 19892 45772 19944 45824
rect 20076 45815 20128 45824
rect 20076 45781 20085 45815
rect 20085 45781 20119 45815
rect 20119 45781 20128 45815
rect 20076 45772 20128 45781
rect 20996 45772 21048 45824
rect 21272 45815 21324 45824
rect 21272 45781 21281 45815
rect 21281 45781 21315 45815
rect 21315 45781 21324 45815
rect 21272 45772 21324 45781
rect 23664 45908 23716 45960
rect 24860 45772 24912 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 1308 45568 1360 45620
rect 16396 45611 16448 45620
rect 8852 45543 8904 45552
rect 8852 45509 8861 45543
rect 8861 45509 8895 45543
rect 8895 45509 8904 45543
rect 8852 45500 8904 45509
rect 9772 45500 9824 45552
rect 14096 45500 14148 45552
rect 16396 45577 16405 45611
rect 16405 45577 16439 45611
rect 16439 45577 16448 45611
rect 16396 45568 16448 45577
rect 19340 45568 19392 45620
rect 15108 45500 15160 45552
rect 19156 45500 19208 45552
rect 21456 45500 21508 45552
rect 9220 45475 9272 45484
rect 9220 45441 9229 45475
rect 9229 45441 9263 45475
rect 9263 45441 9272 45475
rect 9220 45432 9272 45441
rect 10600 45432 10652 45484
rect 23572 45432 23624 45484
rect 24124 45432 24176 45484
rect 9864 45364 9916 45416
rect 12164 45364 12216 45416
rect 14372 45407 14424 45416
rect 14372 45373 14381 45407
rect 14381 45373 14415 45407
rect 14415 45373 14424 45407
rect 14372 45364 14424 45373
rect 16304 45364 16356 45416
rect 18328 45364 18380 45416
rect 20076 45364 20128 45416
rect 20260 45364 20312 45416
rect 21088 45364 21140 45416
rect 10508 45296 10560 45348
rect 12348 45228 12400 45280
rect 16120 45271 16172 45280
rect 16120 45237 16129 45271
rect 16129 45237 16163 45271
rect 16163 45237 16172 45271
rect 16120 45228 16172 45237
rect 18880 45228 18932 45280
rect 20904 45296 20956 45348
rect 21272 45296 21324 45348
rect 24492 45407 24544 45416
rect 24492 45373 24501 45407
rect 24501 45373 24535 45407
rect 24535 45373 24544 45407
rect 24492 45364 24544 45373
rect 23388 45296 23440 45348
rect 22284 45228 22336 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 7380 45024 7432 45076
rect 11244 45024 11296 45076
rect 12072 45024 12124 45076
rect 12808 45024 12860 45076
rect 4712 44956 4764 45008
rect 14372 44956 14424 45008
rect 16672 45024 16724 45076
rect 16948 45024 17000 45076
rect 12624 44888 12676 44940
rect 13728 44888 13780 44940
rect 17684 44956 17736 45008
rect 16764 44888 16816 44940
rect 23020 44888 23072 44940
rect 23572 44888 23624 44940
rect 12348 44863 12400 44872
rect 12348 44829 12357 44863
rect 12357 44829 12391 44863
rect 12391 44829 12400 44863
rect 12348 44820 12400 44829
rect 14372 44820 14424 44872
rect 19524 44863 19576 44872
rect 19524 44829 19533 44863
rect 19533 44829 19567 44863
rect 19567 44829 19576 44863
rect 19524 44820 19576 44829
rect 21088 44820 21140 44872
rect 6644 44684 6696 44736
rect 7104 44727 7156 44736
rect 7104 44693 7113 44727
rect 7113 44693 7147 44727
rect 7147 44693 7156 44727
rect 7104 44684 7156 44693
rect 12532 44752 12584 44804
rect 15108 44752 15160 44804
rect 8484 44684 8536 44736
rect 9772 44727 9824 44736
rect 9772 44693 9781 44727
rect 9781 44693 9815 44727
rect 9815 44693 9824 44727
rect 9772 44684 9824 44693
rect 13360 44727 13412 44736
rect 13360 44693 13369 44727
rect 13369 44693 13403 44727
rect 13403 44693 13412 44727
rect 13360 44684 13412 44693
rect 15292 44684 15344 44736
rect 19800 44795 19852 44804
rect 19800 44761 19809 44795
rect 19809 44761 19843 44795
rect 19843 44761 19852 44795
rect 19800 44752 19852 44761
rect 20260 44752 20312 44804
rect 17132 44727 17184 44736
rect 17132 44693 17141 44727
rect 17141 44693 17175 44727
rect 17175 44693 17184 44727
rect 17132 44684 17184 44693
rect 21272 44727 21324 44736
rect 21272 44693 21281 44727
rect 21281 44693 21315 44727
rect 21315 44693 21324 44727
rect 21272 44684 21324 44693
rect 22284 44863 22336 44872
rect 22284 44829 22293 44863
rect 22293 44829 22327 44863
rect 22327 44829 22336 44863
rect 22284 44820 22336 44829
rect 22560 44795 22612 44804
rect 22560 44761 22569 44795
rect 22569 44761 22603 44795
rect 22603 44761 22612 44795
rect 22560 44752 22612 44761
rect 23020 44752 23072 44804
rect 23388 44684 23440 44736
rect 24492 44684 24544 44736
rect 25504 44727 25556 44736
rect 25504 44693 25513 44727
rect 25513 44693 25547 44727
rect 25547 44693 25556 44727
rect 25504 44684 25556 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 5816 44523 5868 44532
rect 5816 44489 5825 44523
rect 5825 44489 5859 44523
rect 5859 44489 5868 44523
rect 5816 44480 5868 44489
rect 6736 44523 6788 44532
rect 6736 44489 6745 44523
rect 6745 44489 6779 44523
rect 6779 44489 6788 44523
rect 6736 44480 6788 44489
rect 7840 44480 7892 44532
rect 9680 44480 9732 44532
rect 11152 44480 11204 44532
rect 14464 44480 14516 44532
rect 15108 44480 15160 44532
rect 7564 44455 7616 44464
rect 7564 44421 7573 44455
rect 7573 44421 7607 44455
rect 7607 44421 7616 44455
rect 7564 44412 7616 44421
rect 12348 44412 12400 44464
rect 12716 44412 12768 44464
rect 13452 44455 13504 44464
rect 13452 44421 13461 44455
rect 13461 44421 13495 44455
rect 13495 44421 13504 44455
rect 13452 44412 13504 44421
rect 14096 44412 14148 44464
rect 17132 44412 17184 44464
rect 18604 44523 18656 44532
rect 18604 44489 18613 44523
rect 18613 44489 18647 44523
rect 18647 44489 18656 44523
rect 18604 44480 18656 44489
rect 18788 44480 18840 44532
rect 19800 44480 19852 44532
rect 20444 44480 20496 44532
rect 22560 44480 22612 44532
rect 20260 44412 20312 44464
rect 21088 44412 21140 44464
rect 23020 44412 23072 44464
rect 5264 44344 5316 44396
rect 6736 44344 6788 44396
rect 7104 44344 7156 44396
rect 7472 44344 7524 44396
rect 7196 44276 7248 44328
rect 11612 44344 11664 44396
rect 11152 44276 11204 44328
rect 9496 44251 9548 44260
rect 9496 44217 9505 44251
rect 9505 44217 9539 44251
rect 9539 44217 9548 44251
rect 9496 44208 9548 44217
rect 12164 44208 12216 44260
rect 11612 44183 11664 44192
rect 11612 44149 11621 44183
rect 11621 44149 11655 44183
rect 11655 44149 11664 44183
rect 11612 44140 11664 44149
rect 25320 44344 25372 44396
rect 13452 44276 13504 44328
rect 16672 44276 16724 44328
rect 16764 44276 16816 44328
rect 18972 44276 19024 44328
rect 19524 44319 19576 44328
rect 19524 44285 19533 44319
rect 19533 44285 19567 44319
rect 19567 44285 19576 44319
rect 19524 44276 19576 44285
rect 21180 44276 21232 44328
rect 22284 44319 22336 44328
rect 22284 44285 22293 44319
rect 22293 44285 22327 44319
rect 22327 44285 22336 44319
rect 22284 44276 22336 44285
rect 22928 44276 22980 44328
rect 24768 44319 24820 44328
rect 24768 44285 24777 44319
rect 24777 44285 24811 44319
rect 24811 44285 24820 44319
rect 24768 44276 24820 44285
rect 14556 44140 14608 44192
rect 23296 44140 23348 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 9404 43936 9456 43988
rect 9956 43936 10008 43988
rect 18420 43936 18472 43988
rect 21548 43936 21600 43988
rect 23296 43936 23348 43988
rect 23480 43936 23532 43988
rect 23572 43936 23624 43988
rect 24216 43936 24268 43988
rect 7012 43868 7064 43920
rect 16856 43868 16908 43920
rect 9404 43800 9456 43852
rect 9496 43800 9548 43852
rect 18420 43800 18472 43852
rect 22192 43800 22244 43852
rect 23296 43800 23348 43852
rect 9036 43732 9088 43784
rect 8760 43596 8812 43648
rect 10692 43664 10744 43716
rect 10876 43639 10928 43648
rect 10876 43605 10885 43639
rect 10885 43605 10919 43639
rect 10919 43605 10928 43639
rect 10876 43596 10928 43605
rect 11428 43664 11480 43716
rect 21548 43664 21600 43716
rect 16396 43596 16448 43648
rect 17408 43596 17460 43648
rect 19340 43596 19392 43648
rect 21916 43596 21968 43648
rect 25320 43639 25372 43648
rect 25320 43605 25329 43639
rect 25329 43605 25363 43639
rect 25363 43605 25372 43639
rect 25320 43596 25372 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 7748 43435 7800 43444
rect 7748 43401 7757 43435
rect 7757 43401 7791 43435
rect 7791 43401 7800 43435
rect 7748 43392 7800 43401
rect 5356 43324 5408 43376
rect 8668 43392 8720 43444
rect 10416 43392 10468 43444
rect 14740 43392 14792 43444
rect 15568 43392 15620 43444
rect 17408 43435 17460 43444
rect 17408 43401 17417 43435
rect 17417 43401 17451 43435
rect 17451 43401 17460 43435
rect 17408 43392 17460 43401
rect 17500 43435 17552 43444
rect 17500 43401 17509 43435
rect 17509 43401 17543 43435
rect 17543 43401 17552 43435
rect 17500 43392 17552 43401
rect 20076 43435 20128 43444
rect 20076 43401 20085 43435
rect 20085 43401 20119 43435
rect 20119 43401 20128 43435
rect 20076 43392 20128 43401
rect 9128 43324 9180 43376
rect 10692 43324 10744 43376
rect 10968 43324 11020 43376
rect 12624 43367 12676 43376
rect 12624 43333 12633 43367
rect 12633 43333 12667 43367
rect 12667 43333 12676 43367
rect 12624 43324 12676 43333
rect 14096 43324 14148 43376
rect 16212 43324 16264 43376
rect 20904 43392 20956 43444
rect 21088 43392 21140 43444
rect 21640 43435 21692 43444
rect 21640 43401 21649 43435
rect 21649 43401 21683 43435
rect 21683 43401 21692 43435
rect 21640 43392 21692 43401
rect 1308 43256 1360 43308
rect 7656 43256 7708 43308
rect 8392 43256 8444 43308
rect 8760 43256 8812 43308
rect 9772 43256 9824 43308
rect 10324 43256 10376 43308
rect 14648 43256 14700 43308
rect 22376 43392 22428 43444
rect 24216 43392 24268 43444
rect 22192 43324 22244 43376
rect 22744 43324 22796 43376
rect 23572 43324 23624 43376
rect 8852 43188 8904 43240
rect 9312 43188 9364 43240
rect 9496 43188 9548 43240
rect 12348 43231 12400 43240
rect 12348 43197 12357 43231
rect 12357 43197 12391 43231
rect 12391 43197 12400 43231
rect 12348 43188 12400 43197
rect 15660 43188 15712 43240
rect 17684 43231 17736 43240
rect 17684 43197 17693 43231
rect 17693 43197 17727 43231
rect 17727 43197 17736 43231
rect 17684 43188 17736 43197
rect 18328 43231 18380 43240
rect 18328 43197 18337 43231
rect 18337 43197 18371 43231
rect 18371 43197 18380 43231
rect 18328 43188 18380 43197
rect 19616 43188 19668 43240
rect 21272 43188 21324 43240
rect 22744 43188 22796 43240
rect 23480 43188 23532 43240
rect 3976 43120 4028 43172
rect 11152 43120 11204 43172
rect 13728 43120 13780 43172
rect 16764 43120 16816 43172
rect 13912 43052 13964 43104
rect 17040 43095 17092 43104
rect 17040 43061 17049 43095
rect 17049 43061 17083 43095
rect 17083 43061 17092 43095
rect 17040 43052 17092 43061
rect 19248 43052 19300 43104
rect 24952 43052 25004 43104
rect 25136 43052 25188 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 8668 42891 8720 42900
rect 8668 42857 8677 42891
rect 8677 42857 8711 42891
rect 8711 42857 8720 42891
rect 8668 42848 8720 42857
rect 8852 42848 8904 42900
rect 9128 42891 9180 42900
rect 9128 42857 9137 42891
rect 9137 42857 9171 42891
rect 9171 42857 9180 42891
rect 9128 42848 9180 42857
rect 9496 42848 9548 42900
rect 10692 42848 10744 42900
rect 4896 42712 4948 42764
rect 9128 42712 9180 42764
rect 9220 42712 9272 42764
rect 9404 42712 9456 42764
rect 12348 42712 12400 42764
rect 14096 42848 14148 42900
rect 20352 42848 20404 42900
rect 21456 42848 21508 42900
rect 24216 42848 24268 42900
rect 21640 42780 21692 42832
rect 16764 42712 16816 42764
rect 18420 42712 18472 42764
rect 16212 42644 16264 42696
rect 18604 42644 18656 42696
rect 19064 42644 19116 42696
rect 20904 42644 20956 42696
rect 22008 42712 22060 42764
rect 22560 42712 22612 42764
rect 23112 42712 23164 42764
rect 24860 42712 24912 42764
rect 22836 42644 22888 42696
rect 4804 42619 4856 42628
rect 4804 42585 4813 42619
rect 4813 42585 4847 42619
rect 4847 42585 4856 42619
rect 4804 42576 4856 42585
rect 9680 42576 9732 42628
rect 8392 42508 8444 42560
rect 10324 42551 10376 42560
rect 10324 42517 10333 42551
rect 10333 42517 10367 42551
rect 10367 42517 10376 42551
rect 10324 42508 10376 42517
rect 12440 42508 12492 42560
rect 14556 42508 14608 42560
rect 16764 42508 16816 42560
rect 21088 42576 21140 42628
rect 20444 42508 20496 42560
rect 21272 42551 21324 42560
rect 21272 42517 21281 42551
rect 21281 42517 21315 42551
rect 21315 42517 21324 42551
rect 21272 42508 21324 42517
rect 22100 42508 22152 42560
rect 24860 42508 24912 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 4160 42304 4212 42356
rect 5080 42347 5132 42356
rect 5080 42313 5089 42347
rect 5089 42313 5123 42347
rect 5123 42313 5132 42347
rect 5080 42304 5132 42313
rect 5448 42304 5500 42356
rect 8116 42304 8168 42356
rect 9220 42304 9272 42356
rect 9588 42304 9640 42356
rect 11796 42347 11848 42356
rect 11796 42313 11805 42347
rect 11805 42313 11839 42347
rect 11839 42313 11848 42347
rect 11796 42304 11848 42313
rect 13360 42304 13412 42356
rect 15292 42304 15344 42356
rect 20536 42304 20588 42356
rect 20904 42304 20956 42356
rect 22376 42304 22428 42356
rect 23296 42304 23348 42356
rect 4252 42211 4304 42220
rect 4252 42177 4261 42211
rect 4261 42177 4295 42211
rect 4295 42177 4304 42211
rect 4252 42168 4304 42177
rect 7196 42168 7248 42220
rect 9128 42236 9180 42288
rect 11888 42236 11940 42288
rect 15568 42236 15620 42288
rect 17408 42236 17460 42288
rect 7748 42143 7800 42152
rect 7748 42109 7757 42143
rect 7757 42109 7791 42143
rect 7791 42109 7800 42143
rect 9588 42168 9640 42220
rect 11152 42168 11204 42220
rect 16672 42168 16724 42220
rect 20720 42236 20772 42288
rect 24216 42236 24268 42288
rect 7748 42100 7800 42109
rect 6368 41964 6420 42016
rect 7196 42007 7248 42016
rect 7196 41973 7205 42007
rect 7205 41973 7239 42007
rect 7239 41973 7248 42007
rect 7196 41964 7248 41973
rect 7564 41964 7616 42016
rect 9588 42032 9640 42084
rect 12440 42143 12492 42152
rect 12440 42109 12449 42143
rect 12449 42109 12483 42143
rect 12483 42109 12492 42143
rect 12440 42100 12492 42109
rect 14464 42100 14516 42152
rect 20628 42211 20680 42220
rect 20628 42177 20637 42211
rect 20637 42177 20671 42211
rect 20671 42177 20680 42211
rect 20628 42168 20680 42177
rect 13360 42032 13412 42084
rect 9680 41964 9732 42016
rect 10508 41964 10560 42016
rect 14464 41964 14516 42016
rect 19064 42100 19116 42152
rect 19248 42100 19300 42152
rect 20996 42168 21048 42220
rect 19708 42032 19760 42084
rect 21272 42100 21324 42152
rect 22836 42143 22888 42152
rect 22836 42109 22845 42143
rect 22845 42109 22879 42143
rect 22879 42109 22888 42143
rect 23480 42143 23532 42152
rect 22836 42100 22888 42109
rect 23480 42109 23489 42143
rect 23489 42109 23523 42143
rect 23523 42109 23532 42143
rect 23480 42100 23532 42109
rect 25136 42100 25188 42152
rect 20260 42007 20312 42016
rect 20260 41973 20269 42007
rect 20269 41973 20303 42007
rect 20303 41973 20312 42007
rect 20260 41964 20312 41973
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 5172 41803 5224 41812
rect 5172 41769 5181 41803
rect 5181 41769 5215 41803
rect 5215 41769 5224 41803
rect 5172 41760 5224 41769
rect 7748 41760 7800 41812
rect 7840 41760 7892 41812
rect 8116 41803 8168 41812
rect 8116 41769 8125 41803
rect 8125 41769 8159 41803
rect 8159 41769 8168 41803
rect 8116 41760 8168 41769
rect 11060 41760 11112 41812
rect 6184 41624 6236 41676
rect 8300 41692 8352 41744
rect 9128 41692 9180 41744
rect 15292 41692 15344 41744
rect 16120 41692 16172 41744
rect 9220 41624 9272 41676
rect 10600 41624 10652 41676
rect 10784 41624 10836 41676
rect 12348 41624 12400 41676
rect 12808 41667 12860 41676
rect 12808 41633 12817 41667
rect 12817 41633 12851 41667
rect 12851 41633 12860 41667
rect 12808 41624 12860 41633
rect 16580 41624 16632 41676
rect 10508 41556 10560 41608
rect 5908 41420 5960 41472
rect 14004 41488 14056 41540
rect 22928 41760 22980 41812
rect 24216 41760 24268 41812
rect 17776 41692 17828 41744
rect 18512 41624 18564 41676
rect 21180 41735 21232 41744
rect 21180 41701 21189 41735
rect 21189 41701 21223 41735
rect 21223 41701 21232 41735
rect 21180 41692 21232 41701
rect 22560 41692 22612 41744
rect 25044 41692 25096 41744
rect 25412 41692 25464 41744
rect 18972 41624 19024 41676
rect 19708 41667 19760 41676
rect 19708 41633 19717 41667
rect 19717 41633 19751 41667
rect 19751 41633 19760 41667
rect 19708 41624 19760 41633
rect 7748 41420 7800 41472
rect 9680 41420 9732 41472
rect 10784 41420 10836 41472
rect 11060 41463 11112 41472
rect 11060 41429 11069 41463
rect 11069 41429 11103 41463
rect 11103 41429 11112 41463
rect 11060 41420 11112 41429
rect 12808 41420 12860 41472
rect 13636 41420 13688 41472
rect 16212 41463 16264 41472
rect 16212 41429 16221 41463
rect 16221 41429 16255 41463
rect 16255 41429 16264 41463
rect 16212 41420 16264 41429
rect 16488 41420 16540 41472
rect 19248 41556 19300 41608
rect 20904 41624 20956 41676
rect 22468 41624 22520 41676
rect 22652 41624 22704 41676
rect 23480 41624 23532 41676
rect 25320 41599 25372 41608
rect 25320 41565 25329 41599
rect 25329 41565 25363 41599
rect 25363 41565 25372 41599
rect 25320 41556 25372 41565
rect 19156 41488 19208 41540
rect 20996 41488 21048 41540
rect 22192 41488 22244 41540
rect 18420 41420 18472 41472
rect 19984 41420 20036 41472
rect 21640 41420 21692 41472
rect 22008 41463 22060 41472
rect 22008 41429 22017 41463
rect 22017 41429 22051 41463
rect 22051 41429 22060 41463
rect 22008 41420 22060 41429
rect 24860 41463 24912 41472
rect 24860 41429 24869 41463
rect 24869 41429 24903 41463
rect 24903 41429 24912 41463
rect 24860 41420 24912 41429
rect 25320 41420 25372 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 1952 41216 2004 41268
rect 6184 41216 6236 41268
rect 7840 41216 7892 41268
rect 1308 41080 1360 41132
rect 4620 41080 4672 41132
rect 9404 41216 9456 41268
rect 10968 41259 11020 41268
rect 10968 41225 10977 41259
rect 10977 41225 11011 41259
rect 11011 41225 11020 41259
rect 10968 41216 11020 41225
rect 11704 41259 11756 41268
rect 11704 41225 11713 41259
rect 11713 41225 11747 41259
rect 11747 41225 11756 41259
rect 11704 41216 11756 41225
rect 15384 41148 15436 41200
rect 16120 41216 16172 41268
rect 19892 41259 19944 41268
rect 19892 41225 19901 41259
rect 19901 41225 19935 41259
rect 19935 41225 19944 41259
rect 19892 41216 19944 41225
rect 20168 41216 20220 41268
rect 20444 41216 20496 41268
rect 20812 41216 20864 41268
rect 20996 41216 21048 41268
rect 21456 41216 21508 41268
rect 22008 41259 22060 41268
rect 22008 41225 22017 41259
rect 22017 41225 22051 41259
rect 22051 41225 22060 41259
rect 22008 41216 22060 41225
rect 23480 41216 23532 41268
rect 10508 41080 10560 41132
rect 12348 41080 12400 41132
rect 13636 41123 13688 41132
rect 13636 41089 13645 41123
rect 13645 41089 13679 41123
rect 13679 41089 13688 41123
rect 13636 41080 13688 41089
rect 16672 41080 16724 41132
rect 9220 41055 9272 41064
rect 9220 41021 9229 41055
rect 9229 41021 9263 41055
rect 9263 41021 9272 41055
rect 9220 41012 9272 41021
rect 12256 41055 12308 41064
rect 12256 41021 12265 41055
rect 12265 41021 12299 41055
rect 12299 41021 12308 41055
rect 12256 41012 12308 41021
rect 14004 41012 14056 41064
rect 15292 41012 15344 41064
rect 16764 41012 16816 41064
rect 21272 41148 21324 41200
rect 22284 41148 22336 41200
rect 23204 41191 23256 41200
rect 23204 41157 23213 41191
rect 23213 41157 23247 41191
rect 23247 41157 23256 41191
rect 23204 41148 23256 41157
rect 24216 41148 24268 41200
rect 19800 41123 19852 41132
rect 19800 41089 19809 41123
rect 19809 41089 19843 41123
rect 19843 41089 19852 41123
rect 19800 41080 19852 41089
rect 19616 41012 19668 41064
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 20996 41012 21048 41064
rect 21272 41055 21324 41064
rect 21272 41021 21281 41055
rect 21281 41021 21315 41055
rect 21315 41021 21324 41055
rect 21272 41012 21324 41021
rect 15752 40944 15804 40996
rect 18328 40944 18380 40996
rect 18972 40944 19024 40996
rect 19984 40944 20036 40996
rect 22468 41012 22520 41064
rect 22836 41012 22888 41064
rect 23204 41012 23256 41064
rect 24860 41012 24912 41064
rect 1676 40876 1728 40928
rect 9956 40876 10008 40928
rect 10692 40919 10744 40928
rect 10692 40885 10701 40919
rect 10701 40885 10735 40919
rect 10735 40885 10744 40919
rect 10692 40876 10744 40885
rect 18512 40876 18564 40928
rect 19156 40919 19208 40928
rect 19156 40885 19165 40919
rect 19165 40885 19199 40919
rect 19199 40885 19208 40919
rect 19156 40876 19208 40885
rect 19432 40919 19484 40928
rect 19432 40885 19441 40919
rect 19441 40885 19475 40919
rect 19475 40885 19484 40919
rect 19432 40876 19484 40885
rect 19524 40876 19576 40928
rect 20812 40876 20864 40928
rect 21456 40876 21508 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 8576 40715 8628 40724
rect 8576 40681 8585 40715
rect 8585 40681 8619 40715
rect 8619 40681 8628 40715
rect 8576 40672 8628 40681
rect 8668 40672 8720 40724
rect 10232 40604 10284 40656
rect 10600 40715 10652 40724
rect 10600 40681 10609 40715
rect 10609 40681 10643 40715
rect 10643 40681 10652 40715
rect 10600 40672 10652 40681
rect 11244 40672 11296 40724
rect 13912 40672 13964 40724
rect 6552 40536 6604 40588
rect 6184 40511 6236 40520
rect 6184 40477 6193 40511
rect 6193 40477 6227 40511
rect 6227 40477 6236 40511
rect 6184 40468 6236 40477
rect 10324 40536 10376 40588
rect 13636 40536 13688 40588
rect 15844 40579 15896 40588
rect 15844 40545 15853 40579
rect 15853 40545 15887 40579
rect 15887 40545 15896 40579
rect 15844 40536 15896 40545
rect 12440 40468 12492 40520
rect 19524 40672 19576 40724
rect 19616 40672 19668 40724
rect 21088 40672 21140 40724
rect 16948 40604 17000 40656
rect 17040 40536 17092 40588
rect 17316 40604 17368 40656
rect 20168 40604 20220 40656
rect 22560 40672 22612 40724
rect 23020 40672 23072 40724
rect 24216 40672 24268 40724
rect 19616 40536 19668 40588
rect 16580 40468 16632 40520
rect 19156 40468 19208 40520
rect 22100 40536 22152 40588
rect 23388 40536 23440 40588
rect 8576 40400 8628 40452
rect 11244 40400 11296 40452
rect 12256 40400 12308 40452
rect 15936 40400 15988 40452
rect 7288 40332 7340 40384
rect 7748 40332 7800 40384
rect 8300 40375 8352 40384
rect 8300 40341 8309 40375
rect 8309 40341 8343 40375
rect 8343 40341 8352 40375
rect 8300 40332 8352 40341
rect 9496 40332 9548 40384
rect 10324 40375 10376 40384
rect 10324 40341 10333 40375
rect 10333 40341 10367 40375
rect 10367 40341 10376 40375
rect 10324 40332 10376 40341
rect 12164 40375 12216 40384
rect 12164 40341 12173 40375
rect 12173 40341 12207 40375
rect 12207 40341 12216 40375
rect 12164 40332 12216 40341
rect 12624 40375 12676 40384
rect 12624 40341 12633 40375
rect 12633 40341 12667 40375
rect 12667 40341 12676 40375
rect 12624 40332 12676 40341
rect 15384 40332 15436 40384
rect 17500 40400 17552 40452
rect 22468 40468 22520 40520
rect 23020 40468 23072 40520
rect 25320 40511 25372 40520
rect 25320 40477 25329 40511
rect 25329 40477 25363 40511
rect 25363 40477 25372 40511
rect 25320 40468 25372 40477
rect 21732 40400 21784 40452
rect 22008 40400 22060 40452
rect 17040 40375 17092 40384
rect 17040 40341 17049 40375
rect 17049 40341 17083 40375
rect 17083 40341 17092 40375
rect 17040 40332 17092 40341
rect 19800 40332 19852 40384
rect 20444 40332 20496 40384
rect 21272 40375 21324 40384
rect 21272 40341 21281 40375
rect 21281 40341 21315 40375
rect 21315 40341 21324 40375
rect 21272 40332 21324 40341
rect 22652 40332 22704 40384
rect 24768 40400 24820 40452
rect 25228 40400 25280 40452
rect 22928 40332 22980 40384
rect 25780 40332 25832 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 7380 40128 7432 40180
rect 8760 40128 8812 40180
rect 10324 40128 10376 40180
rect 7840 40060 7892 40112
rect 7932 40060 7984 40112
rect 8300 40060 8352 40112
rect 10968 40128 11020 40180
rect 11704 40128 11756 40180
rect 12256 40171 12308 40180
rect 12256 40137 12265 40171
rect 12265 40137 12299 40171
rect 12299 40137 12308 40171
rect 12256 40128 12308 40137
rect 14556 40060 14608 40112
rect 15292 40060 15344 40112
rect 15568 40171 15620 40180
rect 15568 40137 15577 40171
rect 15577 40137 15611 40171
rect 15611 40137 15620 40171
rect 15568 40128 15620 40137
rect 16304 40060 16356 40112
rect 18236 40171 18288 40180
rect 18236 40137 18245 40171
rect 18245 40137 18279 40171
rect 18279 40137 18288 40171
rect 18236 40128 18288 40137
rect 18420 40128 18472 40180
rect 20628 40128 20680 40180
rect 22468 40128 22520 40180
rect 23296 40128 23348 40180
rect 18328 40060 18380 40112
rect 7380 39992 7432 40044
rect 12808 39992 12860 40044
rect 18420 39992 18472 40044
rect 7748 39967 7800 39976
rect 7748 39933 7757 39967
rect 7757 39933 7791 39967
rect 7791 39933 7800 39967
rect 7748 39924 7800 39933
rect 7840 39967 7892 39976
rect 7840 39933 7849 39967
rect 7849 39933 7883 39967
rect 7883 39933 7892 39967
rect 7840 39924 7892 39933
rect 9956 39924 10008 39976
rect 10968 39967 11020 39976
rect 10968 39933 10977 39967
rect 10977 39933 11011 39967
rect 11011 39933 11020 39967
rect 10968 39924 11020 39933
rect 15752 39924 15804 39976
rect 16028 39967 16080 39976
rect 16028 39933 16037 39967
rect 16037 39933 16071 39967
rect 16071 39933 16080 39967
rect 16028 39924 16080 39933
rect 16120 39967 16172 39976
rect 16120 39933 16129 39967
rect 16129 39933 16163 39967
rect 16163 39933 16172 39967
rect 16120 39924 16172 39933
rect 18788 39967 18840 39976
rect 18788 39933 18797 39967
rect 18797 39933 18831 39967
rect 18831 39933 18840 39967
rect 18788 39924 18840 39933
rect 10048 39856 10100 39908
rect 12716 39856 12768 39908
rect 17132 39856 17184 39908
rect 19984 39992 20036 40044
rect 20444 40060 20496 40112
rect 19340 39924 19392 39976
rect 19708 39924 19760 39976
rect 20352 39967 20404 39976
rect 20352 39933 20361 39967
rect 20361 39933 20395 39967
rect 20395 39933 20404 39967
rect 20352 39924 20404 39933
rect 21732 39992 21784 40044
rect 22836 40060 22888 40112
rect 22928 39992 22980 40044
rect 24216 40060 24268 40112
rect 19064 39856 19116 39908
rect 23388 39924 23440 39976
rect 24492 39924 24544 39976
rect 7104 39788 7156 39840
rect 10692 39788 10744 39840
rect 14648 39831 14700 39840
rect 14648 39797 14657 39831
rect 14657 39797 14691 39831
rect 14691 39797 14700 39831
rect 14648 39788 14700 39797
rect 16304 39788 16356 39840
rect 19984 39788 20036 39840
rect 20628 39788 20680 39840
rect 22836 39856 22888 39908
rect 25596 39788 25648 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 6552 39584 6604 39636
rect 7748 39584 7800 39636
rect 10784 39584 10836 39636
rect 16120 39584 16172 39636
rect 18604 39584 18656 39636
rect 19064 39627 19116 39636
rect 19064 39593 19073 39627
rect 19073 39593 19107 39627
rect 19107 39593 19116 39627
rect 19064 39584 19116 39593
rect 22192 39584 22244 39636
rect 12716 39516 12768 39568
rect 16028 39516 16080 39568
rect 25412 39584 25464 39636
rect 6184 39448 6236 39500
rect 10232 39491 10284 39500
rect 10232 39457 10241 39491
rect 10241 39457 10275 39491
rect 10275 39457 10284 39491
rect 10232 39448 10284 39457
rect 8576 39380 8628 39432
rect 12440 39448 12492 39500
rect 12808 39448 12860 39500
rect 13820 39448 13872 39500
rect 15660 39448 15712 39500
rect 17684 39448 17736 39500
rect 19432 39448 19484 39500
rect 20076 39491 20128 39500
rect 20076 39457 20085 39491
rect 20085 39457 20119 39491
rect 20119 39457 20128 39491
rect 20076 39448 20128 39457
rect 21732 39491 21784 39500
rect 21732 39457 21741 39491
rect 21741 39457 21775 39491
rect 21775 39457 21784 39491
rect 21732 39448 21784 39457
rect 12900 39380 12952 39432
rect 14280 39380 14332 39432
rect 14556 39380 14608 39432
rect 7932 39312 7984 39364
rect 11244 39355 11296 39364
rect 11244 39321 11253 39355
rect 11253 39321 11287 39355
rect 11287 39321 11296 39355
rect 11244 39312 11296 39321
rect 15016 39312 15068 39364
rect 5816 39244 5868 39296
rect 7012 39287 7064 39296
rect 7012 39253 7021 39287
rect 7021 39253 7055 39287
rect 7055 39253 7064 39287
rect 7012 39244 7064 39253
rect 8300 39244 8352 39296
rect 10140 39287 10192 39296
rect 10140 39253 10149 39287
rect 10149 39253 10183 39287
rect 10183 39253 10192 39287
rect 10140 39244 10192 39253
rect 12716 39287 12768 39296
rect 12716 39253 12725 39287
rect 12725 39253 12759 39287
rect 12759 39253 12768 39287
rect 12716 39244 12768 39253
rect 13084 39244 13136 39296
rect 13912 39244 13964 39296
rect 17040 39312 17092 39364
rect 17224 39312 17276 39364
rect 21272 39380 21324 39432
rect 18788 39312 18840 39364
rect 15476 39244 15528 39296
rect 16028 39287 16080 39296
rect 16028 39253 16037 39287
rect 16037 39253 16071 39287
rect 16071 39253 16080 39287
rect 16028 39244 16080 39253
rect 18420 39244 18472 39296
rect 18696 39244 18748 39296
rect 20352 39244 20404 39296
rect 20444 39287 20496 39296
rect 20444 39253 20453 39287
rect 20453 39253 20487 39287
rect 20487 39253 20496 39287
rect 20444 39244 20496 39253
rect 20628 39244 20680 39296
rect 21088 39244 21140 39296
rect 21824 39244 21876 39296
rect 23480 39448 23532 39500
rect 22008 39380 22060 39432
rect 25044 39491 25096 39500
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 25136 39491 25188 39500
rect 25136 39457 25145 39491
rect 25145 39457 25179 39491
rect 25179 39457 25188 39491
rect 25136 39448 25188 39457
rect 22284 39287 22336 39296
rect 22284 39253 22293 39287
rect 22293 39253 22327 39287
rect 22327 39253 22336 39287
rect 22284 39244 22336 39253
rect 24308 39244 24360 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 8668 39040 8720 39092
rect 10968 39040 11020 39092
rect 4068 38972 4120 39024
rect 12256 39040 12308 39092
rect 12992 39040 13044 39092
rect 8392 38904 8444 38956
rect 8668 38904 8720 38956
rect 6736 38836 6788 38888
rect 8484 38836 8536 38888
rect 7012 38700 7064 38752
rect 7748 38700 7800 38752
rect 8392 38700 8444 38752
rect 9588 38836 9640 38888
rect 10784 38904 10836 38956
rect 12440 38972 12492 39024
rect 12900 38972 12952 39024
rect 15016 39040 15068 39092
rect 15936 39040 15988 39092
rect 16028 39040 16080 39092
rect 20628 39040 20680 39092
rect 20996 39040 21048 39092
rect 14464 38972 14516 39024
rect 14832 38972 14884 39024
rect 17224 38972 17276 39024
rect 18604 38972 18656 39024
rect 20812 38972 20864 39024
rect 15660 38904 15712 38956
rect 19892 38904 19944 38956
rect 22376 39015 22428 39024
rect 22376 38981 22385 39015
rect 22385 38981 22419 39015
rect 22419 38981 22428 39015
rect 22376 38972 22428 38981
rect 24216 38972 24268 39024
rect 24860 38904 24912 38956
rect 25320 38947 25372 38956
rect 25320 38913 25329 38947
rect 25329 38913 25363 38947
rect 25363 38913 25372 38947
rect 25320 38904 25372 38913
rect 9128 38743 9180 38752
rect 9128 38709 9137 38743
rect 9137 38709 9171 38743
rect 9171 38709 9180 38743
rect 9128 38700 9180 38709
rect 14648 38836 14700 38888
rect 15568 38879 15620 38888
rect 15568 38845 15577 38879
rect 15577 38845 15611 38879
rect 15611 38845 15620 38879
rect 15568 38836 15620 38845
rect 16396 38836 16448 38888
rect 17224 38836 17276 38888
rect 18420 38879 18472 38888
rect 18420 38845 18429 38879
rect 18429 38845 18463 38879
rect 18463 38845 18472 38879
rect 18420 38836 18472 38845
rect 19156 38836 19208 38888
rect 11152 38768 11204 38820
rect 11244 38768 11296 38820
rect 11520 38743 11572 38752
rect 11520 38709 11529 38743
rect 11529 38709 11563 38743
rect 11563 38709 11572 38743
rect 11520 38700 11572 38709
rect 14004 38768 14056 38820
rect 18236 38768 18288 38820
rect 20444 38836 20496 38888
rect 19984 38768 20036 38820
rect 22100 38879 22152 38888
rect 22100 38845 22109 38879
rect 22109 38845 22143 38879
rect 22143 38845 22152 38879
rect 22100 38836 22152 38845
rect 22836 38836 22888 38888
rect 24216 38879 24268 38888
rect 24216 38845 24225 38879
rect 24225 38845 24259 38879
rect 24259 38845 24268 38879
rect 24216 38836 24268 38845
rect 25964 38836 26016 38888
rect 23388 38768 23440 38820
rect 25872 38768 25924 38820
rect 12072 38700 12124 38752
rect 13084 38700 13136 38752
rect 13912 38700 13964 38752
rect 18420 38700 18472 38752
rect 18512 38700 18564 38752
rect 18604 38700 18656 38752
rect 18972 38700 19024 38752
rect 21272 38700 21324 38752
rect 22560 38700 22612 38752
rect 25136 38743 25188 38752
rect 25136 38709 25145 38743
rect 25145 38709 25179 38743
rect 25179 38709 25188 38743
rect 25136 38700 25188 38709
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 7564 38496 7616 38548
rect 11060 38496 11112 38548
rect 11888 38539 11940 38548
rect 11888 38505 11897 38539
rect 11897 38505 11931 38539
rect 11931 38505 11940 38539
rect 11888 38496 11940 38505
rect 12348 38496 12400 38548
rect 12532 38496 12584 38548
rect 14188 38496 14240 38548
rect 17408 38496 17460 38548
rect 22192 38496 22244 38548
rect 22376 38496 22428 38548
rect 8576 38428 8628 38480
rect 9220 38428 9272 38480
rect 6920 38360 6972 38412
rect 7840 38360 7892 38412
rect 1308 38292 1360 38344
rect 1584 38199 1636 38208
rect 1584 38165 1593 38199
rect 1593 38165 1627 38199
rect 1627 38165 1636 38199
rect 1584 38156 1636 38165
rect 7288 38292 7340 38344
rect 7748 38224 7800 38276
rect 8300 38292 8352 38344
rect 9128 38360 9180 38412
rect 12716 38428 12768 38480
rect 9220 38292 9272 38344
rect 12164 38360 12216 38412
rect 10600 38292 10652 38344
rect 14280 38360 14332 38412
rect 17868 38428 17920 38480
rect 15016 38360 15068 38412
rect 18236 38360 18288 38412
rect 15384 38292 15436 38344
rect 15936 38335 15988 38344
rect 15936 38301 15945 38335
rect 15945 38301 15979 38335
rect 15979 38301 15988 38335
rect 15936 38292 15988 38301
rect 17592 38292 17644 38344
rect 20812 38428 20864 38480
rect 22744 38428 22796 38480
rect 18696 38403 18748 38412
rect 18696 38369 18705 38403
rect 18705 38369 18739 38403
rect 18739 38369 18748 38403
rect 18696 38360 18748 38369
rect 19248 38360 19300 38412
rect 20260 38360 20312 38412
rect 21180 38403 21232 38412
rect 21180 38369 21189 38403
rect 21189 38369 21223 38403
rect 21223 38369 21232 38403
rect 21180 38360 21232 38369
rect 21916 38360 21968 38412
rect 22560 38403 22612 38412
rect 22560 38369 22569 38403
rect 22569 38369 22603 38403
rect 22603 38369 22612 38403
rect 22560 38360 22612 38369
rect 23848 38360 23900 38412
rect 18972 38292 19024 38344
rect 6552 38156 6604 38208
rect 7104 38156 7156 38208
rect 8208 38156 8260 38208
rect 8484 38156 8536 38208
rect 9680 38224 9732 38276
rect 10600 38156 10652 38208
rect 10784 38199 10836 38208
rect 10784 38165 10793 38199
rect 10793 38165 10827 38199
rect 10827 38165 10836 38199
rect 10784 38156 10836 38165
rect 10876 38199 10928 38208
rect 10876 38165 10885 38199
rect 10885 38165 10919 38199
rect 10919 38165 10928 38199
rect 10876 38156 10928 38165
rect 12532 38156 12584 38208
rect 13268 38199 13320 38208
rect 13268 38165 13277 38199
rect 13277 38165 13311 38199
rect 13311 38165 13320 38199
rect 13268 38156 13320 38165
rect 13544 38156 13596 38208
rect 13820 38156 13872 38208
rect 19524 38224 19576 38276
rect 19892 38267 19944 38276
rect 19892 38233 19901 38267
rect 19901 38233 19935 38267
rect 19935 38233 19944 38267
rect 19892 38224 19944 38233
rect 17684 38199 17736 38208
rect 17684 38165 17693 38199
rect 17693 38165 17727 38199
rect 17727 38165 17736 38199
rect 17684 38156 17736 38165
rect 19064 38156 19116 38208
rect 20444 38156 20496 38208
rect 21088 38156 21140 38208
rect 24032 38292 24084 38344
rect 24952 38292 25004 38344
rect 23572 38267 23624 38276
rect 23572 38233 23581 38267
rect 23581 38233 23615 38267
rect 23615 38233 23624 38267
rect 23572 38224 23624 38233
rect 24216 38224 24268 38276
rect 23756 38156 23808 38208
rect 24676 38156 24728 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 5264 37995 5316 38004
rect 5264 37961 5273 37995
rect 5273 37961 5307 37995
rect 5307 37961 5316 37995
rect 5264 37952 5316 37961
rect 8944 37952 8996 38004
rect 9312 37952 9364 38004
rect 10508 37952 10560 38004
rect 10784 37952 10836 38004
rect 11796 37952 11848 38004
rect 13268 37952 13320 38004
rect 6920 37884 6972 37936
rect 7840 37884 7892 37936
rect 4988 37816 5040 37868
rect 11336 37927 11388 37936
rect 11336 37893 11345 37927
rect 11345 37893 11379 37927
rect 11379 37893 11388 37927
rect 11336 37884 11388 37893
rect 15384 37952 15436 38004
rect 16304 37952 16356 38004
rect 17224 37995 17276 38004
rect 17224 37961 17233 37995
rect 17233 37961 17267 37995
rect 17267 37961 17276 37995
rect 17224 37952 17276 37961
rect 17592 37952 17644 38004
rect 18696 37952 18748 38004
rect 20904 37952 20956 38004
rect 17868 37927 17920 37936
rect 5816 37791 5868 37800
rect 5816 37757 5825 37791
rect 5825 37757 5859 37791
rect 5859 37757 5868 37791
rect 5816 37748 5868 37757
rect 6552 37791 6604 37800
rect 6552 37757 6561 37791
rect 6561 37757 6595 37791
rect 6595 37757 6604 37791
rect 6552 37748 6604 37757
rect 7288 37748 7340 37800
rect 8392 37748 8444 37800
rect 10508 37791 10560 37800
rect 6644 37612 6696 37664
rect 10508 37757 10517 37791
rect 10517 37757 10551 37791
rect 10551 37757 10560 37791
rect 10508 37748 10560 37757
rect 11336 37680 11388 37732
rect 13452 37748 13504 37800
rect 13544 37791 13596 37800
rect 13544 37757 13553 37791
rect 13553 37757 13587 37791
rect 13587 37757 13596 37791
rect 13544 37748 13596 37757
rect 17868 37893 17877 37927
rect 17877 37893 17911 37927
rect 17911 37893 17920 37927
rect 17868 37884 17920 37893
rect 18236 37884 18288 37936
rect 19248 37884 19300 37936
rect 9588 37612 9640 37664
rect 15568 37748 15620 37800
rect 16120 37748 16172 37800
rect 14280 37680 14332 37732
rect 16396 37723 16448 37732
rect 16396 37689 16405 37723
rect 16405 37689 16439 37723
rect 16439 37689 16448 37723
rect 18604 37816 18656 37868
rect 20076 37884 20128 37936
rect 21088 37816 21140 37868
rect 17776 37748 17828 37800
rect 19616 37791 19668 37800
rect 19616 37757 19625 37791
rect 19625 37757 19659 37791
rect 19659 37757 19668 37791
rect 19616 37748 19668 37757
rect 21824 37952 21876 38004
rect 24676 37952 24728 38004
rect 23388 37884 23440 37936
rect 23848 37927 23900 37936
rect 23848 37893 23857 37927
rect 23857 37893 23891 37927
rect 23891 37893 23900 37927
rect 23848 37884 23900 37893
rect 24860 37884 24912 37936
rect 23204 37859 23256 37868
rect 23204 37825 23213 37859
rect 23213 37825 23247 37859
rect 23247 37825 23256 37859
rect 23204 37816 23256 37825
rect 22836 37748 22888 37800
rect 16396 37680 16448 37689
rect 17408 37680 17460 37732
rect 19800 37680 19852 37732
rect 22008 37680 22060 37732
rect 22100 37680 22152 37732
rect 24492 37748 24544 37800
rect 14372 37612 14424 37664
rect 15200 37612 15252 37664
rect 16304 37612 16356 37664
rect 18328 37612 18380 37664
rect 18604 37655 18656 37664
rect 18604 37621 18613 37655
rect 18613 37621 18647 37655
rect 18647 37621 18656 37655
rect 18604 37612 18656 37621
rect 19294 37612 19346 37664
rect 20076 37612 20128 37664
rect 23572 37612 23624 37664
rect 24032 37612 24084 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 8576 37451 8628 37460
rect 8576 37417 8585 37451
rect 8585 37417 8619 37451
rect 8619 37417 8628 37451
rect 8576 37408 8628 37417
rect 10416 37451 10468 37460
rect 10416 37417 10425 37451
rect 10425 37417 10459 37451
rect 10459 37417 10468 37451
rect 10416 37408 10468 37417
rect 11704 37408 11756 37460
rect 12256 37408 12308 37460
rect 12440 37383 12492 37392
rect 12440 37349 12449 37383
rect 12449 37349 12483 37383
rect 12483 37349 12492 37383
rect 12440 37340 12492 37349
rect 12808 37340 12860 37392
rect 8760 37272 8812 37324
rect 10968 37315 11020 37324
rect 10968 37281 10977 37315
rect 10977 37281 11011 37315
rect 11011 37281 11020 37315
rect 10968 37272 11020 37281
rect 6552 37204 6604 37256
rect 7748 37136 7800 37188
rect 10048 37204 10100 37256
rect 10416 37136 10468 37188
rect 11888 37204 11940 37256
rect 12992 37340 13044 37392
rect 14464 37340 14516 37392
rect 14096 37272 14148 37324
rect 14188 37272 14240 37324
rect 18696 37408 18748 37460
rect 21824 37408 21876 37460
rect 25228 37408 25280 37460
rect 15752 37340 15804 37392
rect 15384 37272 15436 37324
rect 16212 37272 16264 37324
rect 17040 37340 17092 37392
rect 22468 37340 22520 37392
rect 24124 37340 24176 37392
rect 17868 37315 17920 37324
rect 17868 37281 17877 37315
rect 17877 37281 17911 37315
rect 17911 37281 17920 37315
rect 17868 37272 17920 37281
rect 18512 37272 18564 37324
rect 18696 37272 18748 37324
rect 13544 37204 13596 37256
rect 19248 37272 19300 37324
rect 23664 37272 23716 37324
rect 24032 37315 24084 37324
rect 24032 37281 24041 37315
rect 24041 37281 24075 37315
rect 24075 37281 24084 37315
rect 24032 37272 24084 37281
rect 24400 37272 24452 37324
rect 20720 37204 20772 37256
rect 22100 37204 22152 37256
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 12716 37068 12768 37120
rect 13912 37068 13964 37120
rect 14096 37068 14148 37120
rect 15108 37068 15160 37120
rect 15200 37068 15252 37120
rect 15568 37068 15620 37120
rect 17592 37136 17644 37188
rect 18512 37111 18564 37120
rect 18512 37077 18521 37111
rect 18521 37077 18555 37111
rect 18555 37077 18564 37111
rect 18512 37068 18564 37077
rect 19432 37179 19484 37188
rect 19432 37145 19441 37179
rect 19441 37145 19475 37179
rect 19475 37145 19484 37179
rect 19432 37136 19484 37145
rect 19800 37136 19852 37188
rect 20812 37136 20864 37188
rect 20996 37136 21048 37188
rect 20076 37068 20128 37120
rect 20720 37111 20772 37120
rect 20720 37077 20729 37111
rect 20729 37077 20763 37111
rect 20763 37077 20772 37111
rect 20720 37068 20772 37077
rect 21088 37068 21140 37120
rect 24768 37111 24820 37120
rect 24768 37077 24777 37111
rect 24777 37077 24811 37111
rect 24811 37077 24820 37111
rect 24768 37068 24820 37077
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 5540 36864 5592 36916
rect 6552 36864 6604 36916
rect 7472 36907 7524 36916
rect 7472 36873 7481 36907
rect 7481 36873 7515 36907
rect 7515 36873 7524 36907
rect 7472 36864 7524 36873
rect 8484 36864 8536 36916
rect 9036 36907 9088 36916
rect 9036 36873 9045 36907
rect 9045 36873 9079 36907
rect 9079 36873 9088 36907
rect 9036 36864 9088 36873
rect 10784 36864 10836 36916
rect 12256 36864 12308 36916
rect 13728 36864 13780 36916
rect 14464 36864 14516 36916
rect 15384 36864 15436 36916
rect 15844 36864 15896 36916
rect 16948 36864 17000 36916
rect 6092 36796 6144 36848
rect 10416 36796 10468 36848
rect 9128 36728 9180 36780
rect 9312 36728 9364 36780
rect 11060 36728 11112 36780
rect 12716 36796 12768 36848
rect 13544 36796 13596 36848
rect 18512 36864 18564 36916
rect 19892 36864 19944 36916
rect 20536 36864 20588 36916
rect 22836 36864 22888 36916
rect 18788 36796 18840 36848
rect 23296 36864 23348 36916
rect 23848 36864 23900 36916
rect 24768 36796 24820 36848
rect 5448 36660 5500 36712
rect 5816 36660 5868 36712
rect 6000 36660 6052 36712
rect 9588 36703 9640 36712
rect 9588 36669 9597 36703
rect 9597 36669 9631 36703
rect 9631 36669 9640 36703
rect 9588 36660 9640 36669
rect 10968 36703 11020 36712
rect 10968 36669 10977 36703
rect 10977 36669 11011 36703
rect 11011 36669 11020 36703
rect 10968 36660 11020 36669
rect 7840 36592 7892 36644
rect 9496 36592 9548 36644
rect 12256 36592 12308 36644
rect 12808 36728 12860 36780
rect 14096 36728 14148 36780
rect 14832 36728 14884 36780
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 19340 36728 19392 36780
rect 22100 36728 22152 36780
rect 22836 36771 22888 36780
rect 22836 36737 22845 36771
rect 22845 36737 22879 36771
rect 22879 36737 22888 36771
rect 22836 36728 22888 36737
rect 24400 36728 24452 36780
rect 25320 36771 25372 36780
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 12716 36703 12768 36712
rect 12716 36669 12725 36703
rect 12725 36669 12759 36703
rect 12759 36669 12768 36703
rect 12716 36660 12768 36669
rect 14004 36703 14056 36712
rect 14004 36669 14013 36703
rect 14013 36669 14047 36703
rect 14047 36669 14056 36703
rect 14004 36660 14056 36669
rect 15108 36703 15160 36712
rect 15108 36669 15117 36703
rect 15117 36669 15151 36703
rect 15151 36669 15160 36703
rect 15108 36660 15160 36669
rect 15844 36703 15896 36712
rect 15844 36669 15853 36703
rect 15853 36669 15887 36703
rect 15887 36669 15896 36703
rect 15844 36660 15896 36669
rect 17316 36660 17368 36712
rect 18788 36660 18840 36712
rect 19248 36660 19300 36712
rect 22376 36660 22428 36712
rect 25136 36660 25188 36712
rect 16028 36592 16080 36644
rect 19432 36592 19484 36644
rect 6092 36567 6144 36576
rect 6092 36533 6101 36567
rect 6101 36533 6135 36567
rect 6135 36533 6144 36567
rect 6092 36524 6144 36533
rect 8760 36567 8812 36576
rect 8760 36533 8769 36567
rect 8769 36533 8803 36567
rect 8803 36533 8812 36567
rect 8760 36524 8812 36533
rect 9404 36524 9456 36576
rect 14464 36524 14516 36576
rect 14556 36567 14608 36576
rect 14556 36533 14565 36567
rect 14565 36533 14599 36567
rect 14599 36533 14608 36567
rect 14556 36524 14608 36533
rect 17224 36524 17276 36576
rect 20076 36524 20128 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 7656 36363 7708 36372
rect 7656 36329 7665 36363
rect 7665 36329 7699 36363
rect 7699 36329 7708 36363
rect 7656 36320 7708 36329
rect 8944 36320 8996 36372
rect 9772 36320 9824 36372
rect 13360 36320 13412 36372
rect 15476 36320 15528 36372
rect 19524 36320 19576 36372
rect 21732 36320 21784 36372
rect 13084 36252 13136 36304
rect 18972 36252 19024 36304
rect 24400 36252 24452 36304
rect 7564 36184 7616 36236
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 7840 36116 7892 36168
rect 12440 36227 12492 36236
rect 12440 36193 12449 36227
rect 12449 36193 12483 36227
rect 12483 36193 12492 36227
rect 12440 36184 12492 36193
rect 13360 36227 13412 36236
rect 13360 36193 13369 36227
rect 13369 36193 13403 36227
rect 13403 36193 13412 36227
rect 13360 36184 13412 36193
rect 13544 36184 13596 36236
rect 11796 36116 11848 36168
rect 12072 36116 12124 36168
rect 14004 36116 14056 36168
rect 10324 36048 10376 36100
rect 10692 36048 10744 36100
rect 12256 36048 12308 36100
rect 4160 35980 4212 36032
rect 7472 35980 7524 36032
rect 11244 35980 11296 36032
rect 13084 36023 13136 36032
rect 13084 35989 13093 36023
rect 13093 35989 13127 36023
rect 13127 35989 13136 36023
rect 13084 35980 13136 35989
rect 13636 35980 13688 36032
rect 14648 36023 14700 36032
rect 14648 35989 14657 36023
rect 14657 35989 14691 36023
rect 14691 35989 14700 36023
rect 14648 35980 14700 35989
rect 15016 36184 15068 36236
rect 15752 36227 15804 36236
rect 15752 36193 15761 36227
rect 15761 36193 15795 36227
rect 15795 36193 15804 36227
rect 15752 36184 15804 36193
rect 16488 36184 16540 36236
rect 16948 36184 17000 36236
rect 21272 36227 21324 36236
rect 21272 36193 21281 36227
rect 21281 36193 21315 36227
rect 21315 36193 21324 36227
rect 21272 36184 21324 36193
rect 21640 36184 21692 36236
rect 23756 36227 23808 36236
rect 23756 36193 23765 36227
rect 23765 36193 23799 36227
rect 23799 36193 23808 36227
rect 23756 36184 23808 36193
rect 24492 36184 24544 36236
rect 21916 36116 21968 36168
rect 24584 36116 24636 36168
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 20536 35980 20588 36032
rect 20812 36023 20864 36032
rect 20812 35989 20821 36023
rect 20821 35989 20855 36023
rect 20855 35989 20864 36023
rect 20812 35980 20864 35989
rect 21456 35980 21508 36032
rect 22376 35980 22428 36032
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 5540 35776 5592 35828
rect 6000 35819 6052 35828
rect 6000 35785 6009 35819
rect 6009 35785 6043 35819
rect 6043 35785 6052 35819
rect 6000 35776 6052 35785
rect 6092 35640 6144 35692
rect 5816 35572 5868 35624
rect 7656 35436 7708 35488
rect 9588 35572 9640 35624
rect 8852 35436 8904 35488
rect 9588 35436 9640 35488
rect 13452 35776 13504 35828
rect 14648 35776 14700 35828
rect 15016 35776 15068 35828
rect 17132 35776 17184 35828
rect 17684 35776 17736 35828
rect 11888 35708 11940 35760
rect 9772 35436 9824 35488
rect 13360 35640 13412 35692
rect 17776 35708 17828 35760
rect 19248 35776 19300 35828
rect 21548 35776 21600 35828
rect 23296 35776 23348 35828
rect 10968 35572 11020 35624
rect 13820 35572 13872 35624
rect 12532 35436 12584 35488
rect 13544 35504 13596 35556
rect 13728 35479 13780 35488
rect 13728 35445 13737 35479
rect 13737 35445 13771 35479
rect 13771 35445 13780 35479
rect 13728 35436 13780 35445
rect 15936 35436 15988 35488
rect 19248 35640 19300 35692
rect 20260 35615 20312 35624
rect 20260 35581 20269 35615
rect 20269 35581 20303 35615
rect 20303 35581 20312 35615
rect 20260 35572 20312 35581
rect 22192 35640 22244 35692
rect 22836 35640 22888 35692
rect 24492 35640 24544 35692
rect 22468 35615 22520 35624
rect 22468 35581 22477 35615
rect 22477 35581 22511 35615
rect 22511 35581 22520 35615
rect 22468 35572 22520 35581
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 18328 35436 18380 35488
rect 19708 35436 19760 35488
rect 19800 35479 19852 35488
rect 19800 35445 19809 35479
rect 19809 35445 19843 35479
rect 19843 35445 19852 35479
rect 19800 35436 19852 35445
rect 20904 35479 20956 35488
rect 20904 35445 20913 35479
rect 20913 35445 20947 35479
rect 20947 35445 20956 35479
rect 20904 35436 20956 35445
rect 23940 35436 23992 35488
rect 24492 35436 24544 35488
rect 24768 35436 24820 35488
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 7380 35232 7432 35284
rect 11060 35232 11112 35284
rect 16120 35232 16172 35284
rect 19064 35232 19116 35284
rect 21180 35232 21232 35284
rect 7840 35207 7892 35216
rect 7840 35173 7849 35207
rect 7849 35173 7883 35207
rect 7883 35173 7892 35207
rect 7840 35164 7892 35173
rect 8576 35164 8628 35216
rect 5540 35096 5592 35148
rect 6092 35139 6144 35148
rect 6092 35105 6101 35139
rect 6101 35105 6135 35139
rect 6135 35105 6144 35139
rect 6092 35096 6144 35105
rect 9772 35096 9824 35148
rect 16672 35164 16724 35216
rect 19156 35164 19208 35216
rect 11060 35096 11112 35148
rect 15752 35096 15804 35148
rect 16120 35096 16172 35148
rect 19708 35096 19760 35148
rect 20260 35096 20312 35148
rect 20720 35096 20772 35148
rect 20904 35096 20956 35148
rect 21640 35096 21692 35148
rect 8300 35028 8352 35080
rect 12716 35028 12768 35080
rect 14556 35028 14608 35080
rect 22192 35028 22244 35080
rect 7656 34960 7708 35012
rect 8668 34960 8720 35012
rect 14280 34960 14332 35012
rect 7840 34892 7892 34944
rect 13360 34935 13412 34944
rect 13360 34901 13369 34935
rect 13369 34901 13403 34935
rect 13403 34901 13412 34935
rect 13360 34892 13412 34901
rect 16120 34960 16172 35012
rect 19156 34960 19208 35012
rect 19708 35003 19760 35012
rect 19708 34969 19717 35003
rect 19717 34969 19751 35003
rect 19751 34969 19760 35003
rect 19708 34960 19760 34969
rect 19984 34960 20036 35012
rect 22560 35003 22612 35012
rect 22560 34969 22569 35003
rect 22569 34969 22603 35003
rect 22603 34969 22612 35003
rect 22560 34960 22612 34969
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 23388 34892 23440 34944
rect 24492 34935 24544 34944
rect 24492 34901 24501 34935
rect 24501 34901 24535 34935
rect 24535 34901 24544 34935
rect 24492 34892 24544 34901
rect 24768 34892 24820 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 7104 34688 7156 34740
rect 8300 34731 8352 34740
rect 8300 34697 8309 34731
rect 8309 34697 8343 34731
rect 8343 34697 8352 34731
rect 8300 34688 8352 34697
rect 9496 34688 9548 34740
rect 13728 34731 13780 34740
rect 6000 34620 6052 34672
rect 9588 34620 9640 34672
rect 11888 34620 11940 34672
rect 13728 34697 13737 34731
rect 13737 34697 13771 34731
rect 13771 34697 13780 34731
rect 13728 34688 13780 34697
rect 14188 34688 14240 34740
rect 19800 34688 19852 34740
rect 20996 34688 21048 34740
rect 21180 34731 21232 34740
rect 21180 34697 21189 34731
rect 21189 34697 21223 34731
rect 21223 34697 21232 34731
rect 21180 34688 21232 34697
rect 22376 34731 22428 34740
rect 22376 34697 22385 34731
rect 22385 34697 22419 34731
rect 22419 34697 22428 34731
rect 22376 34688 22428 34697
rect 22468 34688 22520 34740
rect 24676 34688 24728 34740
rect 14372 34620 14424 34672
rect 15200 34620 15252 34672
rect 15752 34620 15804 34672
rect 18420 34620 18472 34672
rect 18788 34620 18840 34672
rect 19984 34620 20036 34672
rect 6092 34552 6144 34604
rect 7932 34552 7984 34604
rect 8852 34595 8904 34604
rect 8852 34561 8861 34595
rect 8861 34561 8895 34595
rect 8895 34561 8904 34595
rect 8852 34552 8904 34561
rect 19616 34552 19668 34604
rect 22284 34552 22336 34604
rect 22652 34552 22704 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 7288 34484 7340 34536
rect 8760 34484 8812 34536
rect 9588 34484 9640 34536
rect 9864 34484 9916 34536
rect 10416 34484 10468 34536
rect 10968 34484 11020 34536
rect 13820 34484 13872 34536
rect 14832 34484 14884 34536
rect 4804 34416 4856 34468
rect 5632 34416 5684 34468
rect 10140 34348 10192 34400
rect 11060 34416 11112 34468
rect 15844 34416 15896 34468
rect 19892 34416 19944 34468
rect 22652 34416 22704 34468
rect 23572 34484 23624 34536
rect 23664 34527 23716 34536
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 23848 34416 23900 34468
rect 10968 34391 11020 34400
rect 10968 34357 10977 34391
rect 10977 34357 11011 34391
rect 11011 34357 11020 34391
rect 10968 34348 11020 34357
rect 11796 34348 11848 34400
rect 12072 34348 12124 34400
rect 20720 34391 20772 34400
rect 20720 34357 20729 34391
rect 20729 34357 20763 34391
rect 20763 34357 20772 34391
rect 20720 34348 20772 34357
rect 22008 34391 22060 34400
rect 22008 34357 22017 34391
rect 22017 34357 22051 34391
rect 22051 34357 22060 34391
rect 22008 34348 22060 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 7380 34144 7432 34196
rect 9128 34187 9180 34196
rect 9128 34153 9137 34187
rect 9137 34153 9171 34187
rect 9171 34153 9180 34187
rect 9128 34144 9180 34153
rect 10692 34144 10744 34196
rect 7196 34076 7248 34128
rect 10232 34076 10284 34128
rect 19708 34144 19760 34196
rect 20168 34144 20220 34196
rect 20904 34144 20956 34196
rect 22284 34144 22336 34196
rect 25320 34187 25372 34196
rect 25320 34153 25329 34187
rect 25329 34153 25363 34187
rect 25363 34153 25372 34187
rect 25320 34144 25372 34153
rect 5540 34051 5592 34060
rect 5540 34017 5549 34051
rect 5549 34017 5583 34051
rect 5583 34017 5592 34051
rect 5540 34008 5592 34017
rect 5816 34008 5868 34060
rect 9220 34008 9272 34060
rect 12532 34008 12584 34060
rect 12624 34008 12676 34060
rect 13820 34076 13872 34128
rect 15936 34051 15988 34060
rect 15936 34017 15945 34051
rect 15945 34017 15979 34051
rect 15979 34017 15988 34051
rect 15936 34008 15988 34017
rect 19800 34076 19852 34128
rect 7380 33940 7432 33992
rect 8852 33940 8904 33992
rect 9588 33940 9640 33992
rect 10416 33983 10468 33992
rect 10416 33949 10425 33983
rect 10425 33949 10459 33983
rect 10459 33949 10468 33983
rect 10416 33940 10468 33949
rect 11796 33940 11848 33992
rect 12808 33940 12860 33992
rect 13728 33940 13780 33992
rect 18420 34008 18472 34060
rect 21640 34051 21692 34060
rect 21640 34017 21649 34051
rect 21649 34017 21683 34051
rect 21683 34017 21692 34051
rect 21640 34008 21692 34017
rect 22744 34051 22796 34060
rect 22744 34017 22753 34051
rect 22753 34017 22787 34051
rect 22787 34017 22796 34051
rect 22744 34008 22796 34017
rect 23388 34008 23440 34060
rect 19616 33940 19668 33992
rect 20076 33940 20128 33992
rect 20628 33940 20680 33992
rect 24216 33940 24268 33992
rect 24308 33940 24360 33992
rect 7656 33872 7708 33924
rect 9864 33872 9916 33924
rect 10968 33872 11020 33924
rect 15568 33872 15620 33924
rect 7196 33804 7248 33856
rect 7932 33804 7984 33856
rect 11980 33804 12032 33856
rect 12808 33804 12860 33856
rect 13544 33804 13596 33856
rect 15016 33804 15068 33856
rect 16120 33804 16172 33856
rect 19064 33804 19116 33856
rect 19984 33872 20036 33924
rect 24492 33872 24544 33924
rect 20168 33804 20220 33856
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 21456 33847 21508 33856
rect 21456 33813 21465 33847
rect 21465 33813 21499 33847
rect 21499 33813 21508 33847
rect 21456 33804 21508 33813
rect 22284 33847 22336 33856
rect 22284 33813 22293 33847
rect 22293 33813 22327 33847
rect 22327 33813 22336 33847
rect 22284 33804 22336 33813
rect 22468 33804 22520 33856
rect 24308 33804 24360 33856
rect 24584 33847 24636 33856
rect 24584 33813 24593 33847
rect 24593 33813 24627 33847
rect 24627 33813 24636 33847
rect 24584 33804 24636 33813
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 10324 33600 10376 33652
rect 10784 33600 10836 33652
rect 11244 33600 11296 33652
rect 1308 33464 1360 33516
rect 11612 33464 11664 33516
rect 13268 33507 13320 33516
rect 13268 33473 13277 33507
rect 13277 33473 13311 33507
rect 13311 33473 13320 33507
rect 13268 33464 13320 33473
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 9772 33439 9824 33448
rect 9772 33405 9781 33439
rect 9781 33405 9815 33439
rect 9815 33405 9824 33439
rect 9772 33396 9824 33405
rect 13820 33600 13872 33652
rect 14556 33600 14608 33652
rect 15936 33600 15988 33652
rect 19156 33600 19208 33652
rect 19984 33600 20036 33652
rect 14372 33532 14424 33584
rect 14648 33532 14700 33584
rect 18328 33532 18380 33584
rect 20168 33532 20220 33584
rect 21180 33600 21232 33652
rect 21456 33600 21508 33652
rect 25228 33643 25280 33652
rect 25228 33609 25237 33643
rect 25237 33609 25271 33643
rect 25271 33609 25280 33643
rect 25228 33600 25280 33609
rect 23664 33532 23716 33584
rect 24308 33532 24360 33584
rect 20628 33507 20680 33516
rect 20628 33473 20637 33507
rect 20637 33473 20671 33507
rect 20671 33473 20680 33507
rect 20628 33464 20680 33473
rect 8300 33328 8352 33380
rect 13452 33439 13504 33448
rect 13452 33405 13461 33439
rect 13461 33405 13495 33439
rect 13495 33405 13504 33439
rect 13452 33396 13504 33405
rect 16672 33396 16724 33448
rect 20996 33396 21048 33448
rect 22192 33464 22244 33516
rect 23296 33396 23348 33448
rect 23756 33439 23808 33448
rect 23756 33405 23765 33439
rect 23765 33405 23799 33439
rect 23799 33405 23808 33439
rect 23756 33396 23808 33405
rect 21640 33328 21692 33380
rect 3516 33260 3568 33312
rect 7196 33303 7248 33312
rect 7196 33269 7205 33303
rect 7205 33269 7239 33303
rect 7239 33269 7248 33303
rect 7196 33260 7248 33269
rect 12440 33260 12492 33312
rect 13268 33260 13320 33312
rect 13452 33260 13504 33312
rect 15844 33303 15896 33312
rect 15844 33269 15853 33303
rect 15853 33269 15887 33303
rect 15887 33269 15896 33303
rect 15844 33260 15896 33269
rect 16120 33303 16172 33312
rect 16120 33269 16129 33303
rect 16129 33269 16163 33303
rect 16163 33269 16172 33303
rect 16120 33260 16172 33269
rect 16396 33260 16448 33312
rect 16856 33260 16908 33312
rect 20352 33260 20404 33312
rect 22744 33260 22796 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 7472 33099 7524 33108
rect 7472 33065 7481 33099
rect 7481 33065 7515 33099
rect 7515 33065 7524 33099
rect 7472 33056 7524 33065
rect 9312 33056 9364 33108
rect 10232 33056 10284 33108
rect 7564 32988 7616 33040
rect 5540 32920 5592 32972
rect 7196 32920 7248 32972
rect 9128 32988 9180 33040
rect 8300 32920 8352 32972
rect 10140 32920 10192 32972
rect 9772 32895 9824 32904
rect 9772 32861 9781 32895
rect 9781 32861 9815 32895
rect 9815 32861 9824 32895
rect 9772 32852 9824 32861
rect 7748 32784 7800 32836
rect 10876 33056 10928 33108
rect 12164 33099 12216 33108
rect 12164 33065 12173 33099
rect 12173 33065 12207 33099
rect 12207 33065 12216 33099
rect 12164 33056 12216 33065
rect 11520 32920 11572 32972
rect 14372 33056 14424 33108
rect 15016 33056 15068 33108
rect 20628 33056 20680 33108
rect 20904 33056 20956 33108
rect 12624 32988 12676 33040
rect 13912 32988 13964 33040
rect 17040 32988 17092 33040
rect 17132 33031 17184 33040
rect 17132 32997 17141 33031
rect 17141 32997 17175 33031
rect 17175 32997 17184 33031
rect 17132 32988 17184 32997
rect 14464 32920 14516 32972
rect 14832 32963 14884 32972
rect 14832 32929 14841 32963
rect 14841 32929 14875 32963
rect 14875 32929 14884 32963
rect 14832 32920 14884 32929
rect 16396 32920 16448 32972
rect 16488 32920 16540 32972
rect 16856 32920 16908 32972
rect 20076 32988 20128 33040
rect 15844 32852 15896 32904
rect 16764 32852 16816 32904
rect 17500 32852 17552 32904
rect 19248 32852 19300 32904
rect 11888 32784 11940 32836
rect 14372 32784 14424 32836
rect 22560 32988 22612 33040
rect 21640 32963 21692 32972
rect 21640 32929 21649 32963
rect 21649 32929 21683 32963
rect 21683 32929 21692 32963
rect 21640 32920 21692 32929
rect 24032 32988 24084 33040
rect 20996 32852 21048 32904
rect 21180 32852 21232 32904
rect 21456 32852 21508 32904
rect 22376 32895 22428 32904
rect 22376 32861 22385 32895
rect 22385 32861 22419 32895
rect 22419 32861 22428 32895
rect 22376 32852 22428 32861
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 7840 32759 7892 32768
rect 7840 32725 7849 32759
rect 7849 32725 7883 32759
rect 7883 32725 7892 32759
rect 7840 32716 7892 32725
rect 9496 32716 9548 32768
rect 14648 32759 14700 32768
rect 14648 32725 14657 32759
rect 14657 32725 14691 32759
rect 14691 32725 14700 32759
rect 14648 32716 14700 32725
rect 16120 32759 16172 32768
rect 16120 32725 16129 32759
rect 16129 32725 16163 32759
rect 16163 32725 16172 32759
rect 16120 32716 16172 32725
rect 16396 32716 16448 32768
rect 18604 32716 18656 32768
rect 22468 32784 22520 32836
rect 20076 32716 20128 32768
rect 20904 32716 20956 32768
rect 21272 32716 21324 32768
rect 21640 32716 21692 32768
rect 22376 32716 22428 32768
rect 22560 32716 22612 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 4620 32555 4672 32564
rect 4620 32521 4629 32555
rect 4629 32521 4663 32555
rect 4663 32521 4672 32555
rect 4620 32512 4672 32521
rect 4988 32555 5040 32564
rect 4988 32521 4997 32555
rect 4997 32521 5031 32555
rect 5031 32521 5040 32555
rect 4988 32512 5040 32521
rect 5356 32555 5408 32564
rect 5356 32521 5365 32555
rect 5365 32521 5399 32555
rect 5399 32521 5408 32555
rect 5356 32512 5408 32521
rect 7840 32512 7892 32564
rect 14648 32512 14700 32564
rect 14740 32512 14792 32564
rect 4896 32444 4948 32496
rect 5540 32444 5592 32496
rect 6184 32444 6236 32496
rect 9128 32444 9180 32496
rect 10232 32444 10284 32496
rect 10968 32444 11020 32496
rect 12532 32444 12584 32496
rect 5448 32308 5500 32360
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 12256 32308 12308 32360
rect 14832 32487 14884 32496
rect 14832 32453 14841 32487
rect 14841 32453 14875 32487
rect 14875 32453 14884 32487
rect 14832 32444 14884 32453
rect 16120 32512 16172 32564
rect 17224 32487 17276 32496
rect 17224 32453 17233 32487
rect 17233 32453 17267 32487
rect 17267 32453 17276 32487
rect 17224 32444 17276 32453
rect 14556 32419 14608 32428
rect 14556 32385 14565 32419
rect 14565 32385 14599 32419
rect 14599 32385 14608 32419
rect 14556 32376 14608 32385
rect 18880 32376 18932 32428
rect 19248 32376 19300 32428
rect 20996 32512 21048 32564
rect 21824 32555 21876 32564
rect 21824 32521 21833 32555
rect 21833 32521 21867 32555
rect 21867 32521 21876 32555
rect 21824 32512 21876 32521
rect 20904 32376 20956 32428
rect 22100 32376 22152 32428
rect 22744 32376 22796 32428
rect 25412 32376 25464 32428
rect 7564 32240 7616 32292
rect 12072 32240 12124 32292
rect 16672 32308 16724 32360
rect 17776 32308 17828 32360
rect 18604 32351 18656 32360
rect 18604 32317 18613 32351
rect 18613 32317 18647 32351
rect 18647 32317 18656 32351
rect 18604 32308 18656 32317
rect 9220 32172 9272 32224
rect 10232 32172 10284 32224
rect 12532 32172 12584 32224
rect 13544 32240 13596 32292
rect 15936 32240 15988 32292
rect 12716 32172 12768 32224
rect 14464 32172 14516 32224
rect 14556 32172 14608 32224
rect 15200 32172 15252 32224
rect 16948 32172 17000 32224
rect 17132 32240 17184 32292
rect 20628 32308 20680 32360
rect 21364 32351 21416 32360
rect 21364 32317 21373 32351
rect 21373 32317 21407 32351
rect 21407 32317 21416 32351
rect 21364 32308 21416 32317
rect 17960 32172 18012 32224
rect 18696 32172 18748 32224
rect 20076 32215 20128 32224
rect 20076 32181 20085 32215
rect 20085 32181 20119 32215
rect 20119 32181 20128 32215
rect 20076 32172 20128 32181
rect 21364 32172 21416 32224
rect 21824 32172 21876 32224
rect 22100 32172 22152 32224
rect 22744 32172 22796 32224
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 8300 31968 8352 32020
rect 6184 31875 6236 31884
rect 6184 31841 6193 31875
rect 6193 31841 6227 31875
rect 6227 31841 6236 31875
rect 6184 31832 6236 31841
rect 7104 31832 7156 31884
rect 9128 31968 9180 32020
rect 10140 31968 10192 32020
rect 11612 31968 11664 32020
rect 17960 31968 18012 32020
rect 18420 31968 18472 32020
rect 9220 31900 9272 31952
rect 11244 31900 11296 31952
rect 14096 31900 14148 31952
rect 14280 31943 14332 31952
rect 14280 31909 14289 31943
rect 14289 31909 14323 31943
rect 14323 31909 14332 31943
rect 14280 31900 14332 31909
rect 14648 31900 14700 31952
rect 15108 31900 15160 31952
rect 15936 31900 15988 31952
rect 16120 31900 16172 31952
rect 19432 31943 19484 31952
rect 19432 31909 19441 31943
rect 19441 31909 19475 31943
rect 19475 31909 19484 31943
rect 19432 31900 19484 31909
rect 8300 31807 8352 31816
rect 8300 31773 8309 31807
rect 8309 31773 8343 31807
rect 8343 31773 8352 31807
rect 8300 31764 8352 31773
rect 11428 31832 11480 31884
rect 13820 31832 13872 31884
rect 14648 31764 14700 31816
rect 14740 31807 14792 31816
rect 14740 31773 14749 31807
rect 14749 31773 14783 31807
rect 14783 31773 14792 31807
rect 14740 31764 14792 31773
rect 18236 31875 18288 31884
rect 18236 31841 18245 31875
rect 18245 31841 18279 31875
rect 18279 31841 18288 31875
rect 18236 31832 18288 31841
rect 19156 31832 19208 31884
rect 19984 31875 20036 31884
rect 19984 31841 19993 31875
rect 19993 31841 20027 31875
rect 20027 31841 20036 31875
rect 19984 31832 20036 31841
rect 20260 31900 20312 31952
rect 20904 31968 20956 32020
rect 23296 31968 23348 32020
rect 24216 31968 24268 32020
rect 21640 31900 21692 31952
rect 23388 31900 23440 31952
rect 21364 31832 21416 31884
rect 23480 31832 23532 31884
rect 9588 31696 9640 31748
rect 7380 31628 7432 31680
rect 8300 31628 8352 31680
rect 9128 31671 9180 31680
rect 9128 31637 9137 31671
rect 9137 31637 9171 31671
rect 9171 31637 9180 31671
rect 9128 31628 9180 31637
rect 10140 31696 10192 31748
rect 14464 31696 14516 31748
rect 17132 31764 17184 31816
rect 18052 31764 18104 31816
rect 18880 31764 18932 31816
rect 20812 31764 20864 31816
rect 21640 31764 21692 31816
rect 21916 31764 21968 31816
rect 24308 31764 24360 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 19800 31739 19852 31748
rect 19800 31705 19809 31739
rect 19809 31705 19843 31739
rect 19843 31705 19852 31739
rect 19800 31696 19852 31705
rect 21180 31696 21232 31748
rect 21272 31696 21324 31748
rect 13820 31628 13872 31680
rect 15016 31628 15068 31680
rect 17684 31628 17736 31680
rect 20076 31628 20128 31680
rect 21456 31628 21508 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 7656 31424 7708 31476
rect 8668 31467 8720 31476
rect 8668 31433 8677 31467
rect 8677 31433 8711 31467
rect 8711 31433 8720 31467
rect 8668 31424 8720 31433
rect 9864 31424 9916 31476
rect 13360 31424 13412 31476
rect 18604 31424 18656 31476
rect 18972 31424 19024 31476
rect 1952 31288 2004 31340
rect 7840 31331 7892 31340
rect 7840 31297 7849 31331
rect 7849 31297 7883 31331
rect 7883 31297 7892 31331
rect 7840 31288 7892 31297
rect 1308 31220 1360 31272
rect 5632 31220 5684 31272
rect 8760 31288 8812 31340
rect 11244 31356 11296 31408
rect 15108 31356 15160 31408
rect 18420 31356 18472 31408
rect 18788 31356 18840 31408
rect 8116 31263 8168 31272
rect 8116 31229 8125 31263
rect 8125 31229 8159 31263
rect 8159 31229 8168 31263
rect 8116 31220 8168 31229
rect 8484 31220 8536 31272
rect 9588 31220 9640 31272
rect 5908 31152 5960 31204
rect 13268 31220 13320 31272
rect 14924 31220 14976 31272
rect 18328 31288 18380 31340
rect 18972 31288 19024 31340
rect 17868 31220 17920 31272
rect 18788 31263 18840 31272
rect 18788 31229 18797 31263
rect 18797 31229 18831 31263
rect 18831 31229 18840 31263
rect 18788 31220 18840 31229
rect 18880 31263 18932 31272
rect 18880 31229 18889 31263
rect 18889 31229 18923 31263
rect 18923 31229 18932 31263
rect 18880 31220 18932 31229
rect 15476 31152 15528 31204
rect 19340 31220 19392 31272
rect 20076 31424 20128 31476
rect 21640 31424 21692 31476
rect 22652 31424 22704 31476
rect 23940 31424 23992 31476
rect 21824 31288 21876 31340
rect 24308 31356 24360 31408
rect 24400 31288 24452 31340
rect 25320 31331 25372 31340
rect 25320 31297 25329 31331
rect 25329 31297 25363 31331
rect 25363 31297 25372 31331
rect 25320 31288 25372 31297
rect 20628 31220 20680 31272
rect 22192 31263 22244 31272
rect 22192 31229 22201 31263
rect 22201 31229 22235 31263
rect 22235 31229 22244 31263
rect 22192 31220 22244 31229
rect 14464 31084 14516 31136
rect 14648 31127 14700 31136
rect 14648 31093 14657 31127
rect 14657 31093 14691 31127
rect 14691 31093 14700 31127
rect 14648 31084 14700 31093
rect 15292 31084 15344 31136
rect 17132 31127 17184 31136
rect 17132 31093 17141 31127
rect 17141 31093 17175 31127
rect 17175 31093 17184 31127
rect 17132 31084 17184 31093
rect 21916 31152 21968 31204
rect 23572 31084 23624 31136
rect 24492 31084 24544 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 8116 30880 8168 30932
rect 11980 30880 12032 30932
rect 1676 30744 1728 30796
rect 7840 30744 7892 30796
rect 9588 30787 9640 30796
rect 9588 30753 9597 30787
rect 9597 30753 9631 30787
rect 9631 30753 9640 30787
rect 9588 30744 9640 30753
rect 10600 30744 10652 30796
rect 11428 30676 11480 30728
rect 18512 30880 18564 30932
rect 20444 30923 20496 30932
rect 15200 30744 15252 30796
rect 16488 30787 16540 30796
rect 16488 30753 16497 30787
rect 16497 30753 16531 30787
rect 16531 30753 16540 30787
rect 16488 30744 16540 30753
rect 18880 30744 18932 30796
rect 20444 30889 20453 30923
rect 20453 30889 20487 30923
rect 20487 30889 20496 30923
rect 20444 30880 20496 30889
rect 20536 30880 20588 30932
rect 17500 30676 17552 30728
rect 19984 30787 20036 30796
rect 19984 30753 19993 30787
rect 19993 30753 20027 30787
rect 20027 30753 20036 30787
rect 19984 30744 20036 30753
rect 20444 30744 20496 30796
rect 22836 30880 22888 30932
rect 25320 30880 25372 30932
rect 19432 30676 19484 30728
rect 19708 30676 19760 30728
rect 22284 30676 22336 30728
rect 25504 30676 25556 30728
rect 3792 30608 3844 30660
rect 5908 30608 5960 30660
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 10232 30540 10284 30592
rect 16580 30608 16632 30660
rect 11336 30583 11388 30592
rect 11336 30549 11345 30583
rect 11345 30549 11379 30583
rect 11379 30549 11388 30583
rect 11336 30540 11388 30549
rect 15108 30540 15160 30592
rect 18788 30608 18840 30660
rect 24768 30608 24820 30660
rect 17408 30540 17460 30592
rect 17500 30540 17552 30592
rect 17776 30540 17828 30592
rect 18604 30540 18656 30592
rect 19156 30540 19208 30592
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 21824 30540 21876 30592
rect 22836 30540 22888 30592
rect 24952 30540 25004 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 6368 30268 6420 30320
rect 9588 30268 9640 30320
rect 11796 30268 11848 30320
rect 14280 30268 14332 30320
rect 15200 30268 15252 30320
rect 10508 30132 10560 30184
rect 10692 30132 10744 30184
rect 10600 30064 10652 30116
rect 10416 30039 10468 30048
rect 10416 30005 10425 30039
rect 10425 30005 10459 30039
rect 10459 30005 10468 30039
rect 10416 29996 10468 30005
rect 11888 29996 11940 30048
rect 14372 30200 14424 30252
rect 14464 30243 14516 30252
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 18328 30336 18380 30388
rect 19156 30336 19208 30388
rect 19340 30336 19392 30388
rect 20904 30336 20956 30388
rect 24308 30336 24360 30388
rect 17592 30268 17644 30320
rect 23572 30268 23624 30320
rect 20168 30200 20220 30252
rect 20352 30200 20404 30252
rect 22192 30200 22244 30252
rect 14832 30132 14884 30184
rect 16212 30175 16264 30184
rect 16212 30141 16221 30175
rect 16221 30141 16255 30175
rect 16255 30141 16264 30175
rect 16212 30132 16264 30141
rect 17224 30132 17276 30184
rect 18052 30175 18104 30184
rect 18052 30141 18061 30175
rect 18061 30141 18095 30175
rect 18095 30141 18104 30175
rect 18052 30132 18104 30141
rect 19892 30132 19944 30184
rect 23756 30132 23808 30184
rect 15752 30064 15804 30116
rect 21548 30064 21600 30116
rect 17500 29996 17552 30048
rect 17592 30039 17644 30048
rect 17592 30005 17601 30039
rect 17601 30005 17635 30039
rect 17635 30005 17644 30039
rect 17592 29996 17644 30005
rect 18052 29996 18104 30048
rect 18512 29996 18564 30048
rect 18880 29996 18932 30048
rect 19340 29996 19392 30048
rect 21732 29996 21784 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 4252 29792 4304 29844
rect 7656 29792 7708 29844
rect 7748 29792 7800 29844
rect 9496 29835 9548 29844
rect 9496 29801 9505 29835
rect 9505 29801 9539 29835
rect 9539 29801 9548 29835
rect 9496 29792 9548 29801
rect 12900 29792 12952 29844
rect 11336 29724 11388 29776
rect 1584 29656 1636 29708
rect 7104 29656 7156 29708
rect 9128 29656 9180 29708
rect 7288 29588 7340 29640
rect 7840 29588 7892 29640
rect 14740 29724 14792 29776
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16488 29792 16540 29844
rect 16580 29792 16632 29844
rect 17316 29792 17368 29844
rect 23940 29792 23992 29844
rect 16672 29724 16724 29776
rect 17592 29724 17644 29776
rect 14464 29656 14516 29708
rect 18788 29699 18840 29708
rect 18788 29665 18797 29699
rect 18797 29665 18831 29699
rect 18831 29665 18840 29699
rect 18788 29656 18840 29665
rect 24400 29724 24452 29776
rect 21180 29656 21232 29708
rect 22560 29656 22612 29708
rect 23388 29699 23440 29708
rect 23388 29665 23397 29699
rect 23397 29665 23431 29699
rect 23431 29665 23440 29699
rect 23388 29656 23440 29665
rect 23756 29656 23808 29708
rect 10416 29588 10468 29640
rect 16396 29588 16448 29640
rect 20720 29588 20772 29640
rect 22008 29588 22060 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 3884 29520 3936 29572
rect 6368 29520 6420 29572
rect 7012 29520 7064 29572
rect 9312 29520 9364 29572
rect 9588 29520 9640 29572
rect 11796 29563 11848 29572
rect 11796 29529 11805 29563
rect 11805 29529 11839 29563
rect 11839 29529 11848 29563
rect 11796 29520 11848 29529
rect 12808 29520 12860 29572
rect 16764 29520 16816 29572
rect 17592 29520 17644 29572
rect 20168 29520 20220 29572
rect 7380 29452 7432 29504
rect 7656 29452 7708 29504
rect 9956 29495 10008 29504
rect 9956 29461 9965 29495
rect 9965 29461 9999 29495
rect 9999 29461 10008 29495
rect 9956 29452 10008 29461
rect 10416 29452 10468 29504
rect 10784 29452 10836 29504
rect 11888 29495 11940 29504
rect 11888 29461 11897 29495
rect 11897 29461 11931 29495
rect 11931 29461 11940 29495
rect 11888 29452 11940 29461
rect 14004 29452 14056 29504
rect 14924 29452 14976 29504
rect 16580 29452 16632 29504
rect 17500 29452 17552 29504
rect 18328 29452 18380 29504
rect 20352 29452 20404 29504
rect 20904 29495 20956 29504
rect 20904 29461 20913 29495
rect 20913 29461 20947 29495
rect 20947 29461 20956 29495
rect 20904 29452 20956 29461
rect 21916 29452 21968 29504
rect 22836 29452 22888 29504
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 7656 29248 7708 29300
rect 10232 29180 10284 29232
rect 12900 29291 12952 29300
rect 12900 29257 12909 29291
rect 12909 29257 12943 29291
rect 12943 29257 12952 29291
rect 12900 29248 12952 29257
rect 13544 29248 13596 29300
rect 13728 29248 13780 29300
rect 14188 29291 14240 29300
rect 14188 29257 14197 29291
rect 14197 29257 14231 29291
rect 14231 29257 14240 29291
rect 14188 29248 14240 29257
rect 16120 29248 16172 29300
rect 17224 29291 17276 29300
rect 17224 29257 17233 29291
rect 17233 29257 17267 29291
rect 17267 29257 17276 29291
rect 17224 29248 17276 29257
rect 17500 29248 17552 29300
rect 17592 29248 17644 29300
rect 6552 29044 6604 29096
rect 9404 29044 9456 29096
rect 10876 28976 10928 29028
rect 8668 28908 8720 28960
rect 13728 29112 13780 29164
rect 13452 28976 13504 29028
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 14280 29112 14332 29164
rect 14648 29044 14700 29096
rect 15292 29044 15344 29096
rect 15568 29180 15620 29232
rect 18880 29180 18932 29232
rect 20904 29248 20956 29300
rect 23940 29291 23992 29300
rect 23940 29257 23949 29291
rect 23949 29257 23983 29291
rect 23983 29257 23992 29291
rect 23940 29248 23992 29257
rect 25320 29291 25372 29300
rect 25320 29257 25329 29291
rect 25329 29257 25363 29291
rect 25363 29257 25372 29291
rect 25320 29248 25372 29257
rect 25504 29291 25556 29300
rect 25504 29257 25513 29291
rect 25513 29257 25547 29291
rect 25547 29257 25556 29291
rect 25504 29248 25556 29257
rect 20076 29180 20128 29232
rect 16120 29112 16172 29164
rect 16396 29087 16448 29096
rect 16396 29053 16405 29087
rect 16405 29053 16439 29087
rect 16439 29053 16448 29087
rect 16396 29044 16448 29053
rect 16672 29044 16724 29096
rect 14004 28908 14056 28960
rect 14188 28908 14240 28960
rect 15752 28908 15804 28960
rect 16028 28976 16080 29028
rect 17408 29087 17460 29096
rect 17408 29053 17417 29087
rect 17417 29053 17451 29087
rect 17451 29053 17460 29087
rect 17408 29044 17460 29053
rect 17592 28976 17644 29028
rect 19524 29044 19576 29096
rect 20996 29044 21048 29096
rect 21548 29223 21600 29232
rect 21548 29189 21557 29223
rect 21557 29189 21591 29223
rect 21591 29189 21600 29223
rect 21548 29180 21600 29189
rect 24584 29180 24636 29232
rect 23480 29112 23532 29164
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 23572 29044 23624 29096
rect 18052 29019 18104 29028
rect 18052 28985 18061 29019
rect 18061 28985 18095 29019
rect 18095 28985 18104 29019
rect 18052 28976 18104 28985
rect 18328 28976 18380 29028
rect 18420 28908 18472 28960
rect 18880 28908 18932 28960
rect 20444 28976 20496 29028
rect 21640 28976 21692 29028
rect 23296 28976 23348 29028
rect 23388 28976 23440 29028
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 14096 28704 14148 28756
rect 14832 28704 14884 28756
rect 16764 28747 16816 28756
rect 16764 28713 16773 28747
rect 16773 28713 16807 28747
rect 16807 28713 16816 28747
rect 16764 28704 16816 28713
rect 21272 28704 21324 28756
rect 18420 28636 18472 28688
rect 21180 28679 21232 28688
rect 21180 28645 21189 28679
rect 21189 28645 21223 28679
rect 21223 28645 21232 28679
rect 21180 28636 21232 28645
rect 1308 28568 1360 28620
rect 4160 28568 4212 28620
rect 5632 28611 5684 28620
rect 5632 28577 5641 28611
rect 5641 28577 5675 28611
rect 5675 28577 5684 28611
rect 5632 28568 5684 28577
rect 6552 28611 6604 28620
rect 6552 28577 6561 28611
rect 6561 28577 6595 28611
rect 6595 28577 6604 28611
rect 6552 28568 6604 28577
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 8116 28500 8168 28552
rect 9864 28568 9916 28620
rect 11336 28568 11388 28620
rect 9404 28500 9456 28552
rect 9956 28500 10008 28552
rect 12716 28568 12768 28620
rect 13360 28611 13412 28620
rect 13360 28577 13369 28611
rect 13369 28577 13403 28611
rect 13403 28577 13412 28611
rect 13360 28568 13412 28577
rect 14832 28611 14884 28620
rect 14832 28577 14841 28611
rect 14841 28577 14875 28611
rect 14875 28577 14884 28611
rect 14832 28568 14884 28577
rect 16212 28611 16264 28620
rect 16212 28577 16221 28611
rect 16221 28577 16255 28611
rect 16255 28577 16264 28611
rect 16212 28568 16264 28577
rect 17132 28568 17184 28620
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 22008 28568 22060 28620
rect 22836 28568 22888 28620
rect 15568 28500 15620 28552
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16856 28500 16908 28552
rect 19064 28500 19116 28552
rect 3976 28432 4028 28484
rect 5540 28364 5592 28416
rect 8208 28364 8260 28416
rect 10232 28364 10284 28416
rect 18052 28432 18104 28484
rect 19800 28432 19852 28484
rect 21456 28475 21508 28484
rect 21456 28441 21465 28475
rect 21465 28441 21499 28475
rect 21499 28441 21508 28475
rect 21456 28432 21508 28441
rect 24216 28432 24268 28484
rect 24860 28432 24912 28484
rect 12808 28364 12860 28416
rect 13176 28407 13228 28416
rect 13176 28373 13185 28407
rect 13185 28373 13219 28407
rect 13219 28373 13228 28407
rect 13176 28364 13228 28373
rect 13268 28407 13320 28416
rect 13268 28373 13277 28407
rect 13277 28373 13311 28407
rect 13311 28373 13320 28407
rect 13268 28364 13320 28373
rect 14004 28364 14056 28416
rect 14280 28407 14332 28416
rect 14280 28373 14289 28407
rect 14289 28373 14323 28407
rect 14323 28373 14332 28407
rect 14280 28364 14332 28373
rect 14556 28364 14608 28416
rect 15292 28407 15344 28416
rect 15292 28373 15301 28407
rect 15301 28373 15335 28407
rect 15335 28373 15344 28407
rect 15292 28364 15344 28373
rect 15752 28364 15804 28416
rect 16948 28364 17000 28416
rect 18420 28364 18472 28416
rect 24584 28407 24636 28416
rect 24584 28373 24593 28407
rect 24593 28373 24627 28407
rect 24627 28373 24636 28407
rect 24584 28364 24636 28373
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 1952 28160 2004 28212
rect 3792 28160 3844 28212
rect 10232 28160 10284 28212
rect 13176 28160 13228 28212
rect 15844 28160 15896 28212
rect 18328 28203 18380 28212
rect 18328 28169 18337 28203
rect 18337 28169 18371 28203
rect 18371 28169 18380 28203
rect 18328 28160 18380 28169
rect 20168 28203 20220 28212
rect 20168 28169 20177 28203
rect 20177 28169 20211 28203
rect 20211 28169 20220 28203
rect 20168 28160 20220 28169
rect 22652 28160 22704 28212
rect 3424 28024 3476 28076
rect 3608 28067 3660 28076
rect 3608 28033 3652 28067
rect 3652 28033 3660 28067
rect 3608 28024 3660 28033
rect 8576 27999 8628 28008
rect 8576 27965 8585 27999
rect 8585 27965 8619 27999
rect 8619 27965 8628 27999
rect 8576 27956 8628 27965
rect 8668 27956 8720 28008
rect 11244 27888 11296 27940
rect 9956 27820 10008 27872
rect 13268 28024 13320 28076
rect 16028 27999 16080 28008
rect 16028 27965 16037 27999
rect 16037 27965 16071 27999
rect 16071 27965 16080 27999
rect 16028 27956 16080 27965
rect 16212 27999 16264 28008
rect 16212 27965 16221 27999
rect 16221 27965 16255 27999
rect 16255 27965 16264 27999
rect 18880 28092 18932 28144
rect 17500 28024 17552 28076
rect 20812 28092 20864 28144
rect 21456 28092 21508 28144
rect 24676 28135 24728 28144
rect 24676 28101 24685 28135
rect 24685 28101 24719 28135
rect 24719 28101 24728 28135
rect 24676 28092 24728 28101
rect 16212 27956 16264 27965
rect 18604 27956 18656 28008
rect 12716 27820 12768 27872
rect 14556 27820 14608 27872
rect 15384 27820 15436 27872
rect 15568 27863 15620 27872
rect 15568 27829 15577 27863
rect 15577 27829 15611 27863
rect 15611 27829 15620 27863
rect 15568 27820 15620 27829
rect 19340 28024 19392 28076
rect 22008 28067 22060 28076
rect 22008 28033 22017 28067
rect 22017 28033 22051 28067
rect 22051 28033 22060 28067
rect 22008 28024 22060 28033
rect 19984 27956 20036 28008
rect 24676 27956 24728 28008
rect 18788 27888 18840 27940
rect 17500 27863 17552 27872
rect 17500 27829 17509 27863
rect 17509 27829 17543 27863
rect 17543 27829 17552 27863
rect 17500 27820 17552 27829
rect 18972 27820 19024 27872
rect 19064 27863 19116 27872
rect 19064 27829 19073 27863
rect 19073 27829 19107 27863
rect 19107 27829 19116 27863
rect 19064 27820 19116 27829
rect 25136 27888 25188 27940
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 9864 27616 9916 27668
rect 18328 27616 18380 27668
rect 18788 27616 18840 27668
rect 19340 27616 19392 27668
rect 24216 27659 24268 27668
rect 24216 27625 24225 27659
rect 24225 27625 24259 27659
rect 24259 27625 24268 27659
rect 24216 27616 24268 27625
rect 7840 27548 7892 27600
rect 8300 27591 8352 27600
rect 8300 27557 8309 27591
rect 8309 27557 8343 27591
rect 8343 27557 8352 27591
rect 8300 27548 8352 27557
rect 21088 27548 21140 27600
rect 6552 27480 6604 27532
rect 7564 27412 7616 27464
rect 12808 27480 12860 27532
rect 17132 27480 17184 27532
rect 9956 27412 10008 27464
rect 10968 27412 11020 27464
rect 15476 27412 15528 27464
rect 11428 27387 11480 27396
rect 11428 27353 11437 27387
rect 11437 27353 11471 27387
rect 11471 27353 11480 27387
rect 11428 27344 11480 27353
rect 12716 27344 12768 27396
rect 17040 27412 17092 27464
rect 20536 27523 20588 27532
rect 20536 27489 20545 27523
rect 20545 27489 20579 27523
rect 20579 27489 20588 27523
rect 20536 27480 20588 27489
rect 20628 27523 20680 27532
rect 20628 27489 20637 27523
rect 20637 27489 20671 27523
rect 20671 27489 20680 27523
rect 20628 27480 20680 27489
rect 21916 27523 21968 27532
rect 21916 27489 21925 27523
rect 21925 27489 21959 27523
rect 21959 27489 21968 27523
rect 21916 27480 21968 27489
rect 22744 27480 22796 27532
rect 18236 27344 18288 27396
rect 10232 27276 10284 27328
rect 12900 27319 12952 27328
rect 12900 27285 12909 27319
rect 12909 27285 12943 27319
rect 12943 27285 12952 27319
rect 12900 27276 12952 27285
rect 12992 27276 13044 27328
rect 14096 27276 14148 27328
rect 15016 27276 15068 27328
rect 16396 27319 16448 27328
rect 16396 27285 16405 27319
rect 16405 27285 16439 27319
rect 16439 27285 16448 27319
rect 16396 27276 16448 27285
rect 18604 27276 18656 27328
rect 22192 27387 22244 27396
rect 22192 27353 22201 27387
rect 22201 27353 22235 27387
rect 22235 27353 22244 27387
rect 22192 27344 22244 27353
rect 22284 27344 22336 27396
rect 22652 27344 22704 27396
rect 25044 27344 25096 27396
rect 23020 27276 23072 27328
rect 23112 27276 23164 27328
rect 25228 27319 25280 27328
rect 25228 27285 25237 27319
rect 25237 27285 25271 27319
rect 25271 27285 25280 27319
rect 25228 27276 25280 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 3884 27072 3936 27124
rect 3332 26936 3384 26988
rect 3516 26936 3568 26988
rect 4344 26868 4396 26920
rect 7564 27004 7616 27056
rect 10048 27004 10100 27056
rect 11520 27072 11572 27124
rect 16580 27072 16632 27124
rect 22560 27072 22612 27124
rect 22744 27072 22796 27124
rect 13084 27004 13136 27056
rect 14096 27004 14148 27056
rect 16396 27004 16448 27056
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 10968 26936 11020 26988
rect 18144 27004 18196 27056
rect 18420 27004 18472 27056
rect 21364 27004 21416 27056
rect 24584 27072 24636 27124
rect 23020 27004 23072 27056
rect 23572 27004 23624 27056
rect 24952 27004 25004 27056
rect 3700 26800 3752 26852
rect 7840 26868 7892 26920
rect 8668 26868 8720 26920
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 12808 26911 12860 26920
rect 12808 26877 12817 26911
rect 12817 26877 12851 26911
rect 12851 26877 12860 26911
rect 12808 26868 12860 26877
rect 12900 26868 12952 26920
rect 8300 26843 8352 26852
rect 8300 26809 8309 26843
rect 8309 26809 8343 26843
rect 8343 26809 8352 26843
rect 8300 26800 8352 26809
rect 9680 26800 9732 26852
rect 10324 26800 10376 26852
rect 10508 26732 10560 26784
rect 12992 26732 13044 26784
rect 14372 26732 14424 26784
rect 17408 26800 17460 26852
rect 18144 26868 18196 26920
rect 19340 26868 19392 26920
rect 19800 26868 19852 26920
rect 21180 26868 21232 26920
rect 21456 26868 21508 26920
rect 22008 26868 22060 26920
rect 20628 26800 20680 26852
rect 22560 26800 22612 26852
rect 23204 26868 23256 26920
rect 18328 26732 18380 26784
rect 19524 26775 19576 26784
rect 19524 26741 19533 26775
rect 19533 26741 19567 26775
rect 19567 26741 19576 26775
rect 19524 26732 19576 26741
rect 23848 26732 23900 26784
rect 24584 26775 24636 26784
rect 24584 26741 24593 26775
rect 24593 26741 24627 26775
rect 24627 26741 24636 26775
rect 24584 26732 24636 26741
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 4068 26571 4120 26580
rect 4068 26537 4077 26571
rect 4077 26537 4111 26571
rect 4111 26537 4120 26571
rect 4068 26528 4120 26537
rect 8576 26528 8628 26580
rect 16672 26528 16724 26580
rect 17776 26528 17828 26580
rect 22192 26528 22244 26580
rect 22652 26528 22704 26580
rect 24584 26528 24636 26580
rect 14832 26460 14884 26512
rect 17500 26503 17552 26512
rect 17500 26469 17509 26503
rect 17509 26469 17543 26503
rect 17543 26469 17552 26503
rect 17500 26460 17552 26469
rect 17868 26460 17920 26512
rect 19708 26460 19760 26512
rect 22560 26460 22612 26512
rect 23572 26460 23624 26512
rect 25228 26460 25280 26512
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 8300 26392 8352 26444
rect 9128 26435 9180 26444
rect 9128 26401 9137 26435
rect 9137 26401 9171 26435
rect 9171 26401 9180 26435
rect 9128 26392 9180 26401
rect 10232 26435 10284 26444
rect 10232 26401 10241 26435
rect 10241 26401 10275 26435
rect 10275 26401 10284 26435
rect 10232 26392 10284 26401
rect 11244 26392 11296 26444
rect 13544 26392 13596 26444
rect 13912 26392 13964 26444
rect 18972 26392 19024 26444
rect 20168 26392 20220 26444
rect 20628 26435 20680 26444
rect 20628 26401 20637 26435
rect 20637 26401 20671 26435
rect 20671 26401 20680 26435
rect 20628 26392 20680 26401
rect 21456 26392 21508 26444
rect 21640 26392 21692 26444
rect 24584 26392 24636 26444
rect 2044 26324 2096 26376
rect 9956 26367 10008 26376
rect 9956 26333 9965 26367
rect 9965 26333 9999 26367
rect 9999 26333 10008 26367
rect 9956 26324 10008 26333
rect 14280 26324 14332 26376
rect 15384 26367 15436 26376
rect 15384 26333 15393 26367
rect 15393 26333 15427 26367
rect 15427 26333 15436 26367
rect 15384 26324 15436 26333
rect 20260 26324 20312 26376
rect 22284 26324 22336 26376
rect 24216 26324 24268 26376
rect 2780 26299 2832 26308
rect 2780 26265 2789 26299
rect 2789 26265 2823 26299
rect 2823 26265 2832 26299
rect 2780 26256 2832 26265
rect 7472 26256 7524 26308
rect 8668 26299 8720 26308
rect 8668 26265 8677 26299
rect 8677 26265 8711 26299
rect 8711 26265 8720 26299
rect 8668 26256 8720 26265
rect 8760 26256 8812 26308
rect 13360 26256 13412 26308
rect 13544 26256 13596 26308
rect 15200 26256 15252 26308
rect 7656 26188 7708 26240
rect 12164 26231 12216 26240
rect 12164 26197 12173 26231
rect 12173 26197 12207 26231
rect 12207 26197 12216 26231
rect 12164 26188 12216 26197
rect 12532 26231 12584 26240
rect 12532 26197 12541 26231
rect 12541 26197 12575 26231
rect 12575 26197 12584 26231
rect 12532 26188 12584 26197
rect 14096 26188 14148 26240
rect 14832 26188 14884 26240
rect 17776 26256 17828 26308
rect 21180 26256 21232 26308
rect 21824 26188 21876 26240
rect 24492 26256 24544 26308
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 1768 25984 1820 26036
rect 7564 25984 7616 26036
rect 8760 25984 8812 26036
rect 3516 25916 3568 25968
rect 4068 25916 4120 25968
rect 10508 25984 10560 26036
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 2872 25848 2924 25900
rect 12532 25916 12584 25968
rect 2780 25780 2832 25832
rect 3608 25780 3660 25832
rect 5448 25848 5500 25900
rect 8484 25848 8536 25900
rect 6184 25780 6236 25832
rect 7840 25780 7892 25832
rect 9404 25848 9456 25900
rect 15384 25984 15436 26036
rect 15568 25984 15620 26036
rect 14832 25959 14884 25968
rect 14832 25925 14841 25959
rect 14841 25925 14875 25959
rect 14875 25925 14884 25959
rect 14832 25916 14884 25925
rect 18696 25984 18748 26036
rect 19340 26027 19392 26036
rect 19340 25993 19349 26027
rect 19349 25993 19383 26027
rect 19383 25993 19392 26027
rect 19340 25984 19392 25993
rect 19524 25984 19576 26036
rect 20352 26027 20404 26036
rect 20352 25993 20361 26027
rect 20361 25993 20395 26027
rect 20395 25993 20404 26027
rect 20352 25984 20404 25993
rect 21364 25984 21416 26036
rect 22284 25984 22336 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 21548 25916 21600 25968
rect 25136 25916 25188 25968
rect 25412 25916 25464 25968
rect 3424 25755 3476 25764
rect 3424 25721 3433 25755
rect 3433 25721 3467 25755
rect 3467 25721 3476 25755
rect 3424 25712 3476 25721
rect 8576 25712 8628 25764
rect 9864 25780 9916 25832
rect 11796 25780 11848 25832
rect 14372 25780 14424 25832
rect 14464 25823 14516 25832
rect 14464 25789 14473 25823
rect 14473 25789 14507 25823
rect 14507 25789 14516 25823
rect 14464 25780 14516 25789
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 4252 25687 4304 25696
rect 4252 25653 4261 25687
rect 4261 25653 4295 25687
rect 4295 25653 4304 25687
rect 4252 25644 4304 25653
rect 11336 25644 11388 25696
rect 11428 25644 11480 25696
rect 15476 25712 15528 25764
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 18236 25780 18288 25832
rect 22192 25848 22244 25900
rect 23388 25848 23440 25900
rect 23848 25848 23900 25900
rect 21640 25780 21692 25832
rect 22284 25780 22336 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 18972 25712 19024 25764
rect 22100 25712 22152 25764
rect 22836 25712 22888 25764
rect 23756 25712 23808 25764
rect 15200 25644 15252 25696
rect 21180 25644 21232 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 7472 25440 7524 25492
rect 7656 25440 7708 25492
rect 8760 25440 8812 25492
rect 9036 25440 9088 25492
rect 11520 25440 11572 25492
rect 12440 25440 12492 25492
rect 7656 25304 7708 25356
rect 4068 25279 4120 25288
rect 4068 25245 4086 25279
rect 4086 25245 4120 25279
rect 4068 25236 4120 25245
rect 9404 25347 9456 25356
rect 9404 25313 9413 25347
rect 9413 25313 9447 25347
rect 9447 25313 9456 25347
rect 9404 25304 9456 25313
rect 9680 25304 9732 25356
rect 11428 25304 11480 25356
rect 8392 25236 8444 25288
rect 10784 25236 10836 25288
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 16764 25440 16816 25492
rect 17776 25440 17828 25492
rect 18236 25440 18288 25492
rect 22468 25440 22520 25492
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 25228 25483 25280 25492
rect 25228 25449 25237 25483
rect 25237 25449 25271 25483
rect 25271 25449 25280 25483
rect 25228 25440 25280 25449
rect 25504 25483 25556 25492
rect 25504 25449 25513 25483
rect 25513 25449 25547 25483
rect 25547 25449 25556 25483
rect 25504 25440 25556 25449
rect 12808 25304 12860 25356
rect 13636 25304 13688 25356
rect 15384 25304 15436 25356
rect 24952 25372 25004 25424
rect 16672 25304 16724 25356
rect 19064 25304 19116 25356
rect 20076 25347 20128 25356
rect 20076 25313 20085 25347
rect 20085 25313 20119 25347
rect 20119 25313 20128 25347
rect 20076 25304 20128 25313
rect 21088 25304 21140 25356
rect 22652 25304 22704 25356
rect 23204 25304 23256 25356
rect 12532 25236 12584 25288
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 19432 25236 19484 25288
rect 21640 25236 21692 25288
rect 22836 25236 22888 25288
rect 3976 25100 4028 25152
rect 6644 25100 6696 25152
rect 8576 25143 8628 25152
rect 8576 25109 8585 25143
rect 8585 25109 8619 25143
rect 8619 25109 8628 25143
rect 8576 25100 8628 25109
rect 13636 25168 13688 25220
rect 17776 25168 17828 25220
rect 22376 25168 22428 25220
rect 11980 25100 12032 25152
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 12808 25100 12860 25152
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 16856 25100 16908 25152
rect 17040 25100 17092 25152
rect 17868 25100 17920 25152
rect 18328 25100 18380 25152
rect 18512 25100 18564 25152
rect 18696 25100 18748 25152
rect 19432 25143 19484 25152
rect 19432 25109 19441 25143
rect 19441 25109 19475 25143
rect 19475 25109 19484 25143
rect 19432 25100 19484 25109
rect 23940 25143 23992 25152
rect 23940 25109 23949 25143
rect 23949 25109 23983 25143
rect 23983 25109 23992 25143
rect 23940 25100 23992 25109
rect 24032 25100 24084 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 4252 24896 4304 24948
rect 7840 24896 7892 24948
rect 12624 24896 12676 24948
rect 16856 24939 16908 24948
rect 16856 24905 16865 24939
rect 16865 24905 16899 24939
rect 16899 24905 16908 24939
rect 16856 24896 16908 24905
rect 17684 24896 17736 24948
rect 18512 24939 18564 24948
rect 18512 24905 18521 24939
rect 18521 24905 18555 24939
rect 18555 24905 18564 24939
rect 18512 24896 18564 24905
rect 19892 24939 19944 24948
rect 19892 24905 19901 24939
rect 19901 24905 19935 24939
rect 19935 24905 19944 24939
rect 19892 24896 19944 24905
rect 7472 24828 7524 24880
rect 5816 24760 5868 24812
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 7748 24760 7800 24812
rect 6000 24692 6052 24744
rect 8116 24735 8168 24744
rect 8116 24701 8125 24735
rect 8125 24701 8159 24735
rect 8159 24701 8168 24735
rect 8116 24692 8168 24701
rect 9312 24735 9364 24744
rect 9312 24701 9321 24735
rect 9321 24701 9355 24735
rect 9355 24701 9364 24735
rect 9312 24692 9364 24701
rect 12440 24760 12492 24812
rect 12900 24828 12952 24880
rect 13084 24828 13136 24880
rect 13544 24760 13596 24812
rect 13820 24803 13872 24812
rect 13820 24769 13829 24803
rect 13829 24769 13863 24803
rect 13863 24769 13872 24803
rect 13820 24760 13872 24769
rect 10140 24692 10192 24744
rect 12992 24735 13044 24744
rect 12992 24701 13001 24735
rect 13001 24701 13035 24735
rect 13035 24701 13044 24735
rect 12992 24692 13044 24701
rect 15016 24760 15068 24812
rect 16396 24828 16448 24880
rect 17132 24828 17184 24880
rect 23204 24871 23256 24880
rect 23204 24837 23213 24871
rect 23213 24837 23247 24871
rect 23247 24837 23256 24871
rect 23204 24828 23256 24837
rect 24492 24828 24544 24880
rect 25228 24828 25280 24880
rect 14372 24692 14424 24744
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17868 24760 17920 24812
rect 18328 24760 18380 24812
rect 18880 24760 18932 24812
rect 20628 24760 20680 24812
rect 22836 24760 22888 24812
rect 25504 24760 25556 24812
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 17776 24692 17828 24744
rect 18788 24692 18840 24744
rect 20536 24692 20588 24744
rect 8392 24624 8444 24676
rect 3976 24556 4028 24608
rect 5816 24599 5868 24608
rect 5816 24565 5825 24599
rect 5825 24565 5859 24599
rect 5859 24565 5868 24599
rect 5816 24556 5868 24565
rect 7748 24556 7800 24608
rect 12624 24624 12676 24676
rect 11152 24556 11204 24608
rect 12256 24556 12308 24608
rect 12900 24556 12952 24608
rect 15108 24624 15160 24676
rect 13728 24556 13780 24608
rect 18880 24624 18932 24676
rect 20444 24624 20496 24676
rect 20628 24624 20680 24676
rect 24676 24735 24728 24744
rect 24676 24701 24685 24735
rect 24685 24701 24719 24735
rect 24719 24701 24728 24735
rect 24676 24692 24728 24701
rect 25136 24667 25188 24676
rect 25136 24633 25145 24667
rect 25145 24633 25179 24667
rect 25179 24633 25188 24667
rect 25136 24624 25188 24633
rect 16396 24599 16448 24608
rect 16396 24565 16405 24599
rect 16405 24565 16439 24599
rect 16439 24565 16448 24599
rect 16396 24556 16448 24565
rect 18512 24556 18564 24608
rect 23388 24556 23440 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 3332 24352 3384 24404
rect 4436 24352 4488 24404
rect 6184 24395 6236 24404
rect 6184 24361 6193 24395
rect 6193 24361 6227 24395
rect 6227 24361 6236 24395
rect 6184 24352 6236 24361
rect 8484 24352 8536 24404
rect 9312 24352 9364 24404
rect 10232 24352 10284 24404
rect 6368 24284 6420 24336
rect 8576 24284 8628 24336
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 4252 24216 4304 24225
rect 9864 24216 9916 24268
rect 11060 24216 11112 24268
rect 12164 24284 12216 24336
rect 13728 24284 13780 24336
rect 12808 24216 12860 24268
rect 15384 24352 15436 24404
rect 15936 24352 15988 24404
rect 20720 24352 20772 24404
rect 24676 24284 24728 24336
rect 2780 24148 2832 24200
rect 3516 24148 3568 24200
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 7104 24148 7156 24200
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 12624 24148 12676 24200
rect 4528 24080 4580 24132
rect 5816 24080 5868 24132
rect 6552 24080 6604 24132
rect 9036 24080 9088 24132
rect 16948 24216 17000 24268
rect 17040 24259 17092 24268
rect 17040 24225 17049 24259
rect 17049 24225 17083 24259
rect 17083 24225 17092 24259
rect 17040 24216 17092 24225
rect 17316 24216 17368 24268
rect 22836 24216 22888 24268
rect 24860 24216 24912 24268
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 1860 24012 1912 24064
rect 8760 24012 8812 24064
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 13820 24080 13872 24132
rect 14740 24080 14792 24132
rect 21732 24148 21784 24200
rect 23296 24148 23348 24200
rect 24400 24148 24452 24200
rect 18788 24080 18840 24132
rect 19892 24080 19944 24132
rect 21364 24080 21416 24132
rect 24952 24123 25004 24132
rect 24952 24089 24961 24123
rect 24961 24089 24995 24123
rect 24995 24089 25004 24123
rect 24952 24080 25004 24089
rect 10692 24012 10744 24064
rect 10968 24012 11020 24064
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 12072 24012 12124 24064
rect 16672 24012 16724 24064
rect 17500 24012 17552 24064
rect 20260 24012 20312 24064
rect 22100 24055 22152 24064
rect 22100 24021 22109 24055
rect 22109 24021 22143 24055
rect 22143 24021 22152 24055
rect 22100 24012 22152 24021
rect 22376 24012 22428 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 6000 23851 6052 23860
rect 6000 23817 6009 23851
rect 6009 23817 6043 23851
rect 6043 23817 6052 23851
rect 6000 23808 6052 23817
rect 6552 23808 6604 23860
rect 7656 23808 7708 23860
rect 9956 23808 10008 23860
rect 10692 23808 10744 23860
rect 11244 23808 11296 23860
rect 12072 23808 12124 23860
rect 12348 23808 12400 23860
rect 13544 23808 13596 23860
rect 13912 23851 13964 23860
rect 13912 23817 13921 23851
rect 13921 23817 13955 23851
rect 13955 23817 13964 23851
rect 13912 23808 13964 23817
rect 18696 23808 18748 23860
rect 19892 23808 19944 23860
rect 1768 23715 1820 23724
rect 1768 23681 1777 23715
rect 1777 23681 1811 23715
rect 1811 23681 1820 23715
rect 1768 23672 1820 23681
rect 9772 23740 9824 23792
rect 10508 23740 10560 23792
rect 9036 23672 9088 23724
rect 11244 23672 11296 23724
rect 20536 23808 20588 23860
rect 20628 23740 20680 23792
rect 23480 23740 23532 23792
rect 24492 23740 24544 23792
rect 1308 23604 1360 23656
rect 3976 23604 4028 23656
rect 7564 23604 7616 23656
rect 8576 23604 8628 23656
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 11704 23604 11756 23656
rect 12440 23604 12492 23656
rect 13452 23604 13504 23656
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 18604 23604 18656 23656
rect 19800 23604 19852 23656
rect 9956 23536 10008 23588
rect 16488 23536 16540 23588
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 21364 23672 21416 23724
rect 22008 23672 22060 23724
rect 22836 23672 22888 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 21364 23536 21416 23588
rect 24308 23536 24360 23588
rect 5724 23468 5776 23520
rect 6828 23468 6880 23520
rect 10140 23468 10192 23520
rect 10784 23468 10836 23520
rect 11796 23468 11848 23520
rect 17500 23468 17552 23520
rect 20812 23468 20864 23520
rect 23664 23468 23716 23520
rect 24676 23511 24728 23520
rect 24676 23477 24685 23511
rect 24685 23477 24719 23511
rect 24719 23477 24728 23511
rect 24676 23468 24728 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 2044 23307 2096 23316
rect 2044 23273 2053 23307
rect 2053 23273 2087 23307
rect 2087 23273 2096 23307
rect 2044 23264 2096 23273
rect 2872 23264 2924 23316
rect 7564 23307 7616 23316
rect 7564 23273 7573 23307
rect 7573 23273 7607 23307
rect 7607 23273 7616 23307
rect 7564 23264 7616 23273
rect 2872 23128 2924 23180
rect 3332 23128 3384 23180
rect 5724 23128 5776 23180
rect 6460 23128 6512 23180
rect 3792 22992 3844 23044
rect 3976 23060 4028 23112
rect 4344 23060 4396 23112
rect 7840 23128 7892 23180
rect 9036 23264 9088 23316
rect 14648 23264 14700 23316
rect 16028 23307 16080 23316
rect 16028 23273 16037 23307
rect 16037 23273 16071 23307
rect 16071 23273 16080 23307
rect 16028 23264 16080 23273
rect 20076 23264 20128 23316
rect 20444 23264 20496 23316
rect 21364 23264 21416 23316
rect 19340 23196 19392 23248
rect 24676 23196 24728 23248
rect 12164 23128 12216 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 14280 23171 14332 23180
rect 14280 23137 14289 23171
rect 14289 23137 14323 23171
rect 14323 23137 14332 23171
rect 14280 23128 14332 23137
rect 15292 23128 15344 23180
rect 18604 23128 18656 23180
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 10876 23060 10928 23112
rect 5080 22992 5132 23044
rect 3332 22924 3384 22976
rect 5448 22924 5500 22976
rect 10692 23035 10744 23044
rect 10692 23001 10701 23035
rect 10701 23001 10735 23035
rect 10735 23001 10744 23035
rect 10692 22992 10744 23001
rect 10784 22992 10836 23044
rect 16396 23060 16448 23112
rect 22744 23103 22796 23112
rect 22744 23069 22753 23103
rect 22753 23069 22787 23103
rect 22787 23069 22796 23103
rect 22744 23060 22796 23069
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 12440 22992 12492 23044
rect 7472 22924 7524 22976
rect 9772 22924 9824 22976
rect 11704 22924 11756 22976
rect 12256 22924 12308 22976
rect 13912 22992 13964 23044
rect 13084 22924 13136 22976
rect 15936 22992 15988 23044
rect 16212 22924 16264 22976
rect 16396 22924 16448 22976
rect 19340 22992 19392 23044
rect 19984 22992 20036 23044
rect 21364 22992 21416 23044
rect 23388 22992 23440 23044
rect 23480 22924 23532 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 1768 22720 1820 22772
rect 8760 22720 8812 22772
rect 5908 22652 5960 22704
rect 2872 22584 2924 22636
rect 6920 22584 6972 22636
rect 6000 22516 6052 22568
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 7564 22584 7616 22636
rect 9956 22720 10008 22772
rect 10048 22652 10100 22704
rect 12072 22652 12124 22704
rect 15200 22763 15252 22772
rect 15200 22729 15209 22763
rect 15209 22729 15243 22763
rect 15243 22729 15252 22763
rect 15200 22720 15252 22729
rect 15292 22720 15344 22772
rect 15568 22720 15620 22772
rect 16212 22763 16264 22772
rect 16212 22729 16221 22763
rect 16221 22729 16255 22763
rect 16255 22729 16264 22763
rect 16212 22720 16264 22729
rect 16488 22720 16540 22772
rect 16580 22720 16632 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 15844 22652 15896 22704
rect 16396 22695 16448 22704
rect 16396 22661 16405 22695
rect 16405 22661 16439 22695
rect 16439 22661 16448 22695
rect 16396 22652 16448 22661
rect 20352 22720 20404 22772
rect 23572 22720 23624 22772
rect 18604 22695 18656 22704
rect 18604 22661 18613 22695
rect 18613 22661 18647 22695
rect 18647 22661 18656 22695
rect 18604 22652 18656 22661
rect 19708 22695 19760 22704
rect 19708 22661 19717 22695
rect 19717 22661 19751 22695
rect 19751 22661 19760 22695
rect 19708 22652 19760 22661
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 11152 22516 11204 22568
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 13084 22584 13136 22593
rect 13820 22584 13872 22636
rect 15200 22584 15252 22636
rect 19340 22584 19392 22636
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 23388 22584 23440 22636
rect 4436 22448 4488 22500
rect 6644 22448 6696 22500
rect 9404 22448 9456 22500
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 15936 22516 15988 22568
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 19800 22516 19852 22525
rect 21640 22516 21692 22568
rect 24492 22720 24544 22772
rect 25320 22720 25372 22772
rect 17868 22448 17920 22500
rect 4252 22380 4304 22432
rect 7472 22380 7524 22432
rect 10508 22380 10560 22432
rect 12808 22380 12860 22432
rect 14740 22423 14792 22432
rect 14740 22389 14749 22423
rect 14749 22389 14783 22423
rect 14783 22389 14792 22423
rect 14740 22380 14792 22389
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 13268 22176 13320 22228
rect 13544 22176 13596 22228
rect 16396 22219 16448 22228
rect 16396 22185 16405 22219
rect 16405 22185 16439 22219
rect 16439 22185 16448 22219
rect 16396 22176 16448 22185
rect 11428 22151 11480 22160
rect 11428 22117 11437 22151
rect 11437 22117 11471 22151
rect 11471 22117 11480 22151
rect 11428 22108 11480 22117
rect 11796 22108 11848 22160
rect 12256 22108 12308 22160
rect 14280 22083 14332 22092
rect 14280 22049 14289 22083
rect 14289 22049 14323 22083
rect 14323 22049 14332 22083
rect 14280 22040 14332 22049
rect 14556 22040 14608 22092
rect 14924 22040 14976 22092
rect 16028 22083 16080 22092
rect 16028 22049 16037 22083
rect 16037 22049 16071 22083
rect 16071 22049 16080 22083
rect 16028 22040 16080 22049
rect 16856 22040 16908 22092
rect 13360 21972 13412 22024
rect 4528 21836 4580 21888
rect 10600 21836 10652 21888
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 11520 21836 11572 21888
rect 12900 21836 12952 21888
rect 14188 21904 14240 21956
rect 14648 21904 14700 21956
rect 16396 21904 16448 21956
rect 17040 21972 17092 22024
rect 17776 22040 17828 22092
rect 18512 22083 18564 22092
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 20260 22176 20312 22228
rect 21364 22176 21416 22228
rect 19340 22040 19392 22092
rect 19800 22040 19852 22092
rect 22008 22083 22060 22092
rect 22008 22049 22017 22083
rect 22017 22049 22051 22083
rect 22051 22049 22060 22083
rect 22008 22040 22060 22049
rect 24308 22040 24360 22092
rect 15476 21836 15528 21888
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 23388 21972 23440 22024
rect 24124 21972 24176 22024
rect 19800 21904 19852 21956
rect 21456 21904 21508 21956
rect 22284 21947 22336 21956
rect 22284 21913 22293 21947
rect 22293 21913 22327 21947
rect 22327 21913 22336 21947
rect 22284 21904 22336 21913
rect 19524 21836 19576 21888
rect 19892 21836 19944 21888
rect 21272 21836 21324 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 7104 21675 7156 21684
rect 7104 21641 7113 21675
rect 7113 21641 7147 21675
rect 7147 21641 7156 21675
rect 7104 21632 7156 21641
rect 9772 21632 9824 21684
rect 11980 21632 12032 21684
rect 13820 21632 13872 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 15384 21632 15436 21684
rect 17224 21632 17276 21684
rect 7656 21564 7708 21616
rect 1860 21496 1912 21548
rect 4160 21496 4212 21548
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 8944 21496 8996 21548
rect 1308 21428 1360 21480
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 4068 21428 4120 21480
rect 7656 21471 7708 21480
rect 7656 21437 7665 21471
rect 7665 21437 7699 21471
rect 7699 21437 7708 21471
rect 7656 21428 7708 21437
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 9036 21428 9088 21480
rect 12808 21564 12860 21616
rect 18696 21632 18748 21684
rect 21272 21632 21324 21684
rect 22560 21675 22612 21684
rect 22560 21641 22569 21675
rect 22569 21641 22603 21675
rect 22603 21641 22612 21675
rect 22560 21632 22612 21641
rect 23388 21632 23440 21684
rect 23572 21632 23624 21684
rect 13912 21496 13964 21548
rect 3792 21403 3844 21412
rect 3792 21369 3801 21403
rect 3801 21369 3835 21403
rect 3835 21369 3844 21403
rect 3792 21360 3844 21369
rect 6920 21360 6972 21412
rect 11060 21428 11112 21480
rect 12348 21471 12400 21480
rect 12348 21437 12357 21471
rect 12357 21437 12391 21471
rect 12391 21437 12400 21471
rect 12348 21428 12400 21437
rect 13728 21428 13780 21480
rect 16120 21496 16172 21548
rect 21088 21564 21140 21616
rect 22008 21564 22060 21616
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 14648 21428 14700 21480
rect 15384 21471 15436 21480
rect 15384 21437 15393 21471
rect 15393 21437 15427 21471
rect 15427 21437 15436 21471
rect 15384 21428 15436 21437
rect 10784 21360 10836 21412
rect 5816 21292 5868 21344
rect 7564 21292 7616 21344
rect 8208 21292 8260 21344
rect 11336 21360 11388 21412
rect 17408 21496 17460 21548
rect 23296 21496 23348 21548
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 17592 21428 17644 21480
rect 19524 21428 19576 21480
rect 20628 21428 20680 21480
rect 20996 21428 21048 21480
rect 22284 21428 22336 21480
rect 22468 21360 22520 21412
rect 13820 21292 13872 21344
rect 16028 21335 16080 21344
rect 16028 21301 16037 21335
rect 16037 21301 16071 21335
rect 16071 21301 16080 21335
rect 16028 21292 16080 21301
rect 16396 21292 16448 21344
rect 19524 21292 19576 21344
rect 20444 21335 20496 21344
rect 20444 21301 20453 21335
rect 20453 21301 20487 21335
rect 20487 21301 20496 21335
rect 20444 21292 20496 21301
rect 20812 21292 20864 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 2872 21088 2924 21140
rect 7288 21088 7340 21140
rect 9128 21088 9180 21140
rect 10048 21088 10100 21140
rect 12256 21020 12308 21072
rect 8208 20952 8260 21004
rect 10692 20952 10744 21004
rect 11244 20952 11296 21004
rect 11520 20952 11572 21004
rect 11980 20952 12032 21004
rect 4068 20884 4120 20936
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 1768 20748 1820 20800
rect 2780 20748 2832 20800
rect 4712 20748 4764 20800
rect 8484 20816 8536 20868
rect 10048 20859 10100 20868
rect 10048 20825 10057 20859
rect 10057 20825 10091 20859
rect 10091 20825 10100 20859
rect 10048 20816 10100 20825
rect 15016 20884 15068 20936
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15752 20884 15804 20893
rect 10416 20748 10468 20800
rect 10692 20748 10744 20800
rect 16396 21088 16448 21140
rect 17132 21088 17184 21140
rect 16120 21063 16172 21072
rect 16120 21029 16129 21063
rect 16129 21029 16163 21063
rect 16163 21029 16172 21063
rect 20168 21088 20220 21140
rect 21456 21088 21508 21140
rect 16120 21020 16172 21029
rect 17132 20952 17184 21004
rect 19800 20952 19852 21004
rect 20536 20952 20588 21004
rect 24860 20952 24912 21004
rect 17592 20927 17644 20936
rect 17592 20893 17601 20927
rect 17601 20893 17635 20927
rect 17635 20893 17644 20927
rect 17592 20884 17644 20893
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 21456 20884 21508 20936
rect 25412 20884 25464 20936
rect 12348 20748 12400 20800
rect 15568 20791 15620 20800
rect 15568 20757 15577 20791
rect 15577 20757 15611 20791
rect 15611 20757 15620 20791
rect 15568 20748 15620 20757
rect 19432 20816 19484 20868
rect 24860 20816 24912 20868
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 6552 20544 6604 20596
rect 8852 20544 8904 20596
rect 8944 20544 8996 20596
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 4344 20476 4396 20528
rect 7104 20476 7156 20528
rect 9036 20476 9088 20528
rect 6552 20451 6604 20460
rect 6552 20417 6561 20451
rect 6561 20417 6595 20451
rect 6595 20417 6604 20451
rect 6552 20408 6604 20417
rect 8668 20408 8720 20460
rect 5724 20340 5776 20392
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 5816 20204 5868 20256
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 9036 20204 9088 20256
rect 9220 20383 9272 20392
rect 9220 20349 9229 20383
rect 9229 20349 9263 20383
rect 9263 20349 9272 20383
rect 9220 20340 9272 20349
rect 11520 20476 11572 20528
rect 11796 20476 11848 20528
rect 12532 20476 12584 20528
rect 13912 20476 13964 20528
rect 14280 20476 14332 20528
rect 19340 20544 19392 20596
rect 23388 20476 23440 20528
rect 11704 20408 11756 20460
rect 13636 20408 13688 20460
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 19432 20408 19484 20460
rect 24032 20408 24084 20460
rect 24216 20408 24268 20460
rect 12164 20272 12216 20324
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 21640 20340 21692 20392
rect 23296 20340 23348 20392
rect 13912 20272 13964 20324
rect 14648 20315 14700 20324
rect 14648 20281 14657 20315
rect 14657 20281 14691 20315
rect 14691 20281 14700 20315
rect 14648 20272 14700 20281
rect 20996 20272 21048 20324
rect 13636 20204 13688 20256
rect 14004 20204 14056 20256
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 18788 20204 18840 20256
rect 19800 20204 19852 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 5080 20043 5132 20052
rect 5080 20009 5089 20043
rect 5089 20009 5123 20043
rect 5123 20009 5132 20043
rect 5080 20000 5132 20009
rect 5724 20000 5776 20052
rect 6552 20000 6604 20052
rect 11704 20043 11756 20052
rect 11704 20009 11713 20043
rect 11713 20009 11747 20043
rect 11747 20009 11756 20043
rect 11704 20000 11756 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 18880 20000 18932 20052
rect 19156 20000 19208 20052
rect 20260 20043 20312 20052
rect 20260 20009 20269 20043
rect 20269 20009 20303 20043
rect 20303 20009 20312 20043
rect 20260 20000 20312 20009
rect 8300 19864 8352 19916
rect 8852 19864 8904 19916
rect 11796 19864 11848 19916
rect 7104 19796 7156 19848
rect 7840 19796 7892 19848
rect 8944 19796 8996 19848
rect 11704 19796 11756 19848
rect 12164 19864 12216 19916
rect 13912 19864 13964 19916
rect 12440 19796 12492 19848
rect 18328 19932 18380 19984
rect 19984 19932 20036 19984
rect 16028 19864 16080 19916
rect 19156 19864 19208 19916
rect 24952 19864 25004 19916
rect 17868 19796 17920 19848
rect 18972 19796 19024 19848
rect 20720 19796 20772 19848
rect 25044 19796 25096 19848
rect 7380 19660 7432 19712
rect 7656 19728 7708 19780
rect 8668 19703 8720 19712
rect 8668 19669 8677 19703
rect 8677 19669 8711 19703
rect 8711 19669 8720 19703
rect 8668 19660 8720 19669
rect 8944 19660 8996 19712
rect 11796 19728 11848 19780
rect 11980 19728 12032 19780
rect 14188 19728 14240 19780
rect 10968 19660 11020 19712
rect 13728 19660 13780 19712
rect 17592 19728 17644 19780
rect 18604 19728 18656 19780
rect 23664 19728 23716 19780
rect 14832 19660 14884 19712
rect 18972 19660 19024 19712
rect 19524 19660 19576 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 1492 19456 1544 19508
rect 4160 19456 4212 19508
rect 7840 19456 7892 19508
rect 9404 19456 9456 19508
rect 7104 19388 7156 19440
rect 9312 19388 9364 19440
rect 12808 19456 12860 19508
rect 14096 19456 14148 19508
rect 17316 19456 17368 19508
rect 13728 19388 13780 19440
rect 3608 19320 3660 19372
rect 6276 19320 6328 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8392 19320 8444 19372
rect 8852 19320 8904 19372
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 9220 19252 9272 19304
rect 11980 19320 12032 19372
rect 14648 19320 14700 19372
rect 17592 19388 17644 19440
rect 19248 19388 19300 19440
rect 20260 19456 20312 19508
rect 20536 19388 20588 19440
rect 21180 19499 21232 19508
rect 21180 19465 21189 19499
rect 21189 19465 21223 19499
rect 21223 19465 21232 19499
rect 21180 19456 21232 19465
rect 21916 19456 21968 19508
rect 21456 19388 21508 19440
rect 23572 19388 23624 19440
rect 19524 19320 19576 19372
rect 19892 19320 19944 19372
rect 7564 19116 7616 19168
rect 10232 19116 10284 19168
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 13360 19184 13412 19236
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 13912 19184 13964 19236
rect 17684 19252 17736 19304
rect 19340 19252 19392 19304
rect 21272 19252 21324 19304
rect 21916 19252 21968 19304
rect 22008 19295 22060 19304
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 14832 19184 14884 19236
rect 19248 19184 19300 19236
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 20720 19116 20772 19168
rect 24400 19116 24452 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 5172 18912 5224 18964
rect 10600 18912 10652 18964
rect 11244 18912 11296 18964
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 14188 18912 14240 18964
rect 8944 18887 8996 18896
rect 8944 18853 8953 18887
rect 8953 18853 8987 18887
rect 8987 18853 8996 18887
rect 8944 18844 8996 18853
rect 1308 18776 1360 18828
rect 6184 18776 6236 18828
rect 11060 18776 11112 18828
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 11336 18844 11388 18896
rect 13912 18844 13964 18896
rect 12716 18776 12768 18828
rect 14372 18776 14424 18828
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 13820 18708 13872 18760
rect 17684 18912 17736 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 22284 18912 22336 18964
rect 24400 18955 24452 18964
rect 24400 18921 24409 18955
rect 24409 18921 24443 18955
rect 24443 18921 24452 18955
rect 24400 18912 24452 18921
rect 18972 18844 19024 18896
rect 16488 18776 16540 18828
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 19064 18708 19116 18760
rect 20444 18708 20496 18760
rect 22008 18708 22060 18760
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 8852 18572 8904 18624
rect 10876 18572 10928 18624
rect 11612 18572 11664 18624
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 13728 18572 13780 18624
rect 18420 18640 18472 18692
rect 19432 18640 19484 18692
rect 20904 18640 20956 18692
rect 22560 18683 22612 18692
rect 22560 18649 22569 18683
rect 22569 18649 22603 18683
rect 22603 18649 22612 18683
rect 22560 18640 22612 18649
rect 24400 18640 24452 18692
rect 18328 18572 18380 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 7748 18411 7800 18420
rect 7748 18377 7757 18411
rect 7757 18377 7791 18411
rect 7791 18377 7800 18411
rect 7748 18368 7800 18377
rect 9956 18368 10008 18420
rect 10416 18411 10468 18420
rect 10416 18377 10425 18411
rect 10425 18377 10459 18411
rect 10459 18377 10468 18411
rect 10416 18368 10468 18377
rect 12164 18368 12216 18420
rect 13360 18368 13412 18420
rect 18696 18368 18748 18420
rect 18880 18368 18932 18420
rect 19340 18368 19392 18420
rect 11152 18300 11204 18352
rect 11612 18300 11664 18352
rect 13544 18300 13596 18352
rect 4896 18028 4948 18080
rect 9864 18232 9916 18284
rect 10048 18232 10100 18284
rect 7564 18164 7616 18216
rect 8484 18164 8536 18216
rect 10692 18164 10744 18216
rect 11336 18232 11388 18284
rect 12164 18207 12216 18216
rect 12164 18173 12173 18207
rect 12173 18173 12207 18207
rect 12207 18173 12216 18207
rect 12164 18164 12216 18173
rect 12348 18207 12400 18216
rect 12348 18173 12357 18207
rect 12357 18173 12391 18207
rect 12391 18173 12400 18207
rect 12348 18164 12400 18173
rect 10784 18096 10836 18148
rect 14096 18300 14148 18352
rect 17500 18343 17552 18352
rect 17500 18309 17509 18343
rect 17509 18309 17543 18343
rect 17543 18309 17552 18343
rect 17500 18300 17552 18309
rect 19432 18300 19484 18352
rect 21088 18300 21140 18352
rect 13728 18232 13780 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 13820 18164 13872 18216
rect 15384 18164 15436 18216
rect 16028 18164 16080 18216
rect 16212 18164 16264 18216
rect 16488 18164 16540 18216
rect 20168 18164 20220 18216
rect 21088 18164 21140 18216
rect 23388 18164 23440 18216
rect 24768 18207 24820 18216
rect 24768 18173 24777 18207
rect 24777 18173 24811 18207
rect 24811 18173 24820 18207
rect 24768 18164 24820 18173
rect 8668 18028 8720 18080
rect 11244 18028 11296 18080
rect 22744 18096 22796 18148
rect 13728 18028 13780 18080
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 20168 18028 20220 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 7380 17824 7432 17876
rect 11980 17824 12032 17876
rect 12624 17824 12676 17876
rect 15844 17824 15896 17876
rect 19524 17824 19576 17876
rect 21272 17824 21324 17876
rect 6920 17688 6972 17740
rect 7840 17688 7892 17740
rect 8392 17688 8444 17740
rect 9404 17688 9456 17740
rect 4528 17620 4580 17672
rect 7288 17484 7340 17536
rect 9588 17620 9640 17672
rect 9956 17620 10008 17672
rect 10508 17663 10560 17672
rect 10508 17629 10517 17663
rect 10517 17629 10551 17663
rect 10551 17629 10560 17663
rect 10508 17620 10560 17629
rect 11704 17620 11756 17672
rect 12624 17620 12676 17672
rect 15568 17756 15620 17808
rect 16120 17756 16172 17808
rect 18880 17756 18932 17808
rect 14832 17731 14884 17740
rect 14832 17697 14841 17731
rect 14841 17697 14875 17731
rect 14875 17697 14884 17731
rect 14832 17688 14884 17697
rect 16304 17688 16356 17740
rect 11336 17595 11388 17604
rect 11336 17561 11345 17595
rect 11345 17561 11379 17595
rect 11379 17561 11388 17595
rect 11336 17552 11388 17561
rect 14740 17620 14792 17672
rect 17132 17688 17184 17740
rect 20904 17688 20956 17740
rect 22560 17824 22612 17876
rect 23848 17620 23900 17672
rect 24400 17824 24452 17876
rect 24860 17663 24912 17672
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 14096 17552 14148 17604
rect 8576 17484 8628 17536
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 9496 17527 9548 17536
rect 9496 17493 9505 17527
rect 9505 17493 9539 17527
rect 9539 17493 9548 17527
rect 9496 17484 9548 17493
rect 10140 17484 10192 17536
rect 12716 17484 12768 17536
rect 13544 17484 13596 17536
rect 14648 17527 14700 17536
rect 14648 17493 14657 17527
rect 14657 17493 14691 17527
rect 14691 17493 14700 17527
rect 14648 17484 14700 17493
rect 20168 17595 20220 17604
rect 20168 17561 20177 17595
rect 20177 17561 20211 17595
rect 20211 17561 20220 17595
rect 20168 17552 20220 17561
rect 15568 17484 15620 17536
rect 16580 17527 16632 17536
rect 16580 17493 16589 17527
rect 16589 17493 16623 17527
rect 16623 17493 16632 17527
rect 16580 17484 16632 17493
rect 19432 17484 19484 17536
rect 24216 17484 24268 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 4068 17280 4120 17332
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 6920 17076 6972 17128
rect 9496 17280 9548 17332
rect 10508 17280 10560 17332
rect 12532 17280 12584 17332
rect 9864 17212 9916 17264
rect 12072 17212 12124 17264
rect 13728 17280 13780 17332
rect 13820 17280 13872 17332
rect 16580 17280 16632 17332
rect 8760 17144 8812 17196
rect 9220 17144 9272 17196
rect 12532 17144 12584 17196
rect 10508 17119 10560 17128
rect 10508 17085 10517 17119
rect 10517 17085 10551 17119
rect 10551 17085 10560 17119
rect 10508 17076 10560 17085
rect 10968 17076 11020 17128
rect 11336 17076 11388 17128
rect 13360 17076 13412 17128
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 16672 17144 16724 17196
rect 20904 17280 20956 17332
rect 18420 17212 18472 17264
rect 19432 17212 19484 17264
rect 23848 17280 23900 17332
rect 22468 17212 22520 17264
rect 23756 17144 23808 17196
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 18604 17076 18656 17128
rect 19156 17076 19208 17128
rect 19340 17076 19392 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 24676 17119 24728 17128
rect 24676 17085 24685 17119
rect 24685 17085 24719 17119
rect 24719 17085 24728 17119
rect 24676 17076 24728 17085
rect 8300 17008 8352 17060
rect 8944 17008 8996 17060
rect 14648 17008 14700 17060
rect 7012 16940 7064 16992
rect 7472 16940 7524 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 22652 17008 22704 17060
rect 23296 17008 23348 17060
rect 19064 16940 19116 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6920 16736 6972 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 8300 16736 8352 16788
rect 8392 16668 8444 16720
rect 8576 16736 8628 16788
rect 10140 16736 10192 16788
rect 8760 16668 8812 16720
rect 9312 16668 9364 16720
rect 11612 16736 11664 16788
rect 23848 16779 23900 16788
rect 23848 16745 23857 16779
rect 23857 16745 23891 16779
rect 23891 16745 23900 16779
rect 23848 16736 23900 16745
rect 6644 16600 6696 16652
rect 8484 16600 8536 16652
rect 14280 16668 14332 16720
rect 19340 16711 19392 16720
rect 1492 16532 1544 16584
rect 7472 16532 7524 16584
rect 8300 16532 8352 16584
rect 9220 16532 9272 16584
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 12256 16643 12308 16652
rect 12256 16609 12265 16643
rect 12265 16609 12299 16643
rect 12299 16609 12308 16643
rect 12256 16600 12308 16609
rect 12624 16600 12676 16652
rect 15108 16600 15160 16652
rect 19340 16677 19349 16711
rect 19349 16677 19383 16711
rect 19383 16677 19392 16711
rect 19340 16668 19392 16677
rect 16028 16600 16080 16652
rect 20168 16600 20220 16652
rect 20904 16600 20956 16652
rect 22008 16643 22060 16652
rect 22008 16609 22017 16643
rect 22017 16609 22051 16643
rect 22051 16609 22060 16643
rect 22008 16600 22060 16609
rect 9588 16532 9640 16584
rect 10876 16575 10928 16584
rect 10876 16541 10885 16575
rect 10885 16541 10919 16575
rect 10919 16541 10928 16575
rect 10876 16532 10928 16541
rect 12716 16532 12768 16584
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 23388 16600 23440 16652
rect 1308 16464 1360 16516
rect 10324 16464 10376 16516
rect 12072 16464 12124 16516
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 9956 16396 10008 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 13820 16396 13872 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 15752 16396 15804 16448
rect 16948 16396 17000 16448
rect 22100 16464 22152 16516
rect 21180 16396 21232 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 7288 16192 7340 16244
rect 10508 16192 10560 16244
rect 11428 16192 11480 16244
rect 11520 16192 11572 16244
rect 12532 16192 12584 16244
rect 13360 16192 13412 16244
rect 13452 16192 13504 16244
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19892 16192 19944 16244
rect 20720 16192 20772 16244
rect 4068 16124 4120 16176
rect 7472 16124 7524 16176
rect 11796 16124 11848 16176
rect 13544 16124 13596 16176
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 17132 16167 17184 16176
rect 17132 16133 17141 16167
rect 17141 16133 17175 16167
rect 17175 16133 17184 16167
rect 17132 16124 17184 16133
rect 18420 16124 18472 16176
rect 19340 16124 19392 16176
rect 20996 16124 21048 16176
rect 21640 16124 21692 16176
rect 6644 16099 6696 16108
rect 6644 16065 6653 16099
rect 6653 16065 6687 16099
rect 6687 16065 6696 16099
rect 6644 16056 6696 16065
rect 8300 15988 8352 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 10416 16056 10468 16108
rect 12808 16056 12860 16108
rect 16580 16056 16632 16108
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22468 16056 22520 16108
rect 24124 16099 24176 16108
rect 24124 16065 24133 16099
rect 24133 16065 24167 16099
rect 24167 16065 24176 16099
rect 24124 16056 24176 16065
rect 1768 15852 1820 15904
rect 10232 15920 10284 15972
rect 11152 15988 11204 16040
rect 22284 15988 22336 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 23848 15920 23900 15972
rect 12348 15852 12400 15904
rect 14096 15852 14148 15904
rect 15752 15852 15804 15904
rect 17316 15852 17368 15904
rect 21824 15852 21876 15904
rect 21916 15852 21968 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 10232 15648 10284 15700
rect 11336 15512 11388 15564
rect 12440 15648 12492 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 19340 15580 19392 15632
rect 14372 15512 14424 15564
rect 17408 15512 17460 15564
rect 21180 15512 21232 15564
rect 13452 15487 13504 15496
rect 13452 15453 13461 15487
rect 13461 15453 13495 15487
rect 13495 15453 13504 15487
rect 13452 15444 13504 15453
rect 15292 15444 15344 15496
rect 16396 15444 16448 15496
rect 18696 15444 18748 15496
rect 19248 15444 19300 15496
rect 19892 15444 19944 15496
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 24216 15444 24268 15496
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 10416 15308 10468 15360
rect 10876 15308 10928 15360
rect 11796 15376 11848 15428
rect 16764 15376 16816 15428
rect 11704 15308 11756 15360
rect 12624 15308 12676 15360
rect 15660 15308 15712 15360
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 19616 15308 19668 15360
rect 21824 15419 21876 15428
rect 21824 15385 21833 15419
rect 21833 15385 21867 15419
rect 21867 15385 21876 15419
rect 21824 15376 21876 15385
rect 26056 15376 26108 15428
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 21548 15308 21600 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 8760 15104 8812 15156
rect 9404 15079 9456 15088
rect 9404 15045 9413 15079
rect 9413 15045 9447 15079
rect 9447 15045 9456 15079
rect 9404 15036 9456 15045
rect 12164 15104 12216 15156
rect 17316 15104 17368 15156
rect 18696 15104 18748 15156
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 22376 15104 22428 15156
rect 10876 14900 10928 14952
rect 9956 14764 10008 14816
rect 10508 14764 10560 14816
rect 11796 14764 11848 14816
rect 12532 15036 12584 15088
rect 13452 15079 13504 15088
rect 13452 15045 13461 15079
rect 13461 15045 13495 15079
rect 13495 15045 13504 15079
rect 13452 15036 13504 15045
rect 17040 15036 17092 15088
rect 17224 15079 17276 15088
rect 17224 15045 17233 15079
rect 17233 15045 17267 15079
rect 17267 15045 17276 15079
rect 17224 15036 17276 15045
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 13912 14900 13964 14952
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 15476 14968 15528 15020
rect 18604 14968 18656 15020
rect 16396 14900 16448 14952
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 23664 14968 23716 15020
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 16672 14832 16724 14884
rect 19524 14832 19576 14884
rect 19156 14764 19208 14816
rect 19800 14764 19852 14816
rect 19892 14764 19944 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10784 14560 10836 14612
rect 11336 14492 11388 14544
rect 11796 14492 11848 14544
rect 12808 14560 12860 14612
rect 17132 14603 17184 14612
rect 17132 14569 17141 14603
rect 17141 14569 17175 14603
rect 17175 14569 17184 14603
rect 17132 14560 17184 14569
rect 14556 14492 14608 14544
rect 16948 14492 17000 14544
rect 20812 14492 20864 14544
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 13452 14467 13504 14476
rect 12532 14424 12584 14433
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 14740 14424 14792 14476
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 16396 14424 16448 14476
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 18512 14356 18564 14408
rect 20076 14356 20128 14408
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 22284 14356 22336 14408
rect 23388 14560 23440 14612
rect 10232 14331 10284 14340
rect 10232 14297 10241 14331
rect 10241 14297 10275 14331
rect 10275 14297 10284 14331
rect 10232 14288 10284 14297
rect 10508 14288 10560 14340
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 15936 14288 15988 14340
rect 9864 14220 9916 14272
rect 10968 14220 11020 14272
rect 15568 14220 15620 14272
rect 16396 14220 16448 14272
rect 16488 14220 16540 14272
rect 21180 14288 21232 14340
rect 18420 14220 18472 14272
rect 18512 14220 18564 14272
rect 18972 14220 19024 14272
rect 19984 14263 20036 14272
rect 19984 14229 19993 14263
rect 19993 14229 20027 14263
rect 20027 14229 20036 14263
rect 19984 14220 20036 14229
rect 21824 14220 21876 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 9956 14016 10008 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 8760 13948 8812 14000
rect 11888 13948 11940 14000
rect 13544 14016 13596 14068
rect 18328 14016 18380 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 21088 14016 21140 14068
rect 23388 14016 23440 14068
rect 1308 13812 1360 13864
rect 8760 13812 8812 13864
rect 10232 13880 10284 13932
rect 10508 13880 10560 13932
rect 15292 13948 15344 14000
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 9496 13812 9548 13864
rect 10416 13812 10468 13864
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 18420 13880 18472 13932
rect 19984 13880 20036 13932
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 21088 13880 21140 13932
rect 12808 13812 12860 13864
rect 11796 13744 11848 13796
rect 9864 13676 9916 13728
rect 18972 13812 19024 13864
rect 20352 13812 20404 13864
rect 21732 13948 21784 14000
rect 22744 13948 22796 14000
rect 21456 13880 21508 13932
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 21364 13812 21416 13864
rect 23756 13812 23808 13864
rect 22192 13744 22244 13796
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 7104 13515 7156 13524
rect 7104 13481 7134 13515
rect 7134 13481 7156 13515
rect 7104 13472 7156 13481
rect 7564 13472 7616 13524
rect 8760 13472 8812 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 12808 13472 12860 13524
rect 8484 13336 8536 13388
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 8392 13268 8444 13320
rect 8760 13268 8812 13320
rect 5816 13132 5868 13184
rect 10232 13200 10284 13252
rect 10600 13200 10652 13252
rect 8760 13132 8812 13184
rect 11520 13132 11572 13184
rect 13268 13404 13320 13456
rect 12624 13336 12676 13388
rect 15384 13336 15436 13388
rect 15936 13472 15988 13524
rect 18880 13472 18932 13524
rect 19432 13447 19484 13456
rect 19432 13413 19441 13447
rect 19441 13413 19475 13447
rect 19475 13413 19484 13447
rect 19432 13404 19484 13413
rect 18512 13336 18564 13388
rect 20444 13472 20496 13524
rect 14464 13268 14516 13320
rect 16120 13268 16172 13320
rect 14372 13200 14424 13252
rect 14556 13200 14608 13252
rect 14832 13243 14884 13252
rect 14832 13209 14841 13243
rect 14841 13209 14875 13243
rect 14875 13209 14884 13243
rect 14832 13200 14884 13209
rect 16212 13200 16264 13252
rect 16488 13200 16540 13252
rect 21456 13268 21508 13320
rect 22652 13311 22704 13320
rect 22652 13277 22661 13311
rect 22661 13277 22695 13311
rect 22695 13277 22704 13311
rect 22652 13268 22704 13277
rect 20076 13200 20128 13252
rect 25136 13200 25188 13252
rect 17224 13132 17276 13184
rect 18880 13132 18932 13184
rect 19340 13132 19392 13184
rect 22284 13132 22336 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 6644 12928 6696 12980
rect 8392 12928 8444 12980
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 10600 12928 10652 12980
rect 6552 12792 6604 12844
rect 8668 12792 8720 12844
rect 8852 12792 8904 12844
rect 9680 12860 9732 12912
rect 9956 12860 10008 12912
rect 10232 12860 10284 12912
rect 11796 12928 11848 12980
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 14924 12971 14976 12980
rect 14924 12937 14933 12971
rect 14933 12937 14967 12971
rect 14967 12937 14976 12971
rect 14924 12928 14976 12937
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 17224 12971 17276 12980
rect 17224 12937 17233 12971
rect 17233 12937 17267 12971
rect 17267 12937 17276 12971
rect 17224 12928 17276 12937
rect 17316 12971 17368 12980
rect 17316 12937 17325 12971
rect 17325 12937 17359 12971
rect 17359 12937 17368 12971
rect 17316 12928 17368 12937
rect 11520 12903 11572 12912
rect 11520 12869 11529 12903
rect 11529 12869 11563 12903
rect 11563 12869 11572 12903
rect 11520 12860 11572 12869
rect 15200 12860 15252 12912
rect 19248 12928 19300 12980
rect 13636 12792 13688 12844
rect 13820 12792 13872 12844
rect 15936 12792 15988 12844
rect 8760 12767 8812 12776
rect 8760 12733 8769 12767
rect 8769 12733 8803 12767
rect 8803 12733 8812 12767
rect 8760 12724 8812 12733
rect 14832 12724 14884 12776
rect 18880 12792 18932 12844
rect 19524 12792 19576 12844
rect 18328 12724 18380 12776
rect 20904 12928 20956 12980
rect 21456 12971 21508 12980
rect 21456 12937 21465 12971
rect 21465 12937 21499 12971
rect 21499 12937 21508 12971
rect 21456 12928 21508 12937
rect 22284 12860 22336 12912
rect 22652 12860 22704 12912
rect 22100 12792 22152 12844
rect 23296 12792 23348 12844
rect 21824 12724 21876 12776
rect 22008 12767 22060 12776
rect 22008 12733 22017 12767
rect 22017 12733 22051 12767
rect 22051 12733 22060 12767
rect 22008 12724 22060 12733
rect 24768 12767 24820 12776
rect 24768 12733 24777 12767
rect 24777 12733 24811 12767
rect 24811 12733 24820 12767
rect 24768 12724 24820 12733
rect 14280 12656 14332 12708
rect 14648 12699 14700 12708
rect 14648 12665 14657 12699
rect 14657 12665 14691 12699
rect 14691 12665 14700 12699
rect 14648 12656 14700 12665
rect 16304 12588 16356 12640
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 20536 12588 20588 12640
rect 22560 12588 22612 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 2688 12384 2740 12436
rect 8668 12384 8720 12436
rect 10876 12384 10928 12436
rect 13820 12384 13872 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 9680 12248 9732 12300
rect 10968 12248 11020 12300
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 15936 12248 15988 12300
rect 13636 12180 13688 12232
rect 15844 12180 15896 12232
rect 17408 12384 17460 12436
rect 17500 12384 17552 12436
rect 19616 12316 19668 12368
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 19984 12248 20036 12300
rect 22836 12316 22888 12368
rect 21824 12248 21876 12300
rect 21916 12248 21968 12300
rect 18972 12180 19024 12232
rect 19156 12180 19208 12232
rect 22008 12180 22060 12232
rect 13452 12112 13504 12164
rect 16856 12112 16908 12164
rect 17316 12112 17368 12164
rect 13176 12044 13228 12096
rect 15384 12044 15436 12096
rect 16028 12044 16080 12096
rect 17408 12044 17460 12096
rect 19800 12112 19852 12164
rect 18972 12044 19024 12096
rect 19248 12044 19300 12096
rect 22744 12112 22796 12164
rect 24124 12044 24176 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 13452 11840 13504 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 15200 11840 15252 11892
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 10968 11704 11020 11756
rect 14740 11704 14792 11756
rect 18328 11840 18380 11892
rect 19248 11840 19300 11892
rect 18512 11815 18564 11824
rect 18512 11781 18521 11815
rect 18521 11781 18555 11815
rect 18555 11781 18564 11815
rect 18512 11772 18564 11781
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 22652 11840 22704 11892
rect 20812 11772 20864 11824
rect 22376 11704 22428 11756
rect 13176 11636 13228 11688
rect 21364 11636 21416 11688
rect 15752 11500 15804 11552
rect 16856 11500 16908 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 14372 11296 14424 11348
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 15936 11092 15988 11144
rect 19892 11092 19944 11144
rect 5908 11024 5960 11076
rect 10140 11024 10192 11076
rect 20628 11024 20680 11076
rect 20812 11067 20864 11076
rect 20812 11033 20821 11067
rect 20821 11033 20855 11067
rect 20855 11033 20864 11067
rect 20812 11024 20864 11033
rect 23940 11024 23992 11076
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 10048 10684 10100 10736
rect 16028 10684 16080 10736
rect 19616 10752 19668 10804
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 15752 10616 15804 10668
rect 19524 10616 19576 10668
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 23848 10616 23900 10668
rect 12808 10480 12860 10532
rect 15936 10480 15988 10532
rect 20812 10548 20864 10600
rect 24768 10591 24820 10600
rect 24768 10557 24777 10591
rect 24777 10557 24811 10591
rect 24811 10557 24820 10591
rect 24768 10548 24820 10557
rect 19984 10480 20036 10532
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 20628 10412 20680 10464
rect 23296 10412 23348 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 22468 10140 22520 10192
rect 18236 10072 18288 10124
rect 13360 10004 13412 10056
rect 19432 10004 19484 10056
rect 21272 10004 21324 10056
rect 16948 9979 17000 9988
rect 16948 9945 16957 9979
rect 16957 9945 16991 9979
rect 16991 9945 17000 9979
rect 16948 9936 17000 9945
rect 24952 10004 25004 10056
rect 18788 9868 18840 9920
rect 22744 9936 22796 9988
rect 24032 9868 24084 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 16396 9596 16448 9648
rect 17776 9596 17828 9648
rect 18696 9596 18748 9648
rect 21548 9596 21600 9648
rect 18420 9528 18472 9580
rect 22836 9528 22888 9580
rect 4252 9460 4304 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 17592 9392 17644 9444
rect 17684 9324 17736 9376
rect 22284 9324 22336 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 4068 9120 4120 9172
rect 5540 9120 5592 9172
rect 22652 9052 22704 9104
rect 22560 8984 22612 9036
rect 20628 8916 20680 8968
rect 23388 8916 23440 8968
rect 22836 8780 22888 8832
rect 23480 8780 23532 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 19064 8508 19116 8560
rect 21640 8508 21692 8560
rect 10048 8372 10100 8424
rect 13912 8372 13964 8424
rect 22008 8372 22060 8424
rect 21272 8304 21324 8356
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 22560 8415 22612 8424
rect 22560 8381 22569 8415
rect 22569 8381 22603 8415
rect 22603 8381 22612 8415
rect 22560 8372 22612 8381
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 24860 8304 24912 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 6828 8032 6880 8084
rect 22376 8032 22428 8084
rect 6184 7896 6236 7948
rect 6644 7896 6696 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 19800 7828 19852 7880
rect 20536 7828 20588 7880
rect 23480 7828 23532 7880
rect 25044 7828 25096 7880
rect 4344 7803 4396 7812
rect 4344 7769 4353 7803
rect 4353 7769 4387 7803
rect 4387 7769 4396 7803
rect 4344 7760 4396 7769
rect 20812 7692 20864 7744
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 17316 7420 17368 7472
rect 20904 7352 20956 7404
rect 22008 7352 22060 7404
rect 23296 7352 23348 7404
rect 21640 7284 21692 7336
rect 22284 7284 22336 7336
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 20628 7216 20680 7268
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 22376 6876 22428 6928
rect 22744 6876 22796 6928
rect 5816 6808 5868 6860
rect 10692 6808 10744 6860
rect 4068 6740 4120 6792
rect 6368 6740 6420 6792
rect 16396 6740 16448 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 22836 6783 22888 6792
rect 22836 6749 22845 6783
rect 22845 6749 22879 6783
rect 22879 6749 22888 6783
rect 22836 6740 22888 6749
rect 24124 6740 24176 6792
rect 22008 6715 22060 6724
rect 22008 6681 22017 6715
rect 22017 6681 22051 6715
rect 22051 6681 22060 6715
rect 22008 6672 22060 6681
rect 24952 6672 25004 6724
rect 18512 6604 18564 6656
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 4344 6400 4396 6452
rect 11612 6400 11664 6452
rect 2872 6264 2924 6316
rect 21088 6264 21140 6316
rect 21364 6264 21416 6316
rect 22192 6264 22244 6316
rect 20812 6196 20864 6248
rect 21732 6196 21784 6248
rect 21916 6196 21968 6248
rect 24584 6239 24636 6248
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 20904 5856 20956 5908
rect 20444 5720 20496 5772
rect 21548 5720 21600 5772
rect 7104 5652 7156 5704
rect 11980 5652 12032 5704
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 20352 5652 20404 5704
rect 20628 5652 20680 5704
rect 22468 5652 22520 5704
rect 21088 5584 21140 5636
rect 3424 5516 3476 5568
rect 4712 5516 4764 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 2872 5312 2924 5364
rect 19708 5244 19760 5296
rect 1768 5219 1820 5228
rect 1768 5185 1777 5219
rect 1777 5185 1811 5219
rect 1811 5185 1820 5219
rect 1768 5176 1820 5185
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 21824 5176 21876 5228
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 19616 5108 19668 5160
rect 22468 5151 22520 5160
rect 22468 5117 22477 5151
rect 22477 5117 22511 5151
rect 22511 5117 22520 5151
rect 22468 5108 22520 5117
rect 24768 5151 24820 5160
rect 24768 5117 24777 5151
rect 24777 5117 24811 5151
rect 24811 5117 24820 5151
rect 24768 5108 24820 5117
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 17776 4768 17828 4820
rect 4896 4700 4948 4752
rect 24860 4743 24912 4752
rect 24860 4709 24869 4743
rect 24869 4709 24903 4743
rect 24903 4709 24912 4743
rect 24860 4700 24912 4709
rect 11796 4632 11848 4684
rect 12624 4632 12676 4684
rect 19892 4675 19944 4684
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 20720 4632 20772 4684
rect 18512 4564 18564 4616
rect 18604 4564 18656 4616
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 22744 4564 22796 4616
rect 2044 4496 2096 4548
rect 20628 4496 20680 4548
rect 23296 4496 23348 4548
rect 12624 4428 12676 4480
rect 14188 4428 14240 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 1768 4224 1820 4276
rect 9312 4224 9364 4276
rect 10324 4224 10376 4276
rect 13544 4224 13596 4276
rect 2228 4088 2280 4140
rect 2412 4088 2464 4140
rect 25136 4199 25188 4208
rect 25136 4165 25145 4199
rect 25145 4165 25179 4199
rect 25179 4165 25188 4199
rect 25136 4156 25188 4165
rect 4068 4020 4120 4072
rect 6000 4020 6052 4072
rect 11612 4020 11664 4072
rect 3424 3952 3476 4004
rect 9036 3952 9088 4004
rect 6092 3884 6144 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 10324 3884 10376 3936
rect 13452 4020 13504 4072
rect 12164 3952 12216 4004
rect 16672 4088 16724 4140
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 24676 4088 24728 4140
rect 16396 4020 16448 4072
rect 17500 4020 17552 4072
rect 20076 4020 20128 4072
rect 19708 3952 19760 4004
rect 22100 3952 22152 4004
rect 15936 3884 15988 3936
rect 22192 3884 22244 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 4252 3680 4304 3732
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 9312 3723 9364 3732
rect 9312 3689 9321 3723
rect 9321 3689 9355 3723
rect 9355 3689 9364 3723
rect 9312 3680 9364 3689
rect 10048 3723 10100 3732
rect 10048 3689 10057 3723
rect 10057 3689 10091 3723
rect 10091 3689 10100 3723
rect 10048 3680 10100 3689
rect 18788 3680 18840 3732
rect 3516 3544 3568 3596
rect 12164 3612 12216 3664
rect 8944 3544 8996 3596
rect 15108 3612 15160 3664
rect 20812 3612 20864 3664
rect 24952 3612 25004 3664
rect 12716 3544 12768 3596
rect 14924 3544 14976 3596
rect 16028 3544 16080 3596
rect 17868 3544 17920 3596
rect 2872 3476 2924 3528
rect 1676 3408 1728 3460
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 7840 3476 7892 3528
rect 9496 3476 9548 3528
rect 9772 3476 9824 3528
rect 10876 3476 10928 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 15568 3476 15620 3528
rect 16304 3476 16356 3528
rect 19340 3476 19392 3528
rect 21180 3476 21232 3528
rect 8300 3408 8352 3460
rect 18972 3408 19024 3460
rect 24124 3408 24176 3460
rect 4988 3340 5040 3392
rect 6828 3340 6880 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 11244 3340 11296 3392
rect 11704 3340 11756 3392
rect 22008 3340 22060 3392
rect 22836 3340 22888 3392
rect 24584 3340 24636 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6552 3136 6604 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7196 3136 7248 3188
rect 8852 3136 8904 3188
rect 11336 3136 11388 3188
rect 25044 3136 25096 3188
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 5356 3000 5408 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8208 3000 8260 3052
rect 8668 3000 8720 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9588 3000 9640 3052
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 13636 3068 13688 3120
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 3424 2932 3476 2984
rect 10416 2932 10468 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 14188 2932 14240 2984
rect 15660 2932 15712 2984
rect 17132 2864 17184 2916
rect 20628 2932 20680 2984
rect 23388 2932 23440 2984
rect 19708 2864 19760 2916
rect 20720 2864 20772 2916
rect 20812 2864 20864 2916
rect 22468 2864 22520 2916
rect 4252 2796 4304 2848
rect 16764 2796 16816 2848
rect 17960 2796 18012 2848
rect 18604 2796 18656 2848
rect 19892 2796 19944 2848
rect 21732 2796 21784 2848
rect 22652 2796 22704 2848
rect 24124 2839 24176 2848
rect 24124 2805 24133 2839
rect 24133 2805 24167 2839
rect 24167 2805 24176 2839
rect 24124 2796 24176 2805
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 1584 2592 1636 2644
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 9864 2592 9916 2644
rect 15384 2592 15436 2644
rect 18696 2592 18748 2644
rect 25320 2592 25372 2644
rect 11796 2524 11848 2576
rect 17592 2524 17644 2576
rect 1308 2388 1360 2440
rect 3884 2388 3936 2440
rect 4252 2388 4304 2440
rect 4620 2388 4672 2440
rect 11704 2456 11756 2508
rect 6000 2388 6052 2440
rect 7196 2388 7248 2440
rect 7564 2388 7616 2440
rect 10140 2388 10192 2440
rect 11980 2456 12032 2508
rect 14556 2456 14608 2508
rect 15292 2456 15344 2508
rect 17960 2456 18012 2508
rect 5724 2320 5776 2372
rect 12808 2388 12860 2440
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 12348 2320 12400 2372
rect 13820 2320 13872 2372
rect 18328 2320 18380 2372
rect 24860 2456 24912 2508
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1490 56200 1546 57000
rect 1858 56200 1914 57000
rect 2226 56200 2282 57000
rect 2594 56200 2650 57000
rect 2962 56200 3018 57000
rect 3330 56200 3386 57000
rect 3698 56200 3754 57000
rect 4066 56200 4122 57000
rect 4434 56200 4490 57000
rect 4802 56200 4858 57000
rect 5170 56200 5226 57000
rect 5538 56200 5594 57000
rect 5906 56200 5962 57000
rect 6274 56200 6330 57000
rect 6642 56200 6698 57000
rect 7010 56200 7066 57000
rect 7378 56200 7434 57000
rect 7746 56200 7802 57000
rect 7852 56222 8064 56250
rect 1306 53000 1362 53009
rect 1306 52935 1362 52944
rect 1320 52630 1348 52935
rect 1308 52624 1360 52630
rect 1308 52566 1360 52572
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1320 50386 1348 50487
rect 1308 50380 1360 50386
rect 1308 50322 1360 50328
rect 1504 49298 1532 56200
rect 1676 53100 1728 53106
rect 1676 53042 1728 53048
rect 1688 52154 1716 53042
rect 1872 52970 1900 56200
rect 1860 52964 1912 52970
rect 1860 52906 1912 52912
rect 1768 52896 1820 52902
rect 1768 52838 1820 52844
rect 1676 52148 1728 52154
rect 1676 52090 1728 52096
rect 1780 50930 1808 52838
rect 2240 52698 2268 56200
rect 2320 54188 2372 54194
rect 2320 54130 2372 54136
rect 2228 52692 2280 52698
rect 2228 52634 2280 52640
rect 2332 50998 2360 54130
rect 2608 52986 2636 56200
rect 2976 55214 3004 56200
rect 2884 55186 3004 55214
rect 2608 52958 2820 52986
rect 2320 50992 2372 50998
rect 2320 50934 2372 50940
rect 1768 50924 1820 50930
rect 1768 50866 1820 50872
rect 2792 50862 2820 52958
rect 2884 51474 2912 55186
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 3344 51950 3372 56200
rect 3516 52964 3568 52970
rect 3516 52906 3568 52912
rect 3424 52692 3476 52698
rect 3424 52634 3476 52640
rect 3332 51944 3384 51950
rect 3332 51886 3384 51892
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 2872 51468 2924 51474
rect 2872 51410 2924 51416
rect 2780 50856 2832 50862
rect 2780 50798 2832 50804
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 3436 50386 3464 52634
rect 3424 50380 3476 50386
rect 3424 50322 3476 50328
rect 3528 49910 3556 52906
rect 3712 52562 3740 56200
rect 3974 55448 4030 55457
rect 3974 55383 4030 55392
rect 3988 54330 4016 55383
rect 3976 54324 4028 54330
rect 3976 54266 4028 54272
rect 3792 53984 3844 53990
rect 3792 53926 3844 53932
rect 3804 52630 3832 53926
rect 3988 53582 4016 54266
rect 3976 53576 4028 53582
rect 3976 53518 4028 53524
rect 4080 53258 4108 56200
rect 4080 53230 4384 53258
rect 4160 53100 4212 53106
rect 4160 53042 4212 53048
rect 3792 52624 3844 52630
rect 3792 52566 3844 52572
rect 3700 52556 3752 52562
rect 3700 52498 3752 52504
rect 4172 52154 4200 53042
rect 4160 52148 4212 52154
rect 4160 52090 4212 52096
rect 3976 51400 4028 51406
rect 3976 51342 4028 51348
rect 3988 51066 4016 51342
rect 4252 51264 4304 51270
rect 4252 51206 4304 51212
rect 3976 51060 4028 51066
rect 3976 51002 4028 51008
rect 4160 50788 4212 50794
rect 4160 50730 4212 50736
rect 3516 49904 3568 49910
rect 3516 49846 3568 49852
rect 1952 49836 2004 49842
rect 1952 49778 2004 49784
rect 1492 49292 1544 49298
rect 1492 49234 1544 49240
rect 1306 48104 1362 48113
rect 1306 48039 1308 48048
rect 1360 48039 1362 48048
rect 1308 48010 1360 48016
rect 1308 45960 1360 45966
rect 1308 45902 1360 45908
rect 1320 45665 1348 45902
rect 1306 45656 1362 45665
rect 1306 45591 1308 45600
rect 1360 45591 1362 45600
rect 1308 45562 1360 45568
rect 1308 43308 1360 43314
rect 1308 43250 1360 43256
rect 1320 43217 1348 43250
rect 1306 43208 1362 43217
rect 1306 43143 1362 43152
rect 1964 41274 1992 49778
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 4068 48000 4120 48006
rect 4068 47942 4120 47948
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 3976 43172 4028 43178
rect 3976 43114 4028 43120
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 1952 41268 2004 41274
rect 1952 41210 2004 41216
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 1320 40769 1348 41074
rect 1676 40928 1728 40934
rect 1676 40870 1728 40876
rect 1306 40760 1362 40769
rect 1306 40695 1362 40704
rect 1308 38344 1360 38350
rect 1306 38312 1308 38321
rect 1360 38312 1362 38321
rect 1306 38247 1362 38256
rect 1584 38208 1636 38214
rect 1584 38150 1636 38156
rect 1308 33516 1360 33522
rect 1308 33458 1360 33464
rect 1320 33425 1348 33458
rect 1306 33416 1362 33425
rect 1306 33351 1362 33360
rect 1308 31272 1360 31278
rect 1308 31214 1360 31220
rect 1320 30977 1348 31214
rect 1306 30968 1362 30977
rect 1306 30903 1362 30912
rect 1596 29714 1624 38150
rect 1688 30802 1716 40870
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 1780 35873 1808 36110
rect 1766 35864 1822 35873
rect 1766 35799 1822 35808
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 3516 33312 3568 33318
rect 3516 33254 3568 33260
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1676 30796 1728 30802
rect 1676 30738 1728 30744
rect 1584 29708 1636 29714
rect 1584 29650 1636 29656
rect 1308 28620 1360 28626
rect 1308 28562 1360 28568
rect 1320 28529 1348 28562
rect 1768 28552 1820 28558
rect 1306 28520 1362 28529
rect 1768 28494 1820 28500
rect 1306 28455 1362 28464
rect 1780 26042 1808 28494
rect 1964 28218 1992 31282
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 1952 28212 2004 28218
rect 1952 28154 2004 28160
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 1768 26036 1820 26042
rect 1768 25978 1820 25984
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1768 23724 1820 23730
rect 1768 23666 1820 23672
rect 1308 23656 1360 23662
rect 1306 23624 1308 23633
rect 1360 23624 1362 23633
rect 1306 23559 1362 23568
rect 1780 22778 1808 23666
rect 1768 22772 1820 22778
rect 1768 22714 1820 22720
rect 1872 21554 1900 24006
rect 2056 23322 2084 26318
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2792 26081 2820 26250
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2780 25832 2832 25838
rect 2780 25774 2832 25780
rect 2792 24206 2820 25774
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2884 23322 2912 25842
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3344 24410 3372 26930
rect 3436 25770 3464 28018
rect 3528 26994 3556 33254
rect 3988 31754 4016 43114
rect 4080 39030 4108 47942
rect 4172 42362 4200 50730
rect 4264 49910 4292 51206
rect 4356 50862 4384 53230
rect 4448 53174 4476 56200
rect 4816 55214 4844 56200
rect 4816 55186 4936 55214
rect 4620 53440 4672 53446
rect 4620 53382 4672 53388
rect 4436 53168 4488 53174
rect 4436 53110 4488 53116
rect 4632 52086 4660 53382
rect 4712 53100 4764 53106
rect 4712 53042 4764 53048
rect 4620 52080 4672 52086
rect 4620 52022 4672 52028
rect 4344 50856 4396 50862
rect 4344 50798 4396 50804
rect 4252 49904 4304 49910
rect 4252 49846 4304 49852
rect 4724 45014 4752 53042
rect 4908 51950 4936 55186
rect 5184 53242 5212 56200
rect 5356 54188 5408 54194
rect 5356 54130 5408 54136
rect 5172 53236 5224 53242
rect 5172 53178 5224 53184
rect 5172 52488 5224 52494
rect 5172 52430 5224 52436
rect 4896 51944 4948 51950
rect 4896 51886 4948 51892
rect 4896 51808 4948 51814
rect 4896 51750 4948 51756
rect 4712 45008 4764 45014
rect 4712 44950 4764 44956
rect 4908 42770 4936 51750
rect 5080 50176 5132 50182
rect 5080 50118 5132 50124
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 4804 42628 4856 42634
rect 4804 42570 4856 42576
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4068 39024 4120 39030
rect 4068 38966 4120 38972
rect 4160 36032 4212 36038
rect 4160 35974 4212 35980
rect 3988 31726 4108 31754
rect 3792 30660 3844 30666
rect 3792 30602 3844 30608
rect 3804 28218 3832 30602
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3792 28212 3844 28218
rect 3792 28154 3844 28160
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3516 25968 3568 25974
rect 3516 25910 3568 25916
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 3344 23186 3372 24346
rect 3528 24206 3556 25910
rect 3620 25838 3648 28018
rect 3896 27130 3924 29514
rect 3976 28484 4028 28490
rect 3976 28426 4028 28432
rect 3884 27124 3936 27130
rect 3884 27066 3936 27072
rect 3700 26852 3752 26858
rect 3700 26794 3752 26800
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 2872 23180 2924 23186
rect 2872 23122 2924 23128
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 2884 23066 2912 23122
rect 2792 23038 2912 23066
rect 1860 21548 1912 21554
rect 1860 21490 1912 21496
rect 1308 21480 1360 21486
rect 1308 21422 1360 21428
rect 1320 21185 1348 21422
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 2792 20806 2820 23038
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2884 21146 2912 22578
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18737 1348 18770
rect 1306 18728 1362 18737
rect 1306 18663 1362 18672
rect 1504 16590 1532 19450
rect 1780 18766 1808 20742
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 13938 1808 15846
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1308 13864 1360 13870
rect 1306 13832 1308 13841
rect 1360 13832 1362 13841
rect 1306 13767 1362 13776
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 1950 8392 2006 8401
rect 1950 8327 2006 8336
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1780 4282 1808 5170
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1964 3738 1992 8327
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1596 2650 1624 2994
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1320 1601 1348 2382
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 1688 800 1716 3402
rect 2056 800 2084 4490
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2240 3194 2268 4082
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2424 800 2452 4082
rect 2700 3738 2728 12378
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2884 5370 2912 6258
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2884 3194 2912 3470
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2884 2774 2912 3130
rect 2792 2746 2912 2774
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 2792 800 2820 2746
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3344 2650 3372 22918
rect 3712 22094 3740 26794
rect 3988 25158 4016 28426
rect 4080 26586 4108 31726
rect 4172 28626 4200 35974
rect 4264 29850 4292 42162
rect 4620 41132 4672 41138
rect 4620 41074 4672 41080
rect 4632 32570 4660 41074
rect 4816 34474 4844 42570
rect 5092 42362 5120 50118
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 5184 41818 5212 52430
rect 5368 51074 5396 54130
rect 5552 53718 5580 56200
rect 5920 54126 5948 56200
rect 5908 54120 5960 54126
rect 5908 54062 5960 54068
rect 5540 53712 5592 53718
rect 5540 53654 5592 53660
rect 5540 53576 5592 53582
rect 5540 53518 5592 53524
rect 5276 51046 5396 51074
rect 5276 49722 5304 51046
rect 5448 50924 5500 50930
rect 5448 50866 5500 50872
rect 5276 49694 5396 49722
rect 5264 44396 5316 44402
rect 5264 44338 5316 44344
rect 5172 41812 5224 41818
rect 5172 41754 5224 41760
rect 5276 38010 5304 44338
rect 5368 43382 5396 49694
rect 5356 43376 5408 43382
rect 5356 43318 5408 43324
rect 5460 42362 5488 50866
rect 5552 50522 5580 53518
rect 6184 53236 6236 53242
rect 6184 53178 6236 53184
rect 6000 52488 6052 52494
rect 6000 52430 6052 52436
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 5816 50312 5868 50318
rect 5816 50254 5868 50260
rect 5828 44538 5856 50254
rect 6012 46170 6040 52430
rect 6196 51338 6224 53178
rect 6288 53174 6316 56200
rect 6276 53168 6328 53174
rect 6276 53110 6328 53116
rect 6656 52494 6684 56200
rect 6644 52488 6696 52494
rect 6644 52430 6696 52436
rect 7024 51474 7052 56200
rect 7392 53650 7420 56200
rect 7380 53644 7432 53650
rect 7380 53586 7432 53592
rect 7564 53508 7616 53514
rect 7564 53450 7616 53456
rect 7288 53100 7340 53106
rect 7288 53042 7340 53048
rect 7196 52012 7248 52018
rect 7196 51954 7248 51960
rect 6920 51468 6972 51474
rect 6920 51410 6972 51416
rect 7012 51468 7064 51474
rect 7012 51410 7064 51416
rect 6736 51400 6788 51406
rect 6736 51342 6788 51348
rect 6184 51332 6236 51338
rect 6184 51274 6236 51280
rect 6000 46164 6052 46170
rect 6000 46106 6052 46112
rect 6644 44736 6696 44742
rect 6644 44678 6696 44684
rect 5816 44532 5868 44538
rect 5816 44474 5868 44480
rect 6656 44418 6684 44678
rect 6748 44538 6776 51342
rect 6932 51066 6960 51410
rect 7104 51400 7156 51406
rect 7104 51342 7156 51348
rect 7012 51332 7064 51338
rect 7012 51274 7064 51280
rect 6920 51060 6972 51066
rect 6920 51002 6972 51008
rect 6920 45892 6972 45898
rect 6920 45834 6972 45840
rect 6736 44532 6788 44538
rect 6736 44474 6788 44480
rect 6656 44402 6776 44418
rect 6656 44396 6788 44402
rect 6656 44390 6736 44396
rect 6736 44338 6788 44344
rect 5448 42356 5500 42362
rect 5448 42298 5500 42304
rect 6368 42016 6420 42022
rect 6368 41958 6420 41964
rect 6184 41676 6236 41682
rect 6184 41618 6236 41624
rect 5908 41472 5960 41478
rect 5908 41414 5960 41420
rect 5816 39296 5868 39302
rect 5816 39238 5868 39244
rect 5264 38004 5316 38010
rect 5264 37946 5316 37952
rect 4988 37868 5040 37874
rect 4988 37810 5040 37816
rect 4804 34468 4856 34474
rect 4804 34410 4856 34416
rect 5000 32570 5028 37810
rect 5828 37806 5856 39238
rect 5816 37800 5868 37806
rect 5816 37742 5868 37748
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5448 36712 5500 36718
rect 5448 36654 5500 36660
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 32570 5396 33390
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 4896 32496 4948 32502
rect 4896 32438 4948 32444
rect 4252 29844 4304 29850
rect 4252 29786 4304 29792
rect 4160 28620 4212 28626
rect 4160 28562 4212 28568
rect 4344 26920 4396 26926
rect 4344 26862 4396 26868
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4080 25974 4108 26522
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3988 24206 4016 24550
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3988 23662 4016 24142
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3792 23044 3844 23050
rect 3792 22986 3844 22992
rect 3528 22066 3740 22094
rect 3528 11257 3556 22066
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 19378 3648 21422
rect 3804 21418 3832 22986
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 3988 21026 4016 23054
rect 4080 21486 4108 25230
rect 4264 24954 4292 25638
rect 4252 24948 4304 24954
rect 4252 24890 4304 24896
rect 4264 24274 4292 24890
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4356 23118 4384 26862
rect 4436 24404 4488 24410
rect 4436 24346 4488 24352
rect 4344 23112 4396 23118
rect 4344 23054 4396 23060
rect 4448 22930 4476 24346
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4356 22902 4476 22930
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3988 20998 4108 21026
rect 4080 20942 4108 20998
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 4080 17338 4108 20878
rect 4172 19514 4200 21490
rect 4264 20942 4292 22374
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4356 20534 4384 22902
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 16182 4108 17274
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4448 12434 4476 22442
rect 4540 21894 4568 24074
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4540 21554 4568 21830
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4540 17678 4568 21490
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4172 12406 4476 12434
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 8945 4108 9114
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4080 6497 4108 6734
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 4010 3464 5510
rect 4068 4072 4120 4078
rect 4066 4040 4068 4049
rect 4120 4040 4122 4049
rect 3424 4004 3476 4010
rect 4066 3975 4122 3984
rect 3424 3946 3476 3952
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3160 870 3280 898
rect 3160 800 3188 870
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3252 762 3280 870
rect 3436 762 3464 2926
rect 3528 800 3556 3538
rect 4172 2650 4200 12406
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4264 3738 4292 9454
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 6458 4384 7754
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4724 5574 4752 20742
rect 4908 18086 4936 32438
rect 5460 32366 5488 36654
rect 5552 35834 5580 36858
rect 5828 36718 5856 37742
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5552 35154 5580 35770
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5552 34066 5580 35090
rect 5632 34468 5684 34474
rect 5632 34410 5684 34416
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5552 32978 5580 34002
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5552 32502 5580 32914
rect 5540 32496 5592 32502
rect 5540 32438 5592 32444
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5644 31278 5672 34410
rect 5828 34066 5856 35566
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5632 31272 5684 31278
rect 5632 31214 5684 31220
rect 5920 31210 5948 41414
rect 6196 41274 6224 41618
rect 6184 41268 6236 41274
rect 6184 41210 6236 41216
rect 6196 40526 6224 41210
rect 6184 40520 6236 40526
rect 6184 40462 6236 40468
rect 6196 39506 6224 40462
rect 6184 39500 6236 39506
rect 6184 39442 6236 39448
rect 6092 36848 6144 36854
rect 6092 36790 6144 36796
rect 6000 36712 6052 36718
rect 6000 36654 6052 36660
rect 6012 35834 6040 36654
rect 6104 36582 6132 36790
rect 6092 36576 6144 36582
rect 6092 36518 6144 36524
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 6012 34678 6040 35770
rect 6104 35698 6132 36518
rect 6092 35692 6144 35698
rect 6092 35634 6144 35640
rect 6092 35148 6144 35154
rect 6092 35090 6144 35096
rect 6000 34672 6052 34678
rect 6000 34614 6052 34620
rect 6104 34610 6132 35090
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 6184 32496 6236 32502
rect 6184 32438 6236 32444
rect 6196 31890 6224 32438
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 5908 31204 5960 31210
rect 5908 31146 5960 31152
rect 5908 30660 5960 30666
rect 5908 30602 5960 30608
rect 5632 28620 5684 28626
rect 5552 28580 5632 28608
rect 5552 28422 5580 28580
rect 5632 28562 5684 28568
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 5092 20058 5120 22986
rect 5460 22982 5488 25842
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4908 4758 4936 18022
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4264 2446 4292 2790
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 3896 800 3924 2382
rect 4264 800 4292 2382
rect 4632 800 4660 2382
rect 5000 800 5028 3334
rect 5184 3194 5212 18906
rect 5552 9178 5580 28358
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5828 24614 5856 24754
rect 5816 24608 5868 24614
rect 5816 24550 5868 24556
rect 5828 24138 5856 24550
rect 5816 24132 5868 24138
rect 5816 24074 5868 24080
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 23186 5764 23462
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5736 20398 5764 23122
rect 5920 22710 5948 30602
rect 6380 30326 6408 41958
rect 6748 41414 6776 44338
rect 6656 41386 6776 41414
rect 6932 41414 6960 45834
rect 7024 43926 7052 51274
rect 7116 51074 7144 51342
rect 7208 51338 7236 51954
rect 7196 51332 7248 51338
rect 7196 51274 7248 51280
rect 7116 51046 7236 51074
rect 7104 44736 7156 44742
rect 7104 44678 7156 44684
rect 7116 44402 7144 44678
rect 7104 44396 7156 44402
rect 7104 44338 7156 44344
rect 7012 43920 7064 43926
rect 7012 43862 7064 43868
rect 6932 41386 7052 41414
rect 6552 40588 6604 40594
rect 6552 40530 6604 40536
rect 6564 39642 6592 40530
rect 6552 39636 6604 39642
rect 6552 39578 6604 39584
rect 6552 38208 6604 38214
rect 6552 38150 6604 38156
rect 6564 37806 6592 38150
rect 6552 37800 6604 37806
rect 6552 37742 6604 37748
rect 6564 37262 6592 37742
rect 6656 37670 6684 41386
rect 7024 39386 7052 41386
rect 7116 39846 7144 44338
rect 7208 44334 7236 51046
rect 7300 48142 7328 53042
rect 7380 52488 7432 52494
rect 7380 52430 7432 52436
rect 7288 48136 7340 48142
rect 7288 48078 7340 48084
rect 7392 45082 7420 52430
rect 7472 50856 7524 50862
rect 7472 50798 7524 50804
rect 7484 46714 7512 50798
rect 7472 46708 7524 46714
rect 7472 46650 7524 46656
rect 7472 45960 7524 45966
rect 7472 45902 7524 45908
rect 7380 45076 7432 45082
rect 7380 45018 7432 45024
rect 7484 44554 7512 45902
rect 7392 44526 7512 44554
rect 7196 44328 7248 44334
rect 7196 44270 7248 44276
rect 7196 42220 7248 42226
rect 7196 42162 7248 42168
rect 7208 42022 7236 42162
rect 7196 42016 7248 42022
rect 7196 41958 7248 41964
rect 7104 39840 7156 39846
rect 7104 39782 7156 39788
rect 7024 39358 7144 39386
rect 7012 39296 7064 39302
rect 7012 39238 7064 39244
rect 6736 38888 6788 38894
rect 6736 38830 6788 38836
rect 6644 37664 6696 37670
rect 6644 37606 6696 37612
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6564 36922 6592 37198
rect 6552 36916 6604 36922
rect 6552 36858 6604 36864
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6184 25832 6236 25838
rect 6184 25774 6236 25780
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 23866 6040 24686
rect 6196 24410 6224 25774
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6380 24342 6408 29514
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6564 28626 6592 29038
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 6564 27538 6592 28562
rect 6552 27532 6604 27538
rect 6552 27474 6604 27480
rect 6564 26994 6592 27474
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6564 26466 6592 26930
rect 6472 26450 6592 26466
rect 6460 26444 6592 26450
rect 6512 26438 6592 26444
rect 6460 26386 6512 26392
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 5920 22094 5948 22646
rect 6012 22574 6040 23802
rect 6000 22568 6052 22574
rect 6000 22510 6052 22516
rect 5920 22066 6040 22094
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5736 20058 5764 20334
rect 5828 20262 5856 21286
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5828 13190 5856 20198
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5368 800 5396 2994
rect 5736 2378 5764 2994
rect 5828 2774 5856 6802
rect 5920 3194 5948 11018
rect 6012 4078 6040 22066
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6196 7954 6224 18770
rect 6288 17882 6316 19314
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6380 6798 6408 24278
rect 6472 23186 6500 26386
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6564 23866 6592 24074
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6656 22506 6684 25094
rect 6644 22500 6696 22506
rect 6644 22442 6696 22448
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6564 20466 6592 20538
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 20058 6592 20402
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6564 17134 6592 19314
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16640 6592 17070
rect 6644 16652 6696 16658
rect 6564 16612 6644 16640
rect 6644 16594 6696 16600
rect 6656 16114 6684 16594
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 9450 6592 12786
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6656 7954 6684 12922
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3534 6132 3878
rect 6748 3738 6776 38830
rect 7024 38758 7052 39238
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 6920 38412 6972 38418
rect 6920 38354 6972 38360
rect 6932 37942 6960 38354
rect 7116 38214 7144 39358
rect 7104 38208 7156 38214
rect 7104 38150 7156 38156
rect 6920 37936 6972 37942
rect 6920 37878 6972 37884
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 7116 31890 7144 34682
rect 7208 34134 7236 41958
rect 7288 40384 7340 40390
rect 7288 40326 7340 40332
rect 7300 38350 7328 40326
rect 7392 40186 7420 44526
rect 7576 44470 7604 53450
rect 7760 52562 7788 56200
rect 7852 54262 7880 56222
rect 8036 56114 8064 56222
rect 8114 56200 8170 57000
rect 8482 56200 8538 57000
rect 8850 56200 8906 57000
rect 9218 56200 9274 57000
rect 9586 56200 9642 57000
rect 9954 56200 10010 57000
rect 10322 56200 10378 57000
rect 10690 56200 10746 57000
rect 11058 56200 11114 57000
rect 11426 56200 11482 57000
rect 11794 56200 11850 57000
rect 12162 56200 12218 57000
rect 12530 56200 12586 57000
rect 12898 56200 12954 57000
rect 13266 56200 13322 57000
rect 13634 56200 13690 57000
rect 14002 56200 14058 57000
rect 14370 56200 14426 57000
rect 14738 56200 14794 57000
rect 15106 56200 15162 57000
rect 15474 56200 15530 57000
rect 15842 56200 15898 57000
rect 16210 56200 16266 57000
rect 16578 56200 16634 57000
rect 16946 56200 17002 57000
rect 17314 56200 17370 57000
rect 17682 56200 17738 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 8128 56114 8156 56200
rect 8036 56086 8156 56114
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 7840 54256 7892 54262
rect 7840 54198 7892 54204
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 52556 7800 52562
rect 7748 52498 7800 52504
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8496 51950 8524 56200
rect 8864 53650 8892 56200
rect 8852 53644 8904 53650
rect 8852 53586 8904 53592
rect 9128 53576 9180 53582
rect 9128 53518 9180 53524
rect 8668 52488 8720 52494
rect 8668 52430 8720 52436
rect 8484 51944 8536 51950
rect 8484 51886 8536 51892
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7656 50924 7708 50930
rect 7656 50866 7708 50872
rect 7840 50924 7892 50930
rect 7840 50866 7892 50872
rect 7668 46102 7696 50866
rect 7748 49836 7800 49842
rect 7748 49778 7800 49784
rect 7656 46096 7708 46102
rect 7656 46038 7708 46044
rect 7564 44464 7616 44470
rect 7564 44406 7616 44412
rect 7472 44396 7524 44402
rect 7472 44338 7524 44344
rect 7380 40180 7432 40186
rect 7380 40122 7432 40128
rect 7380 40044 7432 40050
rect 7380 39986 7432 39992
rect 7288 38344 7340 38350
rect 7288 38286 7340 38292
rect 7288 37800 7340 37806
rect 7288 37742 7340 37748
rect 7300 35170 7328 37742
rect 7392 35290 7420 39986
rect 7484 36922 7512 44338
rect 7760 43450 7788 49778
rect 7852 44538 7880 50866
rect 8576 50244 8628 50250
rect 8576 50186 8628 50192
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 8484 44736 8536 44742
rect 8484 44678 8536 44684
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7840 44532 7892 44538
rect 7840 44474 7892 44480
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 7656 43308 7708 43314
rect 7656 43250 7708 43256
rect 8392 43308 8444 43314
rect 8392 43250 8444 43256
rect 7564 42016 7616 42022
rect 7564 41958 7616 41964
rect 7576 38554 7604 41958
rect 7564 38548 7616 38554
rect 7564 38490 7616 38496
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7668 36378 7696 43250
rect 8404 42566 8432 43250
rect 8392 42560 8444 42566
rect 8392 42502 8444 42508
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8116 42356 8168 42362
rect 8116 42298 8168 42304
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 7760 41818 7788 42094
rect 8128 41818 8156 42298
rect 7748 41812 7800 41818
rect 7748 41754 7800 41760
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 8116 41812 8168 41818
rect 8116 41754 8168 41760
rect 7748 41472 7800 41478
rect 7748 41414 7800 41420
rect 7760 40390 7788 41414
rect 7852 41274 7880 41754
rect 8300 41744 8352 41750
rect 8300 41686 8352 41692
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7840 41268 7892 41274
rect 7840 41210 7892 41216
rect 7748 40384 7800 40390
rect 7748 40326 7800 40332
rect 7852 40118 7880 41210
rect 8312 40390 8340 41686
rect 8300 40384 8352 40390
rect 8300 40326 8352 40332
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8312 40118 8340 40326
rect 7840 40112 7892 40118
rect 7840 40054 7892 40060
rect 7932 40112 7984 40118
rect 7932 40054 7984 40060
rect 8300 40112 8352 40118
rect 8300 40054 8352 40060
rect 7748 39976 7800 39982
rect 7748 39918 7800 39924
rect 7840 39976 7892 39982
rect 7840 39918 7892 39924
rect 7760 39642 7788 39918
rect 7748 39636 7800 39642
rect 7748 39578 7800 39584
rect 7748 38752 7800 38758
rect 7748 38694 7800 38700
rect 7760 38282 7788 38694
rect 7852 38418 7880 39918
rect 7944 39370 7972 40054
rect 7932 39364 7984 39370
rect 7932 39306 7984 39312
rect 8300 39296 8352 39302
rect 8300 39238 8352 39244
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7840 38412 7892 38418
rect 7840 38354 7892 38360
rect 8312 38350 8340 39238
rect 8404 38962 8432 42502
rect 8392 38956 8444 38962
rect 8392 38898 8444 38904
rect 8496 38894 8524 44678
rect 8588 40730 8616 50186
rect 8680 43450 8708 52430
rect 9036 52080 9088 52086
rect 9036 52022 9088 52028
rect 8944 49904 8996 49910
rect 8944 49846 8996 49852
rect 8852 49768 8904 49774
rect 8852 49710 8904 49716
rect 8864 45558 8892 49710
rect 8956 46986 8984 49846
rect 9048 47802 9076 52022
rect 9140 50522 9168 53518
rect 9232 53174 9260 56200
rect 9600 53564 9628 56200
rect 9968 54330 9996 56200
rect 9956 54324 10008 54330
rect 9956 54266 10008 54272
rect 9956 54188 10008 54194
rect 9956 54130 10008 54136
rect 9600 53536 9812 53564
rect 9220 53168 9272 53174
rect 9220 53110 9272 53116
rect 9312 53100 9364 53106
rect 9312 53042 9364 53048
rect 9220 51400 9272 51406
rect 9220 51342 9272 51348
rect 9128 50516 9180 50522
rect 9128 50458 9180 50464
rect 9036 47796 9088 47802
rect 9036 47738 9088 47744
rect 8944 46980 8996 46986
rect 8944 46922 8996 46928
rect 9232 46170 9260 51342
rect 9324 49910 9352 53042
rect 9588 52488 9640 52494
rect 9588 52430 9640 52436
rect 9600 50998 9628 52430
rect 9680 52012 9732 52018
rect 9680 51954 9732 51960
rect 9588 50992 9640 50998
rect 9588 50934 9640 50940
rect 9404 50312 9456 50318
rect 9404 50254 9456 50260
rect 9312 49904 9364 49910
rect 9312 49846 9364 49852
rect 9220 46164 9272 46170
rect 9220 46106 9272 46112
rect 9128 46028 9180 46034
rect 9128 45970 9180 45976
rect 8852 45552 8904 45558
rect 8852 45494 8904 45500
rect 8760 43648 8812 43654
rect 8760 43590 8812 43596
rect 8668 43444 8720 43450
rect 8668 43386 8720 43392
rect 8680 42906 8708 43386
rect 8772 43314 8800 43590
rect 8760 43308 8812 43314
rect 8760 43250 8812 43256
rect 8864 43246 8892 45494
rect 9036 43784 9088 43790
rect 9036 43726 9088 43732
rect 8852 43240 8904 43246
rect 8852 43182 8904 43188
rect 8864 42906 8892 43182
rect 8668 42900 8720 42906
rect 8668 42842 8720 42848
rect 8852 42900 8904 42906
rect 8852 42842 8904 42848
rect 8680 40730 8708 42842
rect 8576 40724 8628 40730
rect 8576 40666 8628 40672
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8588 40458 8616 40666
rect 8576 40452 8628 40458
rect 8576 40394 8628 40400
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8484 38888 8536 38894
rect 8484 38830 8536 38836
rect 8392 38752 8444 38758
rect 8392 38694 8444 38700
rect 8300 38344 8352 38350
rect 8206 38312 8262 38321
rect 7748 38276 7800 38282
rect 8300 38286 8352 38292
rect 8206 38247 8262 38256
rect 7748 38218 7800 38224
rect 7760 37890 7788 38218
rect 8220 38214 8248 38247
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 37936 7892 37942
rect 7760 37884 7840 37890
rect 7760 37878 7892 37884
rect 7760 37862 7880 37878
rect 7760 37194 7788 37862
rect 8404 37806 8432 38694
rect 8588 38486 8616 39374
rect 8680 39098 8708 40666
rect 8760 40180 8812 40186
rect 8760 40122 8812 40128
rect 8668 39092 8720 39098
rect 8668 39034 8720 39040
rect 8668 38956 8720 38962
rect 8668 38898 8720 38904
rect 8576 38480 8628 38486
rect 8576 38422 8628 38428
rect 8484 38208 8536 38214
rect 8484 38150 8536 38156
rect 8392 37800 8444 37806
rect 8392 37742 8444 37748
rect 7748 37188 7800 37194
rect 7748 37130 7800 37136
rect 7656 36372 7708 36378
rect 7656 36314 7708 36320
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7300 35142 7420 35170
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7196 34128 7248 34134
rect 7196 34070 7248 34076
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7208 33318 7236 33798
rect 7196 33312 7248 33318
rect 7196 33254 7248 33260
rect 7208 32978 7236 33254
rect 7196 32972 7248 32978
rect 7196 32914 7248 32920
rect 7104 31884 7156 31890
rect 7104 31826 7156 31832
rect 7116 29714 7144 31826
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 7300 29646 7328 34478
rect 7392 34202 7420 35142
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 7392 33998 7420 34138
rect 7380 33992 7432 33998
rect 7380 33934 7432 33940
rect 7392 31686 7420 33934
rect 7484 33114 7512 35974
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7576 33046 7604 36178
rect 7656 35488 7708 35494
rect 7760 35476 7788 37130
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 8496 36922 8524 38150
rect 8588 37466 8616 38422
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8484 36916 8536 36922
rect 8484 36858 8536 36864
rect 7840 36644 7892 36650
rect 7840 36586 7892 36592
rect 7852 36174 7880 36586
rect 7840 36168 7892 36174
rect 7840 36110 7892 36116
rect 7708 35448 7788 35476
rect 7656 35430 7708 35436
rect 7668 35018 7696 35430
rect 7852 35222 7880 36110
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 8588 35222 8616 37402
rect 8680 36258 8708 38898
rect 8772 37330 8800 40122
rect 8944 38004 8996 38010
rect 8944 37946 8996 37952
rect 8760 37324 8812 37330
rect 8760 37266 8812 37272
rect 8772 36582 8800 37266
rect 8760 36576 8812 36582
rect 8760 36518 8812 36524
rect 8956 36378 8984 37946
rect 9048 36922 9076 43726
rect 9140 43382 9168 45970
rect 9220 45484 9272 45490
rect 9220 45426 9272 45432
rect 9128 43376 9180 43382
rect 9128 43318 9180 43324
rect 9140 42906 9168 43318
rect 9128 42900 9180 42906
rect 9128 42842 9180 42848
rect 9232 42770 9260 45426
rect 9416 43994 9444 50254
rect 9588 46572 9640 46578
rect 9588 46514 9640 46520
rect 9494 44296 9550 44305
rect 9494 44231 9496 44240
rect 9548 44231 9550 44240
rect 9496 44202 9548 44208
rect 9404 43988 9456 43994
rect 9404 43930 9456 43936
rect 9404 43852 9456 43858
rect 9404 43794 9456 43800
rect 9496 43852 9548 43858
rect 9496 43794 9548 43800
rect 9312 43240 9364 43246
rect 9312 43182 9364 43188
rect 9128 42764 9180 42770
rect 9128 42706 9180 42712
rect 9220 42764 9272 42770
rect 9220 42706 9272 42712
rect 9140 42294 9168 42706
rect 9232 42362 9260 42706
rect 9220 42356 9272 42362
rect 9220 42298 9272 42304
rect 9128 42288 9180 42294
rect 9128 42230 9180 42236
rect 9140 41750 9168 42230
rect 9128 41744 9180 41750
rect 9128 41686 9180 41692
rect 9232 41682 9260 42298
rect 9220 41676 9272 41682
rect 9220 41618 9272 41624
rect 9220 41064 9272 41070
rect 9220 41006 9272 41012
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9140 38418 9168 38694
rect 9232 38486 9260 41006
rect 9220 38480 9272 38486
rect 9220 38422 9272 38428
rect 9128 38412 9180 38418
rect 9128 38354 9180 38360
rect 9220 38344 9272 38350
rect 9220 38286 9272 38292
rect 9036 36916 9088 36922
rect 9036 36858 9088 36864
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8758 36272 8814 36281
rect 8680 36230 8758 36258
rect 8758 36207 8814 36216
rect 7840 35216 7892 35222
rect 7840 35158 7892 35164
rect 8576 35216 8628 35222
rect 8576 35158 8628 35164
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 7656 35012 7708 35018
rect 7656 34954 7708 34960
rect 7840 34944 7892 34950
rect 7840 34886 7892 34892
rect 7852 34626 7880 34886
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8312 34746 8340 35022
rect 8668 35012 8720 35018
rect 8668 34954 8720 34960
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 7852 34610 7972 34626
rect 7852 34604 7984 34610
rect 7852 34598 7932 34604
rect 7932 34546 7984 34552
rect 7656 33924 7708 33930
rect 7656 33866 7708 33872
rect 7564 33040 7616 33046
rect 7564 32982 7616 32988
rect 7576 32298 7604 32982
rect 7564 32292 7616 32298
rect 7564 32234 7616 32240
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7668 31482 7696 33866
rect 7944 33862 7972 34546
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8300 33380 8352 33386
rect 8300 33322 8352 33328
rect 8312 32978 8340 33322
rect 8300 32972 8352 32978
rect 8300 32914 8352 32920
rect 7748 32836 7800 32842
rect 7748 32778 7800 32784
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7760 29850 7788 32778
rect 7840 32768 7892 32774
rect 7840 32710 7892 32716
rect 7852 32570 7880 32710
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 8312 32026 8340 32914
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8300 31816 8352 31822
rect 8300 31758 8352 31764
rect 8312 31686 8340 31758
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 8312 31362 8340 31622
rect 8680 31482 8708 34954
rect 8772 34542 8800 36207
rect 8852 35488 8904 35494
rect 8852 35430 8904 35436
rect 8864 34610 8892 35430
rect 8852 34604 8904 34610
rect 8852 34546 8904 34552
rect 8760 34536 8812 34542
rect 8760 34478 8812 34484
rect 8864 33998 8892 34546
rect 9140 34202 9168 36722
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9232 34066 9260 38286
rect 9324 38010 9352 43182
rect 9416 42770 9444 43794
rect 9508 43246 9536 43794
rect 9496 43240 9548 43246
rect 9496 43182 9548 43188
rect 9496 42900 9548 42906
rect 9496 42842 9548 42848
rect 9404 42764 9456 42770
rect 9404 42706 9456 42712
rect 9416 41274 9444 42706
rect 9404 41268 9456 41274
rect 9404 41210 9456 41216
rect 9508 40390 9536 42842
rect 9600 42362 9628 46514
rect 9692 44538 9720 51954
rect 9784 51950 9812 53536
rect 9772 51944 9824 51950
rect 9772 51886 9824 51892
rect 9968 51610 9996 54130
rect 10336 53038 10364 56200
rect 10324 53032 10376 53038
rect 10324 52974 10376 52980
rect 10704 52562 10732 56200
rect 11072 53650 11100 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11244 54120 11296 54126
rect 11244 54062 11296 54068
rect 11060 53644 11112 53650
rect 11060 53586 11112 53592
rect 10692 52556 10744 52562
rect 10692 52498 10744 52504
rect 10876 52012 10928 52018
rect 10876 51954 10928 51960
rect 10416 51876 10468 51882
rect 10416 51818 10468 51824
rect 9956 51604 10008 51610
rect 9956 51546 10008 51552
rect 9864 49972 9916 49978
rect 9864 49914 9916 49920
rect 9876 47258 9904 49914
rect 9956 48136 10008 48142
rect 9956 48078 10008 48084
rect 9864 47252 9916 47258
rect 9864 47194 9916 47200
rect 9876 45642 9904 47194
rect 9784 45614 9904 45642
rect 9784 45558 9812 45614
rect 9772 45552 9824 45558
rect 9772 45494 9824 45500
rect 9876 45422 9904 45614
rect 9864 45416 9916 45422
rect 9864 45358 9916 45364
rect 9772 44736 9824 44742
rect 9770 44704 9772 44713
rect 9824 44704 9826 44713
rect 9770 44639 9826 44648
rect 9680 44532 9732 44538
rect 9680 44474 9732 44480
rect 9968 43994 9996 48078
rect 10048 45960 10100 45966
rect 10048 45902 10100 45908
rect 9956 43988 10008 43994
rect 9956 43930 10008 43936
rect 9772 43308 9824 43314
rect 9772 43250 9824 43256
rect 9680 42628 9732 42634
rect 9680 42570 9732 42576
rect 9588 42356 9640 42362
rect 9588 42298 9640 42304
rect 9588 42220 9640 42226
rect 9588 42162 9640 42168
rect 9600 42090 9628 42162
rect 9588 42084 9640 42090
rect 9588 42026 9640 42032
rect 9692 42022 9720 42570
rect 9680 42016 9732 42022
rect 9680 41958 9732 41964
rect 9692 41478 9720 41958
rect 9680 41472 9732 41478
rect 9680 41414 9732 41420
rect 9496 40384 9548 40390
rect 9496 40326 9548 40332
rect 9312 38004 9364 38010
rect 9312 37946 9364 37952
rect 9312 36780 9364 36786
rect 9312 36722 9364 36728
rect 9220 34060 9272 34066
rect 9220 34002 9272 34008
rect 8852 33992 8904 33998
rect 8852 33934 8904 33940
rect 9324 33114 9352 36722
rect 9508 36650 9536 40326
rect 9588 38888 9640 38894
rect 9588 38830 9640 38836
rect 9600 37670 9628 38830
rect 9680 38276 9732 38282
rect 9680 38218 9732 38224
rect 9692 37913 9720 38218
rect 9678 37904 9734 37913
rect 9678 37839 9734 37848
rect 9588 37664 9640 37670
rect 9588 37606 9640 37612
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 9496 36644 9548 36650
rect 9496 36586 9548 36592
rect 9404 36576 9456 36582
rect 9404 36518 9456 36524
rect 9416 35873 9444 36518
rect 9402 35864 9458 35873
rect 9402 35799 9458 35808
rect 9600 35630 9628 36654
rect 9784 36378 9812 43250
rect 9956 40928 10008 40934
rect 9956 40870 10008 40876
rect 9968 39982 9996 40870
rect 9956 39976 10008 39982
rect 9956 39918 10008 39924
rect 10060 39914 10088 45902
rect 10428 43450 10456 51818
rect 10692 49224 10744 49230
rect 10692 49166 10744 49172
rect 10508 46980 10560 46986
rect 10508 46922 10560 46928
rect 10520 45354 10548 46922
rect 10600 46912 10652 46918
rect 10600 46854 10652 46860
rect 10612 45490 10640 46854
rect 10704 46170 10732 49166
rect 10784 49088 10836 49094
rect 10784 49030 10836 49036
rect 10796 46594 10824 49030
rect 10888 46714 10916 51954
rect 10876 46708 10928 46714
rect 10876 46650 10928 46656
rect 10796 46566 10916 46594
rect 10692 46164 10744 46170
rect 10692 46106 10744 46112
rect 10600 45484 10652 45490
rect 10600 45426 10652 45432
rect 10508 45348 10560 45354
rect 10508 45290 10560 45296
rect 10612 43704 10640 45426
rect 10692 43716 10744 43722
rect 10612 43676 10692 43704
rect 10692 43658 10744 43664
rect 10416 43444 10468 43450
rect 10416 43386 10468 43392
rect 10704 43382 10732 43658
rect 10888 43654 10916 46566
rect 11060 46572 11112 46578
rect 11060 46514 11112 46520
rect 10876 43648 10928 43654
rect 10876 43590 10928 43596
rect 10692 43376 10744 43382
rect 10692 43318 10744 43324
rect 10324 43308 10376 43314
rect 10324 43250 10376 43256
rect 10336 42566 10364 43250
rect 10704 42906 10732 43318
rect 10692 42900 10744 42906
rect 10692 42842 10744 42848
rect 10324 42560 10376 42566
rect 10322 42528 10324 42537
rect 10376 42528 10378 42537
rect 10322 42463 10378 42472
rect 10508 42016 10560 42022
rect 10508 41958 10560 41964
rect 10520 41614 10548 41958
rect 10600 41676 10652 41682
rect 10600 41618 10652 41624
rect 10784 41676 10836 41682
rect 10784 41618 10836 41624
rect 10508 41608 10560 41614
rect 10508 41550 10560 41556
rect 10520 41414 10548 41550
rect 10428 41386 10548 41414
rect 10232 40656 10284 40662
rect 10232 40598 10284 40604
rect 10048 39908 10100 39914
rect 10048 39850 10100 39856
rect 10244 39506 10272 40598
rect 10324 40588 10376 40594
rect 10324 40530 10376 40536
rect 10336 40390 10364 40530
rect 10324 40384 10376 40390
rect 10324 40326 10376 40332
rect 10336 40186 10364 40326
rect 10324 40180 10376 40186
rect 10324 40122 10376 40128
rect 10232 39500 10284 39506
rect 10232 39442 10284 39448
rect 10140 39296 10192 39302
rect 10140 39238 10192 39244
rect 10152 39001 10180 39238
rect 10138 38992 10194 39001
rect 10138 38927 10194 38936
rect 10428 37466 10456 41386
rect 10508 41132 10560 41138
rect 10508 41074 10560 41080
rect 10520 38010 10548 41074
rect 10612 40730 10640 41618
rect 10796 41562 10824 41618
rect 10704 41534 10824 41562
rect 10704 40934 10732 41534
rect 10784 41472 10836 41478
rect 10784 41414 10836 41420
rect 10692 40928 10744 40934
rect 10692 40870 10744 40876
rect 10600 40724 10652 40730
rect 10600 40666 10652 40672
rect 10692 39840 10744 39846
rect 10692 39782 10744 39788
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10612 38214 10640 38286
rect 10600 38208 10652 38214
rect 10600 38150 10652 38156
rect 10508 38004 10560 38010
rect 10508 37946 10560 37952
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 10416 37460 10468 37466
rect 10416 37402 10468 37408
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 9954 36816 10010 36825
rect 9954 36751 10010 36760
rect 9772 36372 9824 36378
rect 9772 36314 9824 36320
rect 9588 35624 9640 35630
rect 9508 35572 9588 35578
rect 9508 35566 9640 35572
rect 9508 35550 9628 35566
rect 9508 34746 9536 35550
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9772 35488 9824 35494
rect 9772 35430 9824 35436
rect 9496 34740 9548 34746
rect 9496 34682 9548 34688
rect 9600 34678 9628 35430
rect 9784 35154 9812 35430
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 9588 34672 9640 34678
rect 9588 34614 9640 34620
rect 9600 34542 9628 34614
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9588 33992 9640 33998
rect 9588 33934 9640 33940
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9128 33040 9180 33046
rect 9128 32982 9180 32988
rect 9140 32502 9168 32982
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 9140 32026 9168 32438
rect 9220 32224 9272 32230
rect 9220 32166 9272 32172
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 9232 31958 9260 32166
rect 9220 31952 9272 31958
rect 9220 31894 9272 31900
rect 9128 31680 9180 31686
rect 9232 31668 9260 31894
rect 9180 31640 9260 31668
rect 9128 31622 9180 31628
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 8128 31334 8340 31362
rect 8760 31340 8812 31346
rect 7852 30802 7880 31282
rect 8128 31278 8156 31334
rect 8760 31282 8812 31288
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8484 31272 8536 31278
rect 8484 31214 8536 31220
rect 8128 30938 8156 31214
rect 8116 30932 8168 30938
rect 8116 30874 8168 30880
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 8496 30598 8524 31214
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7656 29844 7708 29850
rect 7656 29786 7708 29792
rect 7748 29844 7800 29850
rect 7748 29786 7800 29792
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 19310 6868 23462
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6932 21418 6960 22578
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6932 17134 6960 17682
rect 7024 17218 7052 29514
rect 7668 29510 7696 29786
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7392 24818 7420 29446
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7576 27062 7604 27406
rect 7564 27056 7616 27062
rect 7564 26998 7616 27004
rect 7576 26330 7604 26998
rect 7484 26314 7604 26330
rect 7472 26308 7604 26314
rect 7524 26302 7604 26308
rect 7472 26250 7524 26256
rect 7576 26042 7604 26302
rect 7668 26246 7696 29242
rect 7852 27606 7880 29582
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8128 28404 8156 28494
rect 8208 28416 8260 28422
rect 8128 28376 8208 28404
rect 8260 28376 8340 28404
rect 8208 28358 8260 28364
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 8312 27606 8340 28376
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 7852 26926 7880 27542
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 26920 7892 26926
rect 7760 26880 7840 26908
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 7564 26036 7616 26042
rect 7564 25978 7616 25984
rect 7668 25498 7696 26182
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 7484 24886 7512 25434
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7472 24880 7524 24886
rect 7472 24822 7524 24828
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7116 21690 7144 24142
rect 7668 23866 7696 25298
rect 7760 24818 7788 26880
rect 7840 26862 7892 26868
rect 8300 26852 8352 26858
rect 8300 26794 8352 26800
rect 8312 26450 8340 26794
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 8496 25906 8524 30534
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8680 28014 8708 28902
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 8668 28008 8720 28014
rect 8668 27950 8720 27956
rect 8588 26586 8616 27950
rect 8668 26920 8720 26926
rect 8772 26908 8800 31282
rect 9140 29714 9168 31622
rect 9508 29850 9536 32710
rect 9600 31754 9628 33934
rect 9876 33930 9904 34478
rect 9864 33924 9916 33930
rect 9864 33866 9916 33872
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9784 32910 9812 33390
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9588 31748 9640 31754
rect 9588 31690 9640 31696
rect 9600 31278 9628 31690
rect 9876 31482 9904 32302
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 9600 30802 9628 31214
rect 9588 30796 9640 30802
rect 9588 30738 9640 30744
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 9600 29578 9628 30262
rect 9312 29572 9364 29578
rect 9312 29514 9364 29520
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 8720 26880 8800 26908
rect 8668 26862 8720 26868
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7852 24954 7880 25774
rect 8588 25770 8616 26522
rect 8680 26314 8708 26862
rect 9140 26450 9168 26930
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 8668 26308 8720 26314
rect 8668 26250 8720 26256
rect 8760 26308 8812 26314
rect 8760 26250 8812 26256
rect 8576 25764 8628 25770
rect 8576 25706 8628 25712
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 8116 24744 8168 24750
rect 8116 24686 8168 24692
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 8128 24562 8156 24686
rect 8404 24682 8432 25230
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7576 23322 7604 23598
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7484 22522 7512 22918
rect 7576 22658 7604 23258
rect 7576 22642 7696 22658
rect 7564 22636 7696 22642
rect 7616 22630 7696 22636
rect 7564 22578 7616 22584
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7300 21146 7328 22510
rect 7484 22494 7604 22522
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7116 19854 7144 20470
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19446 7144 19790
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 7392 17882 7420 19654
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7024 17190 7236 17218
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16794 6960 17070
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 8090 6868 13262
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5828 2746 6040 2774
rect 6012 2446 6040 2746
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5736 800 5764 2314
rect 6104 800 6132 3470
rect 6564 3194 6592 3470
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6564 2774 6592 3130
rect 6840 3058 6868 3334
rect 7024 3194 7052 16934
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7116 9518 7144 13466
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6472 2746 6592 2774
rect 6472 800 6500 2746
rect 6840 800 6868 2994
rect 7116 2650 7144 5646
rect 7208 3194 7236 17190
rect 7300 16250 7328 17478
rect 7484 16998 7512 22374
rect 7576 21350 7604 22494
rect 7668 21622 7696 22630
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7668 19786 7696 21422
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18222 7604 19110
rect 7760 18426 7788 24550
rect 8128 24534 8432 24562
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7852 19854 7880 23122
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 21010 8248 21286
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19922 8340 20198
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7484 16590 7512 16730
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7484 16182 7512 16526
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7576 13530 7604 18158
rect 7852 17746 7880 19450
rect 8404 19378 8432 24534
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8496 20874 8524 24346
rect 8588 24342 8616 25094
rect 8576 24336 8628 24342
rect 8576 24278 8628 24284
rect 8588 23662 8616 24278
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8680 20466 8708 26250
rect 8772 26042 8800 26250
rect 8760 26036 8812 26042
rect 8760 25978 8812 25984
rect 8772 25498 8800 25978
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9048 24138 9076 25434
rect 9324 24750 9352 29514
rect 9968 29510 9996 36751
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9416 28558 9444 29038
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9416 26926 9444 28494
rect 9876 27674 9904 28562
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9968 27878 9996 28494
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9680 26852 9732 26858
rect 9680 26794 9732 26800
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9416 25362 9444 25842
rect 9692 25362 9720 26794
rect 9876 25838 9904 27610
rect 9968 27470 9996 27814
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 26382 9996 27406
rect 10060 27062 10088 37198
rect 10428 37194 10456 37402
rect 10416 37188 10468 37194
rect 10416 37130 10468 37136
rect 10428 36854 10456 37130
rect 10416 36848 10468 36854
rect 10416 36790 10468 36796
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10152 32978 10180 34342
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 10244 33114 10272 34070
rect 10336 33658 10364 36042
rect 10416 34536 10468 34542
rect 10416 34478 10468 34484
rect 10428 33998 10456 34478
rect 10416 33992 10468 33998
rect 10416 33934 10468 33940
rect 10324 33652 10376 33658
rect 10324 33594 10376 33600
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10152 32026 10180 32914
rect 10232 32496 10284 32502
rect 10232 32438 10284 32444
rect 10244 32230 10272 32438
rect 10232 32224 10284 32230
rect 10232 32166 10284 32172
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10244 31906 10272 32166
rect 10152 31878 10272 31906
rect 10152 31754 10180 31878
rect 10140 31748 10192 31754
rect 10140 31690 10192 31696
rect 10152 30580 10180 31690
rect 10232 30592 10284 30598
rect 10152 30552 10232 30580
rect 10232 30534 10284 30540
rect 10244 29238 10272 30534
rect 10520 30190 10548 37742
rect 10704 36106 10732 39782
rect 10796 39642 10824 41414
rect 10784 39636 10836 39642
rect 10784 39578 10836 39584
rect 10796 38962 10824 39578
rect 10784 38956 10836 38962
rect 10784 38898 10836 38904
rect 10888 38570 10916 43590
rect 10968 43376 11020 43382
rect 10968 43318 11020 43324
rect 10980 41274 11008 43318
rect 11072 41818 11100 46514
rect 11152 45824 11204 45830
rect 11152 45766 11204 45772
rect 11164 44538 11192 45766
rect 11256 45082 11284 54062
rect 11808 53038 11836 56200
rect 12176 53650 12204 56200
rect 12348 54188 12400 54194
rect 12348 54130 12400 54136
rect 12256 53984 12308 53990
rect 12256 53926 12308 53932
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 12072 53576 12124 53582
rect 12072 53518 12124 53524
rect 11888 53100 11940 53106
rect 11888 53042 11940 53048
rect 11796 53032 11848 53038
rect 11796 52974 11848 52980
rect 11900 52154 11928 53042
rect 11888 52148 11940 52154
rect 11888 52090 11940 52096
rect 11980 52012 12032 52018
rect 11980 51954 12032 51960
rect 11992 49434 12020 51954
rect 11980 49428 12032 49434
rect 11980 49370 12032 49376
rect 11796 47660 11848 47666
rect 11796 47602 11848 47608
rect 11704 45892 11756 45898
rect 11704 45834 11756 45840
rect 11244 45076 11296 45082
rect 11244 45018 11296 45024
rect 11152 44532 11204 44538
rect 11152 44474 11204 44480
rect 11612 44396 11664 44402
rect 11612 44338 11664 44344
rect 11152 44328 11204 44334
rect 11152 44270 11204 44276
rect 11164 43178 11192 44270
rect 11624 44198 11652 44338
rect 11612 44192 11664 44198
rect 11612 44134 11664 44140
rect 11428 43716 11480 43722
rect 11428 43658 11480 43664
rect 11152 43172 11204 43178
rect 11152 43114 11204 43120
rect 11152 42220 11204 42226
rect 11152 42162 11204 42168
rect 11060 41812 11112 41818
rect 11060 41754 11112 41760
rect 11060 41472 11112 41478
rect 11060 41414 11112 41420
rect 10968 41268 11020 41274
rect 10968 41210 11020 41216
rect 10980 40186 11008 41210
rect 10968 40180 11020 40186
rect 10968 40122 11020 40128
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 10980 39098 11008 39918
rect 10968 39092 11020 39098
rect 10968 39034 11020 39040
rect 10888 38542 11008 38570
rect 11072 38554 11100 41414
rect 11164 38826 11192 42162
rect 11244 40724 11296 40730
rect 11244 40666 11296 40672
rect 11256 40458 11284 40666
rect 11244 40452 11296 40458
rect 11244 40394 11296 40400
rect 11256 39658 11284 40394
rect 11256 39630 11376 39658
rect 11244 39364 11296 39370
rect 11244 39306 11296 39312
rect 11256 38826 11284 39306
rect 11152 38820 11204 38826
rect 11152 38762 11204 38768
rect 11244 38820 11296 38826
rect 11244 38762 11296 38768
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 10876 38208 10928 38214
rect 10876 38150 10928 38156
rect 10796 38010 10824 38150
rect 10784 38004 10836 38010
rect 10784 37946 10836 37952
rect 10784 36916 10836 36922
rect 10784 36858 10836 36864
rect 10692 36100 10744 36106
rect 10692 36042 10744 36048
rect 10692 34196 10744 34202
rect 10692 34138 10744 34144
rect 10704 31754 10732 34138
rect 10796 33658 10824 36858
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10888 33114 10916 38150
rect 10980 37330 11008 38542
rect 11060 38548 11112 38554
rect 11060 38490 11112 38496
rect 11242 38312 11298 38321
rect 11242 38247 11298 38256
rect 11256 37618 11284 38247
rect 11348 37942 11376 39630
rect 11336 37936 11388 37942
rect 11336 37878 11388 37884
rect 11348 37738 11376 37878
rect 11336 37732 11388 37738
rect 11336 37674 11388 37680
rect 11256 37590 11376 37618
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 10968 36712 11020 36718
rect 10968 36654 11020 36660
rect 10980 35630 11008 36654
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10980 34542 11008 35566
rect 11072 35290 11100 36722
rect 11244 36032 11296 36038
rect 11244 35974 11296 35980
rect 11060 35284 11112 35290
rect 11060 35226 11112 35232
rect 11060 35148 11112 35154
rect 11060 35090 11112 35096
rect 10968 34536 11020 34542
rect 10968 34478 11020 34484
rect 11072 34474 11100 35090
rect 11060 34468 11112 34474
rect 11060 34410 11112 34416
rect 10968 34400 11020 34406
rect 10968 34342 11020 34348
rect 10980 33930 11008 34342
rect 10968 33924 11020 33930
rect 10968 33866 11020 33872
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10980 32502 11008 33866
rect 11256 33658 11284 35974
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 11348 33538 11376 37590
rect 11256 33510 11376 33538
rect 11256 33436 11284 33510
rect 11072 33408 11284 33436
rect 10968 32496 11020 32502
rect 10968 32438 11020 32444
rect 10612 31726 10732 31754
rect 10612 30802 10640 31726
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10612 30122 10640 30738
rect 10692 30184 10744 30190
rect 10692 30126 10744 30132
rect 10600 30116 10652 30122
rect 10600 30058 10652 30064
rect 10416 30048 10468 30054
rect 10704 30002 10732 30126
rect 10416 29990 10468 29996
rect 10428 29646 10456 29990
rect 10612 29974 10732 30002
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10232 29232 10284 29238
rect 10232 29174 10284 29180
rect 10244 28422 10272 29174
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 28218 10272 28358
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10048 27056 10100 27062
rect 10048 26998 10100 27004
rect 10244 26450 10272 27270
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 9956 26376 10008 26382
rect 9956 26318 10008 26324
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9324 24410 9352 24686
rect 9312 24404 9364 24410
rect 9312 24346 9364 24352
rect 9862 24304 9918 24313
rect 9862 24239 9864 24248
rect 9916 24239 9918 24248
rect 9864 24210 9916 24216
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8772 22778 8800 24006
rect 9048 23730 9076 24074
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23798 9812 24006
rect 9968 23866 9996 26318
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9048 23322 9076 23666
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9968 23118 9996 23530
rect 10152 23526 10180 24686
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8680 19718 8708 20402
rect 8772 20330 8800 21422
rect 8864 20602 8892 22510
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8956 20602 8984 21490
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8864 19922 8892 20538
rect 9048 20534 9076 21422
rect 9128 21140 9180 21146
rect 9128 21082 9180 21088
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9048 20262 9076 20470
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8956 19718 8984 19790
rect 8668 19712 8720 19718
rect 8666 19680 8668 19689
rect 8944 19712 8996 19718
rect 8720 19680 8722 19689
rect 8944 19654 8996 19660
rect 8666 19615 8722 19624
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8864 18630 8892 19314
rect 8956 18902 8984 19654
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8496 18222 8524 18566
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16794 8340 17002
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16726 8432 17682
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16046 8340 16526
rect 8404 16046 8432 16662
rect 8496 16658 8524 18158
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 16794 8616 17478
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16454 8524 16594
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8496 15366 8524 16390
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 8496 13394 8524 15302
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8404 12986 8432 13262
rect 8680 12986 8708 18022
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8772 17202 8800 17478
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8772 15706 8800 16662
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 15162 8800 15642
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 14006 8800 15098
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8772 13870 8800 13942
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8772 13530 8800 13806
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8772 13326 8800 13466
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12442 8708 12786
rect 8772 12782 8800 13126
rect 8864 12850 8892 18566
rect 8956 17066 8984 18838
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8942 16144 8998 16153
rect 8942 16079 8998 16088
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8956 12594 8984 16079
rect 8864 12566 8984 12594
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8206 4176 8262 4185
rect 8206 4111 8262 4120
rect 8220 3738 8248 4111
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7208 800 7236 2382
rect 7576 800 7604 2382
rect 7852 1986 7880 3470
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8208 3052 8260 3058
rect 8312 3040 8340 3402
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3058 8708 3334
rect 8864 3194 8892 12566
rect 9140 12458 9168 21082
rect 9220 20392 9272 20398
rect 9272 20352 9352 20380
rect 9220 20334 9272 20340
rect 9324 19446 9352 20352
rect 9416 19514 9444 22442
rect 9784 21690 9812 22918
rect 9968 22778 9996 23054
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 17202 9260 19246
rect 9968 18426 9996 22714
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 10060 21146 10088 22646
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10244 20890 10272 24346
rect 10060 20874 10272 20890
rect 10048 20868 10272 20874
rect 10100 20862 10272 20868
rect 10048 20810 10100 20816
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16590 9260 17138
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9324 16726 9352 16934
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9416 15094 9444 17682
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9508 17338 9536 17478
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9600 16590 9628 17614
rect 9876 17270 9904 18226
rect 9968 17678 9996 18362
rect 10060 18290 10088 20810
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 10152 16794 10180 17478
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10244 16674 10272 19110
rect 10152 16646 10272 16674
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 15706 9996 16390
rect 9956 15700 10008 15706
rect 10008 15660 10088 15688
rect 9956 15642 10008 15648
rect 9404 15088 9456 15094
rect 9456 15048 9536 15076
rect 9404 15030 9456 15036
rect 9508 13870 9536 15048
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14482 9996 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9876 13734 9904 14214
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9864 13388 9916 13394
rect 9968 13376 9996 14010
rect 9916 13348 9996 13376
rect 9864 13330 9916 13336
rect 9968 12918 9996 13348
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 8956 12430 9168 12458
rect 8956 3602 8984 12430
rect 9692 12306 9720 12854
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 10060 10742 10088 15660
rect 10152 11082 10180 16646
rect 10336 16522 10364 26794
rect 10428 22953 10456 29446
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10520 26042 10548 26726
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 10508 23792 10560 23798
rect 10508 23734 10560 23740
rect 10414 22944 10470 22953
rect 10414 22879 10470 22888
rect 10520 22438 10548 23734
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10612 21894 10640 29974
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10796 25294 10824 29446
rect 10876 29028 10928 29034
rect 10876 28970 10928 28976
rect 10888 26042 10916 28970
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10980 26994 11008 27406
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 11072 24698 11100 33408
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 11256 31414 11284 31894
rect 11440 31890 11468 43658
rect 11520 38752 11572 38758
rect 11518 38720 11520 38729
rect 11572 38720 11574 38729
rect 11518 38655 11574 38664
rect 11624 35034 11652 44134
rect 11716 41274 11744 45834
rect 11808 42362 11836 47602
rect 11888 46368 11940 46374
rect 11888 46310 11940 46316
rect 11900 46034 11928 46310
rect 11888 46028 11940 46034
rect 11888 45970 11940 45976
rect 12084 45082 12112 53518
rect 12164 46912 12216 46918
rect 12164 46854 12216 46860
rect 12176 46034 12204 46854
rect 12164 46028 12216 46034
rect 12164 45970 12216 45976
rect 12164 45416 12216 45422
rect 12164 45358 12216 45364
rect 12072 45076 12124 45082
rect 12072 45018 12124 45024
rect 12176 44266 12204 45358
rect 12164 44260 12216 44266
rect 12164 44202 12216 44208
rect 11796 42356 11848 42362
rect 11796 42298 11848 42304
rect 11888 42288 11940 42294
rect 11888 42230 11940 42236
rect 11704 41268 11756 41274
rect 11704 41210 11756 41216
rect 11704 40180 11756 40186
rect 11704 40122 11756 40128
rect 11716 37466 11744 40122
rect 11900 38554 11928 42230
rect 12176 41290 12204 44202
rect 12268 41426 12296 53926
rect 12360 52154 12388 54130
rect 12544 54126 12572 56200
rect 12912 54262 12940 56200
rect 13280 55214 13308 56200
rect 13280 55186 13400 55214
rect 12900 54256 12952 54262
rect 12900 54198 12952 54204
rect 12532 54120 12584 54126
rect 12532 54062 12584 54068
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12624 53576 12676 53582
rect 12624 53518 12676 53524
rect 12636 52698 12664 53518
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12624 52692 12676 52698
rect 12624 52634 12676 52640
rect 12808 52488 12860 52494
rect 12808 52430 12860 52436
rect 12348 52148 12400 52154
rect 12348 52090 12400 52096
rect 12820 48890 12848 52430
rect 13372 52426 13400 55186
rect 13648 53174 13676 56200
rect 14016 53582 14044 56200
rect 14004 53576 14056 53582
rect 14004 53518 14056 53524
rect 13636 53168 13688 53174
rect 13636 53110 13688 53116
rect 13648 52698 13676 53110
rect 14384 53106 14412 56200
rect 14752 54330 14780 56200
rect 14740 54324 14792 54330
rect 14740 54266 14792 54272
rect 15120 54176 15148 56200
rect 15200 54188 15252 54194
rect 15120 54148 15200 54176
rect 15200 54130 15252 54136
rect 14924 53984 14976 53990
rect 14924 53926 14976 53932
rect 15200 53984 15252 53990
rect 15200 53926 15252 53932
rect 14464 53440 14516 53446
rect 14464 53382 14516 53388
rect 14372 53100 14424 53106
rect 14372 53042 14424 53048
rect 14004 52964 14056 52970
rect 14004 52906 14056 52912
rect 13636 52692 13688 52698
rect 13636 52634 13688 52640
rect 14016 52601 14044 52906
rect 14476 52601 14504 53382
rect 14740 52896 14792 52902
rect 14740 52838 14792 52844
rect 14002 52592 14058 52601
rect 14002 52527 14058 52536
rect 14462 52592 14518 52601
rect 14462 52527 14518 52536
rect 13544 52488 13596 52494
rect 13544 52430 13596 52436
rect 13360 52420 13412 52426
rect 13360 52362 13412 52368
rect 13372 52154 13400 52362
rect 13360 52148 13412 52154
rect 13360 52090 13412 52096
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12808 48884 12860 48890
rect 12808 48826 12860 48832
rect 12808 48748 12860 48754
rect 12808 48690 12860 48696
rect 12624 46980 12676 46986
rect 12624 46922 12676 46928
rect 12636 46628 12664 46922
rect 12716 46640 12768 46646
rect 12636 46600 12716 46628
rect 12636 46034 12664 46600
rect 12716 46582 12768 46588
rect 12716 46368 12768 46374
rect 12716 46310 12768 46316
rect 12624 46028 12676 46034
rect 12624 45970 12676 45976
rect 12636 45898 12664 45970
rect 12624 45892 12676 45898
rect 12624 45834 12676 45840
rect 12348 45280 12400 45286
rect 12348 45222 12400 45228
rect 12360 44878 12388 45222
rect 12624 44940 12676 44946
rect 12624 44882 12676 44888
rect 12348 44872 12400 44878
rect 12348 44814 12400 44820
rect 12532 44804 12584 44810
rect 12532 44746 12584 44752
rect 12348 44464 12400 44470
rect 12348 44406 12400 44412
rect 12360 43246 12388 44406
rect 12348 43240 12400 43246
rect 12348 43182 12400 43188
rect 12360 42770 12388 43182
rect 12348 42764 12400 42770
rect 12348 42706 12400 42712
rect 12360 41682 12388 42706
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 12452 42158 12480 42502
rect 12440 42152 12492 42158
rect 12440 42094 12492 42100
rect 12348 41676 12400 41682
rect 12348 41618 12400 41624
rect 12268 41398 12480 41426
rect 12176 41262 12296 41290
rect 12268 41070 12296 41262
rect 12348 41132 12400 41138
rect 12348 41074 12400 41080
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 12256 40452 12308 40458
rect 12256 40394 12308 40400
rect 12164 40384 12216 40390
rect 12164 40326 12216 40332
rect 12072 38752 12124 38758
rect 12072 38694 12124 38700
rect 11888 38548 11940 38554
rect 11888 38490 11940 38496
rect 11796 38004 11848 38010
rect 11796 37946 11848 37952
rect 11704 37460 11756 37466
rect 11704 37402 11756 37408
rect 11808 36174 11836 37946
rect 11886 37360 11942 37369
rect 11886 37295 11942 37304
rect 11900 37262 11928 37295
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 12084 36258 12112 38694
rect 12176 38418 12204 40326
rect 12268 40186 12296 40394
rect 12256 40180 12308 40186
rect 12256 40122 12308 40128
rect 12254 39128 12310 39137
rect 12254 39063 12256 39072
rect 12308 39063 12310 39072
rect 12256 39034 12308 39040
rect 12360 38842 12388 41074
rect 12452 40526 12480 41398
rect 12440 40520 12492 40526
rect 12440 40462 12492 40468
rect 12440 39500 12492 39506
rect 12440 39442 12492 39448
rect 12452 39030 12480 39442
rect 12440 39024 12492 39030
rect 12440 38966 12492 38972
rect 12268 38814 12388 38842
rect 12164 38412 12216 38418
rect 12164 38354 12216 38360
rect 12268 37466 12296 38814
rect 12346 38720 12402 38729
rect 12402 38678 12480 38706
rect 12346 38655 12402 38664
rect 12348 38548 12400 38554
rect 12348 38490 12400 38496
rect 12256 37460 12308 37466
rect 12256 37402 12308 37408
rect 12360 37233 12388 38490
rect 12452 37398 12480 38678
rect 12544 38554 12572 44746
rect 12636 43382 12664 44882
rect 12728 44470 12756 46310
rect 12820 45082 12848 48690
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 13452 45824 13504 45830
rect 13452 45766 13504 45772
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12808 45076 12860 45082
rect 12808 45018 12860 45024
rect 13360 44736 13412 44742
rect 13360 44678 13412 44684
rect 12716 44464 12768 44470
rect 12716 44406 12768 44412
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12624 43376 12676 43382
rect 12624 43318 12676 43324
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 13372 42362 13400 44678
rect 13464 44470 13492 45766
rect 13452 44464 13504 44470
rect 13452 44406 13504 44412
rect 13464 44334 13492 44406
rect 13452 44328 13504 44334
rect 13452 44270 13504 44276
rect 13360 42356 13412 42362
rect 13360 42298 13412 42304
rect 13360 42084 13412 42090
rect 13360 42026 13412 42032
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12808 41676 12860 41682
rect 12808 41618 12860 41624
rect 12820 41478 12848 41618
rect 12808 41472 12860 41478
rect 12808 41414 12860 41420
rect 12624 40384 12676 40390
rect 12624 40326 12676 40332
rect 12532 38548 12584 38554
rect 12532 38490 12584 38496
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12346 37224 12402 37233
rect 12346 37159 12402 37168
rect 12256 36916 12308 36922
rect 12256 36858 12308 36864
rect 12268 36650 12296 36858
rect 12256 36644 12308 36650
rect 12256 36586 12308 36592
rect 12084 36230 12204 36258
rect 11796 36168 11848 36174
rect 11796 36110 11848 36116
rect 12072 36168 12124 36174
rect 12072 36110 12124 36116
rect 11888 35760 11940 35766
rect 11888 35702 11940 35708
rect 11532 35006 11652 35034
rect 11532 32978 11560 35006
rect 11900 34678 11928 35702
rect 11888 34672 11940 34678
rect 11808 34632 11888 34660
rect 11808 34406 11836 34632
rect 11888 34614 11940 34620
rect 12084 34406 12112 36110
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 11808 33998 11836 34342
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11980 33856 12032 33862
rect 11980 33798 12032 33804
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11624 32026 11652 33458
rect 11888 32836 11940 32842
rect 11888 32778 11940 32784
rect 11612 32020 11664 32026
rect 11612 31962 11664 31968
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 11244 31408 11296 31414
rect 11244 31350 11296 31356
rect 11428 30728 11480 30734
rect 11426 30696 11428 30705
rect 11480 30696 11482 30705
rect 11426 30631 11482 30640
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11348 29782 11376 30534
rect 11796 30320 11848 30326
rect 11796 30262 11848 30268
rect 11336 29776 11388 29782
rect 11336 29718 11388 29724
rect 11348 28626 11376 29718
rect 11808 29578 11836 30262
rect 11900 30138 11928 32778
rect 11992 30938 12020 33798
rect 12084 32298 12112 34342
rect 12176 33114 12204 36230
rect 12360 36224 12388 37159
rect 12440 36236 12492 36242
rect 12360 36196 12440 36224
rect 12440 36178 12492 36184
rect 12452 36145 12480 36178
rect 12438 36136 12494 36145
rect 12256 36100 12308 36106
rect 12438 36071 12494 36080
rect 12256 36042 12308 36048
rect 12164 33108 12216 33114
rect 12164 33050 12216 33056
rect 12268 32366 12296 36042
rect 12544 35578 12572 38150
rect 12452 35550 12572 35578
rect 12452 33538 12480 35550
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12544 34066 12572 35430
rect 12636 34066 12664 40326
rect 12820 40050 12848 41414
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12716 39908 12768 39914
rect 12716 39850 12768 39856
rect 12728 39574 12756 39850
rect 12716 39568 12768 39574
rect 12716 39510 12768 39516
rect 12820 39506 12848 39986
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12808 39500 12860 39506
rect 12808 39442 12860 39448
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12728 38486 12756 39238
rect 12912 39030 12940 39374
rect 13084 39296 13136 39302
rect 13084 39238 13136 39244
rect 12990 39128 13046 39137
rect 12990 39063 12992 39072
rect 13044 39063 13046 39072
rect 12992 39034 13044 39040
rect 12900 39024 12952 39030
rect 12900 38966 12952 38972
rect 13096 38758 13124 39238
rect 13084 38752 13136 38758
rect 13084 38694 13136 38700
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12716 38480 12768 38486
rect 12716 38422 12768 38428
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 13280 38049 13308 38150
rect 13266 38040 13322 38049
rect 13266 37975 13268 37984
rect 13320 37975 13322 37984
rect 13268 37946 13320 37952
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12808 37392 12860 37398
rect 12992 37392 13044 37398
rect 12860 37352 12992 37380
rect 12808 37334 12860 37340
rect 12992 37334 13044 37340
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12728 36854 12756 37062
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 12808 36780 12860 36786
rect 12808 36722 12860 36728
rect 12716 36712 12768 36718
rect 12716 36654 12768 36660
rect 12728 35086 12756 36654
rect 12716 35080 12768 35086
rect 12716 35022 12768 35028
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12452 33510 12572 33538
rect 12438 33416 12494 33425
rect 12438 33351 12494 33360
rect 12452 33318 12480 33351
rect 12440 33312 12492 33318
rect 12440 33254 12492 33260
rect 12256 32360 12308 32366
rect 12254 32328 12256 32337
rect 12308 32328 12310 32337
rect 12072 32292 12124 32298
rect 12254 32263 12310 32272
rect 12072 32234 12124 32240
rect 11980 30932 12032 30938
rect 11980 30874 12032 30880
rect 11900 30110 12020 30138
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11900 29510 11928 29990
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11244 27940 11296 27946
rect 11244 27882 11296 27888
rect 11256 26450 11284 27882
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11440 25702 11468 27338
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11336 25696 11388 25702
rect 11336 25638 11388 25644
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11072 24670 11284 24698
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10692 24064 10744 24070
rect 10968 24064 11020 24070
rect 10744 24024 10824 24052
rect 10692 24006 10744 24012
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10704 23050 10732 23802
rect 10796 23526 10824 24024
rect 10968 24006 11020 24012
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10888 23118 10916 23598
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10692 23044 10744 23050
rect 10692 22986 10744 22992
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10428 18426 10456 20742
rect 10612 18970 10640 21830
rect 10704 21010 10732 22986
rect 10796 22953 10824 22986
rect 10782 22944 10838 22953
rect 10782 22879 10838 22888
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10704 18306 10732 20742
rect 10428 18278 10732 18306
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10428 16402 10456 18278
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10520 17338 10548 17614
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10336 16374 10456 16402
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10244 15706 10272 15914
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10244 14346 10272 15642
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 13258 10272 13874
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10244 12918 10272 13194
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9586 5672 9642 5681
rect 9586 5607 9642 5616
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9048 3058 9076 3946
rect 9324 3738 9352 4218
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9508 3534 9536 3878
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 8260 3012 8340 3040
rect 8208 2994 8260 3000
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 7852 1958 7972 1986
rect 7944 800 7972 1958
rect 8312 800 8340 3012
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8680 800 8708 2994
rect 9048 800 9076 2994
rect 9508 2774 9536 3470
rect 9600 3058 9628 5607
rect 9862 5536 9918 5545
rect 9862 5471 9918 5480
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9784 3534 9812 3878
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9416 2746 9536 2774
rect 9416 800 9444 2746
rect 9784 800 9812 3470
rect 9876 2650 9904 5471
rect 10060 3738 10088 8366
rect 10336 4282 10364 16374
rect 10520 16250 10548 17070
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10428 15366 10456 16050
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10428 13870 10456 15302
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10520 14346 10548 14758
rect 10704 14600 10732 18158
rect 10796 18154 10824 21354
rect 10980 19718 11008 24006
rect 11072 21486 11100 24210
rect 11164 24206 11192 24550
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11256 23866 11284 24670
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11164 21894 11192 22510
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11256 21010 11284 23666
rect 11348 21418 11376 25638
rect 11440 25362 11468 25638
rect 11532 25498 11560 27066
rect 11796 25832 11848 25838
rect 11796 25774 11848 25780
rect 11520 25492 11572 25498
rect 11520 25434 11572 25440
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11808 25294 11836 25774
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11900 25140 11928 29446
rect 11992 25158 12020 30110
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 11808 25112 11928 25140
rect 11980 25152 12032 25158
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11716 22982 11744 23598
rect 11808 23526 11836 25112
rect 11980 25094 12032 25100
rect 12176 24342 12204 26182
rect 12452 25498 12480 33254
rect 12544 32502 12572 33510
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12532 32496 12584 32502
rect 12532 32438 12584 32444
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12544 26353 12572 32166
rect 12530 26344 12586 26353
rect 12530 26279 12586 26288
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25974 12572 26182
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12636 25378 12664 32982
rect 12728 32230 12756 35022
rect 12820 33998 12848 36722
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 13372 36378 13400 42026
rect 13556 38214 13584 52430
rect 14464 46708 14516 46714
rect 14464 46650 14516 46656
rect 13728 46368 13780 46374
rect 13728 46310 13780 46316
rect 13740 44946 13768 46310
rect 14096 46028 14148 46034
rect 14096 45970 14148 45976
rect 14108 45558 14136 45970
rect 14096 45552 14148 45558
rect 14096 45494 14148 45500
rect 13728 44940 13780 44946
rect 13728 44882 13780 44888
rect 14108 44470 14136 45494
rect 14372 45416 14424 45422
rect 14372 45358 14424 45364
rect 14384 45014 14412 45358
rect 14372 45008 14424 45014
rect 14372 44950 14424 44956
rect 14372 44872 14424 44878
rect 14372 44814 14424 44820
rect 14096 44464 14148 44470
rect 14096 44406 14148 44412
rect 14108 43382 14136 44406
rect 14096 43376 14148 43382
rect 14096 43318 14148 43324
rect 13728 43172 13780 43178
rect 13728 43114 13780 43120
rect 13636 41472 13688 41478
rect 13636 41414 13688 41420
rect 13648 41138 13676 41414
rect 13636 41132 13688 41138
rect 13636 41074 13688 41080
rect 13636 40588 13688 40594
rect 13636 40530 13688 40536
rect 13544 38208 13596 38214
rect 13544 38150 13596 38156
rect 13452 37800 13504 37806
rect 13452 37742 13504 37748
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13360 36372 13412 36378
rect 13360 36314 13412 36320
rect 13084 36304 13136 36310
rect 13084 36246 13136 36252
rect 13096 36038 13124 36246
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13084 36032 13136 36038
rect 13084 35974 13136 35980
rect 13372 35698 13400 36178
rect 13464 35834 13492 37742
rect 13556 37262 13584 37742
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 13544 36848 13596 36854
rect 13544 36790 13596 36796
rect 13556 36242 13584 36790
rect 13544 36236 13596 36242
rect 13544 36178 13596 36184
rect 13648 36122 13676 40530
rect 13740 36922 13768 43114
rect 13912 43104 13964 43110
rect 13912 43046 13964 43052
rect 13924 40730 13952 43046
rect 14108 42906 14136 43318
rect 14096 42900 14148 42906
rect 14096 42842 14148 42848
rect 14004 41540 14056 41546
rect 14004 41482 14056 41488
rect 14016 41154 14044 41482
rect 14016 41126 14228 41154
rect 14004 41064 14056 41070
rect 14056 41024 14136 41052
rect 14004 41006 14056 41012
rect 13912 40724 13964 40730
rect 13912 40666 13964 40672
rect 13820 39500 13872 39506
rect 13820 39442 13872 39448
rect 13832 38321 13860 39442
rect 13924 39302 13952 40666
rect 13912 39296 13964 39302
rect 13912 39238 13964 39244
rect 14004 38820 14056 38826
rect 14004 38762 14056 38768
rect 13912 38752 13964 38758
rect 13912 38694 13964 38700
rect 13818 38312 13874 38321
rect 13818 38247 13874 38256
rect 13820 38208 13872 38214
rect 13820 38150 13872 38156
rect 13728 36916 13780 36922
rect 13728 36858 13780 36864
rect 13556 36094 13676 36122
rect 13452 35828 13504 35834
rect 13452 35770 13504 35776
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 13360 34944 13412 34950
rect 13360 34886 13412 34892
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12808 33856 12860 33862
rect 12808 33798 12860 33804
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12820 29578 12848 33798
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 13280 33318 13308 33458
rect 13268 33312 13320 33318
rect 13268 33254 13320 33260
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31482 13400 34886
rect 13464 33454 13492 35770
rect 13556 35562 13584 36094
rect 13636 36032 13688 36038
rect 13636 35974 13688 35980
rect 13544 35556 13596 35562
rect 13544 35498 13596 35504
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13452 33448 13504 33454
rect 13452 33390 13504 33396
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13268 31272 13320 31278
rect 13464 31260 13492 33254
rect 13556 32298 13584 33798
rect 13544 32292 13596 32298
rect 13544 32234 13596 32240
rect 13320 31232 13492 31260
rect 13268 31214 13320 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12900 29844 12952 29850
rect 12900 29786 12952 29792
rect 12808 29572 12860 29578
rect 12808 29514 12860 29520
rect 12912 29306 12940 29786
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13372 28626 13400 31232
rect 13544 29300 13596 29306
rect 13544 29242 13596 29248
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 13360 28620 13412 28626
rect 13360 28562 13412 28568
rect 12728 27878 12756 28562
rect 12808 28416 12860 28422
rect 12808 28358 12860 28364
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 12716 27872 12768 27878
rect 12716 27814 12768 27820
rect 12728 27402 12756 27814
rect 12820 27538 12848 28358
rect 13188 28218 13216 28358
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13280 28082 13308 28358
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 13280 27962 13308 28018
rect 13280 27934 13400 27962
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12716 27396 12768 27402
rect 12716 27338 12768 27344
rect 12820 26926 12848 27474
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 12912 26926 12940 27270
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12452 25350 12664 25378
rect 12820 25362 12848 26862
rect 13004 26790 13032 27270
rect 13372 27146 13400 27934
rect 13096 27118 13400 27146
rect 13096 27062 13124 27118
rect 13084 27056 13136 27062
rect 13084 26998 13136 27004
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13372 26314 13400 27118
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13464 25378 13492 28970
rect 13556 26450 13584 29242
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 12808 25356 12860 25362
rect 12452 24818 12480 25350
rect 12808 25298 12860 25304
rect 13372 25350 13492 25378
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 12164 24336 12216 24342
rect 12164 24278 12216 24284
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11808 23066 11836 23462
rect 11808 23038 11928 23066
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11428 22160 11480 22166
rect 11428 22102 11480 22108
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 11256 19310 11284 20946
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18834 11100 19110
rect 11256 18970 11284 19246
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10888 16590 10916 18566
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10980 16640 11008 17070
rect 11060 16652 11112 16658
rect 10980 16612 11060 16640
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 14958 10916 15302
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14612 10836 14618
rect 10704 14572 10784 14600
rect 10784 14554 10836 14560
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10520 13938 10548 14282
rect 10796 14226 10824 14554
rect 10704 14198 10824 14226
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10336 3058 10364 3878
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10336 2774 10364 2994
rect 10428 2990 10456 13806
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10612 12986 10640 13194
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10704 6866 10732 14198
rect 10888 12442 10916 14894
rect 10980 14278 11008 16612
rect 11060 16594 11112 16600
rect 11164 16046 11192 18294
rect 11348 18290 11376 18838
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10876 12436 10928 12442
rect 11256 12434 11284 18022
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11348 17134 11376 17546
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11348 15570 11376 17070
rect 11440 16250 11468 22102
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11532 21010 11560 21830
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11808 20534 11836 22102
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11532 16250 11560 20470
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11716 20058 11744 20402
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11808 19922 11836 20470
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11716 19394 11744 19790
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11624 19366 11744 19394
rect 11624 18630 11652 19366
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11624 18358 11652 18566
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11704 17672 11756 17678
rect 11808 17660 11836 19722
rect 11756 17632 11836 17660
rect 11704 17614 11756 17620
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 14550 11376 15506
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11624 13530 11652 16730
rect 11716 15366 11744 17614
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16182 11836 16390
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11808 14822 11836 15370
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 14550 11836 14758
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11900 14006 11928 23038
rect 11992 21690 12020 24006
rect 12084 23866 12112 24006
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12268 23474 12296 24550
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12084 23446 12296 23474
rect 12084 22710 12112 23446
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11992 19786 12020 20946
rect 12176 20330 12204 23122
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12268 22166 12296 22918
rect 12360 22642 12388 23802
rect 12452 23662 12480 24754
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 11978 19544 12034 19553
rect 11978 19479 12034 19488
rect 11992 19378 12020 19479
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12918 11560 13126
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11256 12406 11376 12434
rect 10876 12378 10928 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 11762 11008 12242
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10336 2746 10548 2774
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 800 10180 2382
rect 10520 800 10548 2746
rect 10888 800 10916 3470
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 800 11284 3334
rect 11348 3194 11376 12406
rect 11624 6458 11652 13466
rect 11808 12986 11836 13738
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 12306 11836 12922
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11992 5710 12020 17818
rect 12084 17270 12112 20198
rect 12176 19922 12204 20266
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12162 19408 12218 19417
rect 12162 19343 12218 19352
rect 12176 18970 12204 19343
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12176 18426 12204 18906
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11624 800 11652 4014
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3058 11744 3334
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11808 2938 11836 4626
rect 11716 2910 11836 2938
rect 11716 2514 11744 2910
rect 12084 2774 12112 16458
rect 12176 15162 12204 18158
rect 12268 16658 12296 21014
rect 12360 20806 12388 21422
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12360 18222 12388 20742
rect 12452 19854 12480 22986
rect 12544 22094 12572 25230
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12636 24954 12664 25094
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 12636 24206 12664 24618
rect 12820 24274 12848 25094
rect 13096 24886 13124 25230
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 12912 24614 12940 24822
rect 12992 24744 13044 24750
rect 12990 24712 12992 24721
rect 13044 24712 13046 24721
rect 12990 24647 13046 24656
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22642 13124 22918
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12544 22066 12664 22094
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12544 17338 12572 20470
rect 12636 17882 12664 22066
rect 12820 21622 12848 22374
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12912 21434 12940 21830
rect 12820 21406 12940 21434
rect 13280 21434 13308 22170
rect 13372 22030 13400 25350
rect 13556 24818 13584 26250
rect 13648 25362 13676 35974
rect 13832 35714 13860 38150
rect 13924 37126 13952 38694
rect 13912 37120 13964 37126
rect 13912 37062 13964 37068
rect 14016 36718 14044 38762
rect 14108 37330 14136 41024
rect 14200 38554 14228 41126
rect 14280 39432 14332 39438
rect 14280 39374 14332 39380
rect 14188 38548 14240 38554
rect 14188 38490 14240 38496
rect 14292 38457 14320 39374
rect 14278 38448 14334 38457
rect 14278 38383 14280 38392
rect 14332 38383 14334 38392
rect 14280 38354 14332 38360
rect 14280 37732 14332 37738
rect 14280 37674 14332 37680
rect 14292 37369 14320 37674
rect 14384 37670 14412 44814
rect 14476 44538 14504 46650
rect 14464 44532 14516 44538
rect 14464 44474 14516 44480
rect 14476 42158 14504 44474
rect 14556 44192 14608 44198
rect 14556 44134 14608 44140
rect 14568 42566 14596 44134
rect 14752 43450 14780 52838
rect 14740 43444 14792 43450
rect 14740 43386 14792 43392
rect 14648 43308 14700 43314
rect 14648 43250 14700 43256
rect 14556 42560 14608 42566
rect 14556 42502 14608 42508
rect 14464 42152 14516 42158
rect 14464 42094 14516 42100
rect 14464 42016 14516 42022
rect 14464 41958 14516 41964
rect 14476 39030 14504 41958
rect 14556 40112 14608 40118
rect 14556 40054 14608 40060
rect 14568 39438 14596 40054
rect 14660 39846 14688 43250
rect 14648 39840 14700 39846
rect 14648 39782 14700 39788
rect 14556 39432 14608 39438
rect 14556 39374 14608 39380
rect 14464 39024 14516 39030
rect 14464 38966 14516 38972
rect 14372 37664 14424 37670
rect 14372 37606 14424 37612
rect 14476 37398 14504 38966
rect 14660 38894 14688 39782
rect 14832 39024 14884 39030
rect 14832 38966 14884 38972
rect 14648 38888 14700 38894
rect 14648 38830 14700 38836
rect 14464 37392 14516 37398
rect 14278 37360 14334 37369
rect 14096 37324 14148 37330
rect 14096 37266 14148 37272
rect 14188 37324 14240 37330
rect 14464 37334 14516 37340
rect 14278 37295 14334 37304
rect 14188 37266 14240 37272
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14108 36786 14136 37062
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14004 36712 14056 36718
rect 14004 36654 14056 36660
rect 14016 36174 14044 36654
rect 14004 36168 14056 36174
rect 14004 36110 14056 36116
rect 14200 35873 14228 37266
rect 14476 36922 14504 37334
rect 14464 36916 14516 36922
rect 14464 36858 14516 36864
rect 14844 36786 14872 38966
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14464 36576 14516 36582
rect 14464 36518 14516 36524
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14186 35864 14242 35873
rect 14186 35799 14242 35808
rect 13832 35686 13952 35714
rect 13820 35624 13872 35630
rect 13820 35566 13872 35572
rect 13728 35488 13780 35494
rect 13728 35430 13780 35436
rect 13740 34746 13768 35430
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13832 34542 13860 35566
rect 13820 34536 13872 34542
rect 13820 34478 13872 34484
rect 13820 34128 13872 34134
rect 13820 34070 13872 34076
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13740 29306 13768 33934
rect 13832 33658 13860 34070
rect 13820 33652 13872 33658
rect 13820 33594 13872 33600
rect 13924 33046 13952 35686
rect 14200 34898 14228 35799
rect 14280 35012 14332 35018
rect 14280 34954 14332 34960
rect 14108 34870 14228 34898
rect 13912 33040 13964 33046
rect 13912 32982 13964 32988
rect 14108 31958 14136 34870
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 14096 31952 14148 31958
rect 14096 31894 14148 31900
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13832 31686 13860 31826
rect 13820 31680 13872 31686
rect 13820 31622 13872 31628
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13556 23866 13584 24754
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13452 23656 13504 23662
rect 13452 23598 13504 23604
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13280 21406 13400 21434
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 18834 12756 20334
rect 12820 19514 12848 21406
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12898 19952 12954 19961
rect 12898 19887 12954 19896
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12636 17678 12664 17818
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12256 16652 12308 16658
rect 12544 16640 12572 17138
rect 12624 16652 12676 16658
rect 12544 16612 12624 16640
rect 12256 16594 12308 16600
rect 12624 16594 12676 16600
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12360 13530 12388 15846
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 12176 3670 12204 3946
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12452 3534 12480 15642
rect 12544 15094 12572 16186
rect 12636 15366 12664 16594
rect 12728 16590 12756 17478
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12820 16436 12848 19450
rect 12912 19281 12940 19887
rect 12898 19272 12954 19281
rect 13372 19242 13400 21406
rect 12898 19207 12954 19216
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18426 13400 18566
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12728 16408 12848 16436
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 6914 12572 14418
rect 12636 13394 12664 15302
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12728 12434 12756 16408
rect 13372 16250 13400 17070
rect 13464 16250 13492 23598
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13556 22234 13584 23122
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 20466 13676 25162
rect 13740 24614 13768 29106
rect 14016 28966 14044 29446
rect 14200 29306 14228 34682
rect 14292 31958 14320 34954
rect 14372 34672 14424 34678
rect 14372 34614 14424 34620
rect 14384 33590 14412 34614
rect 14372 33584 14424 33590
rect 14372 33526 14424 33532
rect 14372 33108 14424 33114
rect 14372 33050 14424 33056
rect 14384 32842 14412 33050
rect 14476 32978 14504 36518
rect 14568 35086 14596 36518
rect 14648 36032 14700 36038
rect 14648 35974 14700 35980
rect 14660 35834 14688 35974
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 14372 32836 14424 32842
rect 14372 32778 14424 32784
rect 14384 32609 14412 32778
rect 14370 32600 14426 32609
rect 14370 32535 14426 32544
rect 14568 32434 14596 33594
rect 14648 33584 14700 33590
rect 14700 33544 14780 33572
rect 14648 33526 14700 33532
rect 14752 33289 14780 33544
rect 14738 33280 14794 33289
rect 14738 33215 14794 33224
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14660 32570 14688 32710
rect 14752 32570 14780 33215
rect 14844 32978 14872 34478
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14740 32564 14792 32570
rect 14740 32506 14792 32512
rect 14832 32496 14884 32502
rect 14832 32438 14884 32444
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14568 32230 14596 32370
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14280 31952 14332 31958
rect 14280 31894 14332 31900
rect 14476 31754 14504 32166
rect 14648 31952 14700 31958
rect 14648 31894 14700 31900
rect 14660 31822 14688 31894
rect 14648 31816 14700 31822
rect 14648 31758 14700 31764
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14464 31748 14516 31754
rect 14464 31690 14516 31696
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 14370 30288 14426 30297
rect 14188 29300 14240 29306
rect 14188 29242 14240 29248
rect 14292 29170 14320 30262
rect 14476 30258 14504 31078
rect 14370 30223 14372 30232
rect 14424 30223 14426 30232
rect 14464 30252 14516 30258
rect 14372 30194 14424 30200
rect 14464 30194 14516 30200
rect 14464 29708 14516 29714
rect 14464 29650 14516 29656
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14280 29164 14332 29170
rect 14280 29106 14332 29112
rect 14004 28960 14056 28966
rect 14004 28902 14056 28908
rect 14016 28422 14044 28902
rect 14108 28762 14136 29106
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13912 26444 13964 26450
rect 13912 26386 13964 26392
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13740 21486 13768 24278
rect 13832 24138 13860 24754
rect 13924 24721 13952 26386
rect 13910 24712 13966 24721
rect 13910 24647 13966 24656
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13924 23050 13952 23802
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 13832 21690 13860 22578
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21690 13952 22510
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 18358 13584 19110
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 14618 12848 16050
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13464 15502 13492 16186
rect 13556 16182 13584 17478
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13372 14346 13400 14962
rect 13464 14482 13492 15030
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 12806 13968 12862 13977
rect 12806 13903 12862 13912
rect 12820 13870 12848 13903
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13530 12848 13806
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13280 12986 13308 13398
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13280 12832 13308 12922
rect 13280 12804 13492 12832
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12728 12406 13400 12434
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11694 13216 12038
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12544 6886 12664 6914
rect 12636 4690 12664 6886
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12636 3058 12664 4422
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 11808 2746 12112 2774
rect 11808 2582 11836 2746
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11992 800 12020 2450
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12360 800 12388 2314
rect 12728 800 12756 3538
rect 12820 2446 12848 10474
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13372 10062 13400 12406
rect 13464 12170 13492 12804
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11898 13492 12106
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13556 4282 13584 14010
rect 13648 12850 13676 20198
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19446 13768 19654
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13832 18766 13860 21286
rect 13924 20534 13952 21490
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 13924 20074 13952 20266
rect 14016 20262 14044 28358
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 27062 14136 27270
rect 14096 27056 14148 27062
rect 14096 26998 14148 27004
rect 14108 26246 14136 26998
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14200 22094 14228 28902
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14292 26382 14320 28358
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14280 26376 14332 26382
rect 14280 26318 14332 26324
rect 14384 25838 14412 26726
rect 14476 25838 14504 29650
rect 14660 29102 14688 31078
rect 14752 29866 14780 31758
rect 14844 30190 14872 32438
rect 14936 31278 14964 53926
rect 15108 46640 15160 46646
rect 15108 46582 15160 46588
rect 15120 45558 15148 46582
rect 15108 45552 15160 45558
rect 15108 45494 15160 45500
rect 15120 44810 15148 45494
rect 15108 44804 15160 44810
rect 15108 44746 15160 44752
rect 15120 44538 15148 44746
rect 15108 44532 15160 44538
rect 15108 44474 15160 44480
rect 15016 39364 15068 39370
rect 15016 39306 15068 39312
rect 15028 39098 15056 39306
rect 15212 39250 15240 53926
rect 15488 53582 15516 56200
rect 15568 54052 15620 54058
rect 15568 53994 15620 54000
rect 15476 53576 15528 53582
rect 15476 53518 15528 53524
rect 15292 44736 15344 44742
rect 15292 44678 15344 44684
rect 15304 42362 15332 44678
rect 15580 43450 15608 53994
rect 15856 53106 15884 56200
rect 16224 54330 16252 56200
rect 16212 54324 16264 54330
rect 16212 54266 16264 54272
rect 16592 53786 16620 56200
rect 16960 54194 16988 56200
rect 16948 54188 17000 54194
rect 16948 54130 17000 54136
rect 17040 53984 17092 53990
rect 17038 53952 17040 53961
rect 17092 53952 17094 53961
rect 17038 53887 17094 53896
rect 16580 53780 16632 53786
rect 16580 53722 16632 53728
rect 16592 53582 16620 53722
rect 17328 53582 17356 56200
rect 17696 54262 17724 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17684 54256 17736 54262
rect 17684 54198 17736 54204
rect 18340 53582 18368 56222
rect 18418 56200 18474 57000
rect 18786 56200 18842 57000
rect 19154 56200 19210 57000
rect 19522 56200 19578 57000
rect 19890 56200 19946 57000
rect 20258 56200 20314 57000
rect 20626 56200 20682 57000
rect 20994 56200 21050 57000
rect 21362 56200 21418 57000
rect 21730 56200 21786 57000
rect 22098 56200 22154 57000
rect 22466 56200 22522 57000
rect 22834 56200 22890 57000
rect 23202 56200 23258 57000
rect 23570 56200 23626 57000
rect 18432 54126 18460 56200
rect 18420 54120 18472 54126
rect 18420 54062 18472 54068
rect 18420 53984 18472 53990
rect 18420 53926 18472 53932
rect 16580 53576 16632 53582
rect 16580 53518 16632 53524
rect 17316 53576 17368 53582
rect 17316 53518 17368 53524
rect 18328 53576 18380 53582
rect 18328 53518 18380 53524
rect 16396 53508 16448 53514
rect 16396 53450 16448 53456
rect 15844 53100 15896 53106
rect 15844 53042 15896 53048
rect 15936 52896 15988 52902
rect 15936 52838 15988 52844
rect 15948 47802 15976 52838
rect 16408 52601 16436 53450
rect 16856 53440 16908 53446
rect 16856 53382 16908 53388
rect 16394 52592 16450 52601
rect 16394 52527 16450 52536
rect 16868 49774 16896 53382
rect 17328 53242 17356 53518
rect 17408 53440 17460 53446
rect 17408 53382 17460 53388
rect 17316 53236 17368 53242
rect 17316 53178 17368 53184
rect 16028 49768 16080 49774
rect 16028 49710 16080 49716
rect 16856 49768 16908 49774
rect 16856 49710 16908 49716
rect 15936 47796 15988 47802
rect 15936 47738 15988 47744
rect 15568 43444 15620 43450
rect 15488 43404 15568 43432
rect 15292 42356 15344 42362
rect 15292 42298 15344 42304
rect 15292 41744 15344 41750
rect 15292 41686 15344 41692
rect 15304 41070 15332 41686
rect 15384 41200 15436 41206
rect 15384 41142 15436 41148
rect 15292 41064 15344 41070
rect 15292 41006 15344 41012
rect 15396 40474 15424 41142
rect 15304 40446 15424 40474
rect 15304 40118 15332 40446
rect 15384 40384 15436 40390
rect 15384 40326 15436 40332
rect 15292 40112 15344 40118
rect 15292 40054 15344 40060
rect 15212 39222 15332 39250
rect 15016 39092 15068 39098
rect 15016 39034 15068 39040
rect 15016 38412 15068 38418
rect 15016 38354 15068 38360
rect 15028 36242 15056 38354
rect 15200 37664 15252 37670
rect 15200 37606 15252 37612
rect 15212 37126 15240 37606
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15200 37120 15252 37126
rect 15200 37062 15252 37068
rect 15120 36718 15148 37062
rect 15108 36712 15160 36718
rect 15108 36654 15160 36660
rect 15016 36236 15068 36242
rect 15016 36178 15068 36184
rect 15016 35828 15068 35834
rect 15016 35770 15068 35776
rect 15028 33862 15056 35770
rect 15016 33856 15068 33862
rect 15016 33798 15068 33804
rect 15016 33108 15068 33114
rect 15016 33050 15068 33056
rect 15028 31686 15056 33050
rect 15120 31958 15148 36654
rect 15212 34678 15240 37062
rect 15200 34672 15252 34678
rect 15200 34614 15252 34620
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15108 31952 15160 31958
rect 15108 31894 15160 31900
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 14924 31272 14976 31278
rect 14924 31214 14976 31220
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 14752 29838 14872 29866
rect 14740 29776 14792 29782
rect 14740 29718 14792 29724
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14556 28416 14608 28422
rect 14556 28358 14608 28364
rect 14568 27878 14596 28358
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14372 25832 14424 25838
rect 14372 25774 14424 25780
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14384 24750 14412 25774
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22098 14320 23122
rect 14568 22098 14596 27814
rect 14752 24138 14780 29718
rect 14844 28762 14872 29838
rect 14936 29510 14964 31214
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 15028 29322 15056 31622
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 15120 30598 15148 31350
rect 15212 30802 15240 32166
rect 15304 31754 15332 39222
rect 15396 38350 15424 40326
rect 15488 39386 15516 43404
rect 15568 43386 15620 43392
rect 15660 43240 15712 43246
rect 15660 43182 15712 43188
rect 15568 42288 15620 42294
rect 15568 42230 15620 42236
rect 15580 40186 15608 42230
rect 15568 40180 15620 40186
rect 15568 40122 15620 40128
rect 15672 39506 15700 43182
rect 16040 41414 16068 49710
rect 17420 47802 17448 53382
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 18432 48006 18460 53926
rect 18512 53508 18564 53514
rect 18512 53450 18564 53456
rect 17592 48000 17644 48006
rect 17592 47942 17644 47948
rect 18420 48000 18472 48006
rect 18420 47942 18472 47948
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 17604 47666 17632 47942
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 18524 47666 18552 53450
rect 18800 53106 18828 56200
rect 18880 54256 18932 54262
rect 18880 54198 18932 54204
rect 18892 53786 18920 54198
rect 18880 53780 18932 53786
rect 18880 53722 18932 53728
rect 19168 53582 19196 56200
rect 19536 54194 19564 56200
rect 19524 54188 19576 54194
rect 19524 54130 19576 54136
rect 19708 54120 19760 54126
rect 19708 54062 19760 54068
rect 19340 53984 19392 53990
rect 19340 53926 19392 53932
rect 19156 53576 19208 53582
rect 19156 53518 19208 53524
rect 19168 53242 19196 53518
rect 19156 53236 19208 53242
rect 19156 53178 19208 53184
rect 18788 53100 18840 53106
rect 18788 53042 18840 53048
rect 18604 52896 18656 52902
rect 18604 52838 18656 52844
rect 17592 47660 17644 47666
rect 17592 47602 17644 47608
rect 18512 47660 18564 47666
rect 18512 47602 18564 47608
rect 16304 47524 16356 47530
rect 16304 47466 16356 47472
rect 16316 46374 16344 47466
rect 16580 47456 16632 47462
rect 16580 47398 16632 47404
rect 17500 47456 17552 47462
rect 17500 47398 17552 47404
rect 16396 46980 16448 46986
rect 16396 46922 16448 46928
rect 16408 46646 16436 46922
rect 16396 46640 16448 46646
rect 16396 46582 16448 46588
rect 16304 46368 16356 46374
rect 16304 46310 16356 46316
rect 16316 45422 16344 46310
rect 16408 45830 16436 46582
rect 16396 45824 16448 45830
rect 16396 45766 16448 45772
rect 16408 45626 16436 45766
rect 16396 45620 16448 45626
rect 16396 45562 16448 45568
rect 16304 45416 16356 45422
rect 16304 45358 16356 45364
rect 16120 45280 16172 45286
rect 16120 45222 16172 45228
rect 16132 41750 16160 45222
rect 16396 43648 16448 43654
rect 16396 43590 16448 43596
rect 16212 43376 16264 43382
rect 16212 43318 16264 43324
rect 16224 42702 16252 43318
rect 16212 42696 16264 42702
rect 16212 42638 16264 42644
rect 16120 41744 16172 41750
rect 16120 41686 16172 41692
rect 16224 41562 16252 42638
rect 15948 41386 16068 41414
rect 16132 41534 16252 41562
rect 15752 40996 15804 41002
rect 15752 40938 15804 40944
rect 15764 39982 15792 40938
rect 15844 40588 15896 40594
rect 15844 40530 15896 40536
rect 15752 39976 15804 39982
rect 15752 39918 15804 39924
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15488 39358 15700 39386
rect 15476 39296 15528 39302
rect 15476 39238 15528 39244
rect 15384 38344 15436 38350
rect 15384 38286 15436 38292
rect 15384 38004 15436 38010
rect 15384 37946 15436 37952
rect 15396 37330 15424 37946
rect 15384 37324 15436 37330
rect 15384 37266 15436 37272
rect 15396 36922 15424 37266
rect 15384 36916 15436 36922
rect 15384 36858 15436 36864
rect 15488 36378 15516 39238
rect 15672 38962 15700 39358
rect 15660 38956 15712 38962
rect 15660 38898 15712 38904
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15580 37806 15608 38830
rect 15568 37800 15620 37806
rect 15568 37742 15620 37748
rect 15568 37120 15620 37126
rect 15568 37062 15620 37068
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15580 35737 15608 37062
rect 15566 35728 15622 35737
rect 15566 35663 15622 35672
rect 15568 33924 15620 33930
rect 15568 33866 15620 33872
rect 15580 32824 15608 33866
rect 15488 32796 15608 32824
rect 15304 31726 15424 31754
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15200 30796 15252 30802
rect 15200 30738 15252 30744
rect 15304 30705 15332 31078
rect 15290 30696 15346 30705
rect 15290 30631 15346 30640
rect 15108 30592 15160 30598
rect 15108 30534 15160 30540
rect 15120 30308 15148 30534
rect 15200 30320 15252 30326
rect 15120 30280 15200 30308
rect 15200 30262 15252 30268
rect 14936 29294 15056 29322
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14832 28620 14884 28626
rect 14832 28562 14884 28568
rect 14844 26518 14872 28562
rect 14832 26512 14884 26518
rect 14832 26454 14884 26460
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14844 25974 14872 26182
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 14740 24132 14792 24138
rect 14740 24074 14792 24080
rect 14648 23316 14700 23322
rect 14648 23258 14700 23264
rect 14108 22066 14228 22094
rect 14280 22092 14332 22098
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13924 20046 14044 20074
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13924 19242 13952 19858
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13924 18902 13952 19178
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13740 18290 13768 18566
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13740 18193 13768 18226
rect 13820 18216 13872 18222
rect 13726 18184 13782 18193
rect 13820 18158 13872 18164
rect 13726 18119 13782 18128
rect 13832 18086 13860 18158
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13740 17338 13768 18022
rect 13832 17338 13860 18022
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13832 16454 13860 17274
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13924 14958 13952 18838
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12442 13860 12786
rect 13820 12436 13872 12442
rect 14016 12434 14044 20046
rect 14108 19514 14136 22066
rect 14280 22034 14332 22040
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14660 21962 14688 23258
rect 14936 22930 14964 29294
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 15028 24818 15056 27270
rect 15212 26314 15240 30262
rect 15304 29102 15332 30631
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15304 28422 15332 29038
rect 15292 28416 15344 28422
rect 15290 28384 15292 28393
rect 15344 28384 15346 28393
rect 15290 28319 15346 28328
rect 15396 27878 15424 31726
rect 15488 31210 15516 32796
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15580 28558 15608 29174
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15384 26376 15436 26382
rect 15384 26318 15436 26324
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15396 26042 15424 26318
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15396 25752 15424 25978
rect 15488 25922 15516 27406
rect 15580 26042 15608 27814
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15488 25894 15608 25922
rect 15476 25764 15528 25770
rect 15396 25724 15476 25752
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 15120 24682 15148 25094
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 14936 22902 15056 22930
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14200 21486 14228 21898
rect 14646 21720 14702 21729
rect 14646 21655 14702 21664
rect 14660 21486 14688 21655
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14292 20058 14320 20470
rect 14660 20330 14688 21422
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14108 18358 14136 19450
rect 14200 18970 14228 19722
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14660 19174 14688 19314
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 14108 17610 14136 18294
rect 14096 17604 14148 17610
rect 14096 17546 14148 17552
rect 14384 17134 14412 18770
rect 14660 17542 14688 19110
rect 14752 17678 14780 22374
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 14832 19712 14884 19718
rect 14830 19680 14832 19689
rect 14884 19680 14886 19689
rect 14830 19615 14886 19624
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14844 18834 14872 19178
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14844 17746 14872 18770
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 13820 12378 13872 12384
rect 13924 12406 14044 12434
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13096 870 13216 898
rect 13096 800 13124 870
rect 3252 734 3464 762
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13188 762 13216 870
rect 13372 762 13400 2926
rect 13464 800 13492 4014
rect 13648 3126 13676 12174
rect 13924 8430 13952 12406
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 14108 6914 14136 15846
rect 14292 15706 14320 16662
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14384 15570 14412 17070
rect 14660 17066 14688 17478
rect 14844 17202 14872 17682
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14738 16280 14794 16289
rect 14738 16215 14740 16224
rect 14792 16215 14794 16224
rect 14740 16186 14792 16192
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14844 15450 14872 17138
rect 14752 15422 14872 15450
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14550 14596 14962
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14752 14482 14780 15422
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14108 6886 14228 6914
rect 14200 4486 14228 6886
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 14292 3058 14320 12650
rect 14384 11354 14412 13194
rect 14476 12442 14504 13262
rect 14844 13258 14872 14894
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14568 11898 14596 13194
rect 14936 12986 14964 22034
rect 15028 20942 15056 22902
rect 15212 22778 15240 25638
rect 15396 25362 15424 25724
rect 15476 25706 15528 25712
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15396 24970 15424 25298
rect 15304 24942 15424 24970
rect 15304 23186 15332 24942
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 13832 800 13860 2314
rect 14200 800 14228 2926
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14568 800 14596 2450
rect 14660 2446 14688 12650
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11218 14780 11698
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14844 10674 14872 12718
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15120 3670 15148 16594
rect 15212 12918 15240 22578
rect 15304 19417 15332 22714
rect 15396 21690 15424 24346
rect 15580 22778 15608 25894
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15672 22094 15700 38898
rect 15764 37398 15792 39918
rect 15752 37392 15804 37398
rect 15752 37334 15804 37340
rect 15856 36922 15884 40530
rect 15948 40458 15976 41386
rect 16132 41274 16160 41534
rect 16212 41472 16264 41478
rect 16212 41414 16264 41420
rect 16120 41268 16172 41274
rect 16120 41210 16172 41216
rect 15936 40452 15988 40458
rect 15936 40394 15988 40400
rect 15948 40089 15976 40394
rect 15934 40080 15990 40089
rect 15934 40015 15990 40024
rect 16028 39976 16080 39982
rect 16028 39918 16080 39924
rect 16120 39976 16172 39982
rect 16120 39918 16172 39924
rect 16040 39574 16068 39918
rect 16132 39642 16160 39918
rect 16120 39636 16172 39642
rect 16120 39578 16172 39584
rect 16028 39568 16080 39574
rect 16028 39510 16080 39516
rect 16040 39386 16068 39510
rect 15948 39358 16068 39386
rect 15948 39098 15976 39358
rect 16028 39296 16080 39302
rect 16028 39238 16080 39244
rect 16040 39098 16068 39238
rect 15936 39092 15988 39098
rect 15936 39034 15988 39040
rect 16028 39092 16080 39098
rect 16028 39034 16080 39040
rect 15936 38344 15988 38350
rect 15936 38286 15988 38292
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 15844 36712 15896 36718
rect 15842 36680 15844 36689
rect 15896 36680 15898 36689
rect 15842 36615 15898 36624
rect 15750 36272 15806 36281
rect 15750 36207 15752 36216
rect 15804 36207 15806 36216
rect 15752 36178 15804 36184
rect 15948 35494 15976 38286
rect 16120 37800 16172 37806
rect 16120 37742 16172 37748
rect 16028 36644 16080 36650
rect 16028 36586 16080 36592
rect 15936 35488 15988 35494
rect 15936 35430 15988 35436
rect 15948 35170 15976 35430
rect 15764 35154 15976 35170
rect 15752 35148 15976 35154
rect 15804 35142 15976 35148
rect 15752 35090 15804 35096
rect 15752 34672 15804 34678
rect 15752 34614 15804 34620
rect 15764 30122 15792 34614
rect 15844 34468 15896 34474
rect 15844 34410 15896 34416
rect 15856 33318 15884 34410
rect 15948 34066 15976 35142
rect 15936 34060 15988 34066
rect 15936 34002 15988 34008
rect 15948 33658 15976 34002
rect 15936 33652 15988 33658
rect 15936 33594 15988 33600
rect 15844 33312 15896 33318
rect 15844 33254 15896 33260
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 15856 31754 15884 32846
rect 15936 32292 15988 32298
rect 15936 32234 15988 32240
rect 15948 31958 15976 32234
rect 15936 31952 15988 31958
rect 15936 31894 15988 31900
rect 15856 31726 15976 31754
rect 15752 30116 15804 30122
rect 15752 30058 15804 30064
rect 15764 28966 15792 30058
rect 15752 28960 15804 28966
rect 15752 28902 15804 28908
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15488 22066 15700 22094
rect 15488 21894 15516 22066
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15290 19408 15346 19417
rect 15290 19343 15346 19352
rect 15396 18222 15424 21422
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 15502 15332 16390
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15488 15026 15516 21830
rect 15764 20942 15792 28358
rect 15842 28248 15898 28257
rect 15842 28183 15844 28192
rect 15896 28183 15898 28192
rect 15844 28154 15896 28160
rect 15856 22710 15884 28154
rect 15948 24410 15976 31726
rect 16040 29850 16068 36586
rect 16132 35290 16160 37742
rect 16224 37330 16252 41414
rect 16304 40112 16356 40118
rect 16304 40054 16356 40060
rect 16316 39846 16344 40054
rect 16304 39840 16356 39846
rect 16304 39782 16356 39788
rect 16316 38010 16344 39782
rect 16408 38894 16436 43590
rect 16592 41682 16620 47398
rect 16672 47116 16724 47122
rect 16724 47076 16804 47104
rect 16672 47058 16724 47064
rect 16776 46510 16804 47076
rect 17408 46912 17460 46918
rect 17408 46854 17460 46860
rect 17420 46646 17448 46854
rect 17408 46640 17460 46646
rect 17408 46582 17460 46588
rect 16764 46504 16816 46510
rect 16764 46446 16816 46452
rect 16672 46368 16724 46374
rect 16672 46310 16724 46316
rect 16684 45082 16712 46310
rect 16672 45076 16724 45082
rect 16672 45018 16724 45024
rect 16776 44946 16804 46446
rect 17420 46170 17448 46582
rect 17408 46164 17460 46170
rect 17408 46106 17460 46112
rect 16948 45076 17000 45082
rect 16948 45018 17000 45024
rect 16764 44940 16816 44946
rect 16764 44882 16816 44888
rect 16776 44334 16804 44882
rect 16672 44328 16724 44334
rect 16672 44270 16724 44276
rect 16764 44328 16816 44334
rect 16764 44270 16816 44276
rect 16684 42226 16712 44270
rect 16776 43178 16804 44270
rect 16856 43920 16908 43926
rect 16856 43862 16908 43868
rect 16764 43172 16816 43178
rect 16764 43114 16816 43120
rect 16776 42770 16804 43114
rect 16764 42764 16816 42770
rect 16764 42706 16816 42712
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 16580 41676 16632 41682
rect 16580 41618 16632 41624
rect 16670 41576 16726 41585
rect 16670 41511 16726 41520
rect 16488 41472 16540 41478
rect 16488 41414 16540 41420
rect 16396 38888 16448 38894
rect 16396 38830 16448 38836
rect 16304 38004 16356 38010
rect 16304 37946 16356 37952
rect 16316 37670 16344 37946
rect 16394 37768 16450 37777
rect 16394 37703 16396 37712
rect 16448 37703 16450 37712
rect 16396 37674 16448 37680
rect 16304 37664 16356 37670
rect 16356 37612 16436 37618
rect 16304 37606 16436 37612
rect 16316 37590 16436 37606
rect 16212 37324 16264 37330
rect 16212 37266 16264 37272
rect 16120 35284 16172 35290
rect 16120 35226 16172 35232
rect 16120 35148 16172 35154
rect 16120 35090 16172 35096
rect 16132 35018 16160 35090
rect 16120 35012 16172 35018
rect 16120 34954 16172 34960
rect 16132 33862 16160 34954
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 16132 33318 16160 33798
rect 16408 33318 16436 37590
rect 16500 36242 16528 41414
rect 16684 41138 16712 41511
rect 16672 41132 16724 41138
rect 16672 41074 16724 41080
rect 16776 41070 16804 42502
rect 16764 41064 16816 41070
rect 16764 41006 16816 41012
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 16488 36236 16540 36242
rect 16488 36178 16540 36184
rect 16120 33312 16172 33318
rect 16118 33280 16120 33289
rect 16396 33312 16448 33318
rect 16172 33280 16174 33289
rect 16396 33254 16448 33260
rect 16118 33215 16174 33224
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 16488 32972 16540 32978
rect 16488 32914 16540 32920
rect 16408 32774 16436 32914
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16132 32570 16160 32710
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16120 31952 16172 31958
rect 16120 31894 16172 31900
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16132 29306 16160 31894
rect 16500 30802 16528 32914
rect 16592 31754 16620 40462
rect 16868 38978 16896 43862
rect 16960 40662 16988 45018
rect 17132 44736 17184 44742
rect 17132 44678 17184 44684
rect 17144 44470 17172 44678
rect 17132 44464 17184 44470
rect 17132 44406 17184 44412
rect 17408 43648 17460 43654
rect 17408 43590 17460 43596
rect 17420 43450 17448 43590
rect 17512 43450 17540 47398
rect 17408 43444 17460 43450
rect 17408 43386 17460 43392
rect 17500 43444 17552 43450
rect 17500 43386 17552 43392
rect 17040 43104 17092 43110
rect 17040 43046 17092 43052
rect 16948 40656 17000 40662
rect 16948 40598 17000 40604
rect 17052 40594 17080 43046
rect 17408 42288 17460 42294
rect 17408 42230 17460 42236
rect 17316 40656 17368 40662
rect 17316 40598 17368 40604
rect 17040 40588 17092 40594
rect 17040 40530 17092 40536
rect 17040 40384 17092 40390
rect 17040 40326 17092 40332
rect 17052 39370 17080 40326
rect 17132 39908 17184 39914
rect 17132 39850 17184 39856
rect 17040 39364 17092 39370
rect 17040 39306 17092 39312
rect 16776 38950 16896 38978
rect 16670 36816 16726 36825
rect 16670 36751 16672 36760
rect 16724 36751 16726 36760
rect 16672 36722 16724 36728
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16684 33454 16712 35158
rect 16672 33448 16724 33454
rect 16672 33390 16724 33396
rect 16684 32366 16712 33390
rect 16776 32910 16804 38950
rect 17038 37904 17094 37913
rect 17038 37839 17094 37848
rect 17052 37398 17080 37839
rect 17040 37392 17092 37398
rect 17040 37334 17092 37340
rect 16948 36916 17000 36922
rect 16948 36858 17000 36864
rect 16960 36242 16988 36858
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 17144 35834 17172 39850
rect 17224 39364 17276 39370
rect 17224 39306 17276 39312
rect 17236 39030 17264 39306
rect 17224 39024 17276 39030
rect 17224 38966 17276 38972
rect 17224 38888 17276 38894
rect 17224 38830 17276 38836
rect 17236 38010 17264 38830
rect 17224 38004 17276 38010
rect 17224 37946 17276 37952
rect 17328 36718 17356 40598
rect 17420 38554 17448 42230
rect 17500 40452 17552 40458
rect 17500 40394 17552 40400
rect 17408 38548 17460 38554
rect 17408 38490 17460 38496
rect 17406 38040 17462 38049
rect 17406 37975 17462 37984
rect 17420 37738 17448 37975
rect 17408 37732 17460 37738
rect 17408 37674 17460 37680
rect 17316 36712 17368 36718
rect 17316 36654 17368 36660
rect 17224 36576 17276 36582
rect 17224 36518 17276 36524
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 16856 33312 16908 33318
rect 16856 33254 16908 33260
rect 17130 33280 17186 33289
rect 16868 32978 16896 33254
rect 17130 33215 17186 33224
rect 17144 33046 17172 33215
rect 17040 33040 17092 33046
rect 17040 32982 17092 32988
rect 17132 33040 17184 33046
rect 17132 32982 17184 32988
rect 16856 32972 16908 32978
rect 16856 32914 16908 32920
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16960 31754 16988 32166
rect 16592 31726 16712 31754
rect 16488 30796 16540 30802
rect 16488 30738 16540 30744
rect 16580 30660 16632 30666
rect 16580 30602 16632 30608
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16028 29028 16080 29034
rect 16028 28970 16080 28976
rect 16040 28558 16068 28970
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 16028 28008 16080 28014
rect 16026 27976 16028 27985
rect 16080 27976 16082 27985
rect 16026 27911 16082 27920
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16040 23322 16068 25774
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15948 22574 15976 22986
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 15948 22094 15976 22510
rect 16028 22094 16080 22098
rect 15948 22092 16080 22094
rect 15948 22066 16028 22092
rect 16132 22094 16160 29106
rect 16224 28626 16252 30126
rect 16592 29850 16620 30602
rect 16488 29844 16540 29850
rect 16488 29786 16540 29792
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16394 29744 16450 29753
rect 16394 29679 16450 29688
rect 16408 29646 16436 29679
rect 16396 29640 16448 29646
rect 16396 29582 16448 29588
rect 16408 29102 16436 29582
rect 16396 29096 16448 29102
rect 16394 29064 16396 29073
rect 16448 29064 16450 29073
rect 16394 28999 16450 29008
rect 16212 28620 16264 28626
rect 16212 28562 16264 28568
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16224 22982 16252 27950
rect 16396 27328 16448 27334
rect 16396 27270 16448 27276
rect 16408 27062 16436 27270
rect 16396 27056 16448 27062
rect 16316 27004 16396 27010
rect 16316 26998 16448 27004
rect 16316 26982 16436 26998
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16224 22778 16252 22918
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16132 22066 16252 22094
rect 16028 22034 16080 22040
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15580 17814 15608 20742
rect 16040 19922 16068 21286
rect 16132 21078 16160 21490
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16224 18850 16252 22066
rect 16316 18952 16344 26982
rect 16396 24880 16448 24886
rect 16396 24822 16448 24828
rect 16408 24614 16436 24822
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16408 24313 16436 24550
rect 16394 24304 16450 24313
rect 16394 24239 16450 24248
rect 16500 23594 16528 29786
rect 16684 29782 16712 31726
rect 16868 31726 16988 31754
rect 16672 29776 16724 29782
rect 16672 29718 16724 29724
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16592 27130 16620 29446
rect 16684 29102 16712 29718
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16776 28762 16804 29514
rect 16764 28756 16816 28762
rect 16764 28698 16816 28704
rect 16868 28558 16896 31726
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16948 28416 17000 28422
rect 16948 28358 17000 28364
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 25362 16712 26522
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16776 24206 16804 25434
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16868 24954 16896 25094
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16854 24712 16910 24721
rect 16854 24647 16910 24656
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16672 24064 16724 24070
rect 16868 24052 16896 24647
rect 16960 24274 16988 28358
rect 17052 27470 17080 32982
rect 17236 32502 17264 36518
rect 17512 32910 17540 40394
rect 17604 38729 17632 47602
rect 18420 47524 18472 47530
rect 18420 47466 18472 47472
rect 18432 47258 18460 47466
rect 18420 47252 18472 47258
rect 18420 47194 18472 47200
rect 17684 47116 17736 47122
rect 17684 47058 17736 47064
rect 17696 45014 17724 47058
rect 18328 46980 18380 46986
rect 18328 46922 18380 46928
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 18340 46594 18368 46922
rect 18432 46714 18460 47194
rect 18512 47184 18564 47190
rect 18512 47126 18564 47132
rect 18420 46708 18472 46714
rect 18420 46650 18472 46656
rect 18340 46566 18460 46594
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 17684 45008 17736 45014
rect 17684 44950 17736 44956
rect 17696 43246 17724 44950
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 18340 43246 18368 45358
rect 18432 43994 18460 46566
rect 18420 43988 18472 43994
rect 18420 43930 18472 43936
rect 18420 43852 18472 43858
rect 18420 43794 18472 43800
rect 17684 43240 17736 43246
rect 17684 43182 17736 43188
rect 18328 43240 18380 43246
rect 18328 43182 18380 43188
rect 18432 42770 18460 43794
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17776 41744 17828 41750
rect 17776 41686 17828 41692
rect 17684 39500 17736 39506
rect 17684 39442 17736 39448
rect 17590 38720 17646 38729
rect 17590 38655 17646 38664
rect 17590 38448 17646 38457
rect 17590 38383 17646 38392
rect 17604 38350 17632 38383
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 17604 38010 17632 38286
rect 17696 38214 17724 39442
rect 17684 38208 17736 38214
rect 17684 38150 17736 38156
rect 17592 38004 17644 38010
rect 17592 37946 17644 37952
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17224 32496 17276 32502
rect 17224 32438 17276 32444
rect 17132 32292 17184 32298
rect 17132 32234 17184 32240
rect 17144 31822 17172 32234
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17144 28626 17172 31078
rect 17500 30728 17552 30734
rect 17420 30688 17500 30716
rect 17420 30598 17448 30688
rect 17500 30670 17552 30676
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17236 29306 17264 30126
rect 17512 30054 17540 30534
rect 17604 30326 17632 37130
rect 17696 35834 17724 38150
rect 17788 37806 17816 41686
rect 18524 41682 18552 47126
rect 18616 47122 18644 52838
rect 19064 49088 19116 49094
rect 19064 49030 19116 49036
rect 18696 47660 18748 47666
rect 18696 47602 18748 47608
rect 18604 47116 18656 47122
rect 18604 47058 18656 47064
rect 18604 46504 18656 46510
rect 18604 46446 18656 46452
rect 18616 44538 18644 46446
rect 18604 44532 18656 44538
rect 18604 44474 18656 44480
rect 18604 42696 18656 42702
rect 18604 42638 18656 42644
rect 18512 41676 18564 41682
rect 18512 41618 18564 41624
rect 18420 41472 18472 41478
rect 18420 41414 18472 41420
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 18328 40996 18380 41002
rect 18328 40938 18380 40944
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 18236 40180 18288 40186
rect 18236 40122 18288 40128
rect 18248 40089 18276 40122
rect 18340 40118 18368 40938
rect 18432 40186 18460 41414
rect 18512 40928 18564 40934
rect 18512 40870 18564 40876
rect 18420 40180 18472 40186
rect 18420 40122 18472 40128
rect 18328 40112 18380 40118
rect 18234 40080 18290 40089
rect 18328 40054 18380 40060
rect 18234 40015 18290 40024
rect 18420 40044 18472 40050
rect 18420 39986 18472 39992
rect 18432 39386 18460 39986
rect 18340 39358 18460 39386
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17866 38992 17922 39001
rect 17866 38927 17922 38936
rect 17880 38486 17908 38927
rect 18236 38820 18288 38826
rect 18236 38762 18288 38768
rect 17868 38480 17920 38486
rect 17868 38422 17920 38428
rect 18248 38418 18276 38762
rect 18236 38412 18288 38418
rect 18236 38354 18288 38360
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17868 37936 17920 37942
rect 17868 37878 17920 37884
rect 18236 37936 18288 37942
rect 18236 37878 18288 37884
rect 17776 37800 17828 37806
rect 17776 37742 17828 37748
rect 17880 37330 17908 37878
rect 18248 37482 18276 37878
rect 18340 37670 18368 39358
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38894 18460 39238
rect 18420 38888 18472 38894
rect 18418 38856 18420 38865
rect 18472 38856 18474 38865
rect 18418 38791 18474 38800
rect 18524 38758 18552 40870
rect 18616 39642 18644 42638
rect 18604 39636 18656 39642
rect 18604 39578 18656 39584
rect 18616 39030 18644 39578
rect 18708 39302 18736 47602
rect 18972 46708 19024 46714
rect 18972 46650 19024 46656
rect 18880 45280 18932 45286
rect 18880 45222 18932 45228
rect 18788 44532 18840 44538
rect 18788 44474 18840 44480
rect 18800 39982 18828 44474
rect 18788 39976 18840 39982
rect 18788 39918 18840 39924
rect 18788 39364 18840 39370
rect 18788 39306 18840 39312
rect 18696 39296 18748 39302
rect 18696 39238 18748 39244
rect 18604 39024 18656 39030
rect 18604 38966 18656 38972
rect 18420 38752 18472 38758
rect 18420 38694 18472 38700
rect 18512 38752 18564 38758
rect 18512 38694 18564 38700
rect 18604 38752 18656 38758
rect 18604 38694 18656 38700
rect 18328 37664 18380 37670
rect 18328 37606 18380 37612
rect 17972 37454 18276 37482
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17972 37210 18000 37454
rect 17788 37182 18000 37210
rect 17684 35828 17736 35834
rect 17684 35770 17736 35776
rect 17788 35766 17816 37182
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17776 35760 17828 35766
rect 17776 35702 17828 35708
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33590 18368 35430
rect 18432 34678 18460 38694
rect 18616 38026 18644 38694
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 18524 37998 18644 38026
rect 18708 38010 18736 38354
rect 18696 38004 18748 38010
rect 18524 37330 18552 37998
rect 18696 37946 18748 37952
rect 18604 37868 18656 37874
rect 18604 37810 18656 37816
rect 18616 37670 18644 37810
rect 18604 37664 18656 37670
rect 18604 37606 18656 37612
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 18512 37120 18564 37126
rect 18512 37062 18564 37068
rect 18524 36922 18552 37062
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 18616 35714 18644 37606
rect 18708 37466 18736 37946
rect 18696 37460 18748 37466
rect 18696 37402 18748 37408
rect 18696 37324 18748 37330
rect 18696 37266 18748 37272
rect 18524 35686 18644 35714
rect 18420 34672 18472 34678
rect 18420 34614 18472 34620
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 18326 33144 18382 33153
rect 18326 33079 18382 33088
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17776 32360 17828 32366
rect 17776 32302 17828 32308
rect 17684 31680 17736 31686
rect 17684 31622 17736 31628
rect 17592 30320 17644 30326
rect 17592 30262 17644 30268
rect 17500 30048 17552 30054
rect 17420 29996 17500 30002
rect 17420 29990 17552 29996
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17420 29974 17540 29990
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24274 17080 25094
rect 17144 24886 17172 27474
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 16672 24006 16724 24012
rect 16776 24024 16896 24052
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23474 16528 23530
rect 16500 23446 16620 23474
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16408 22982 16436 23054
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22710 16436 22918
rect 16592 22778 16620 23446
rect 16488 22772 16540 22778
rect 16488 22714 16540 22720
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16408 22234 16436 22646
rect 16396 22228 16448 22234
rect 16396 22170 16448 22176
rect 16408 21962 16436 22170
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21146 16436 21286
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16316 18924 16436 18952
rect 16224 18822 16344 18850
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18222 16252 18702
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15304 12434 15332 13942
rect 15396 13394 15424 14418
rect 15580 14278 15608 17478
rect 15750 16824 15806 16833
rect 15750 16759 15806 16768
rect 15764 16454 15792 16759
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15672 12442 15700 15302
rect 15212 12406 15332 12434
rect 15660 12436 15712 12442
rect 15212 11898 15240 12406
rect 15660 12378 15712 12384
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14936 800 14964 3538
rect 15396 2650 15424 12038
rect 15764 11642 15792 15846
rect 15856 12238 15884 17818
rect 16040 16658 16068 18158
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16132 17490 16160 17750
rect 16316 17746 16344 18822
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16132 17462 16344 17490
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15934 16280 15990 16289
rect 15934 16215 15990 16224
rect 15948 16182 15976 16215
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 13530 15976 14282
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15948 12850 15976 13466
rect 16040 13025 16068 16594
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16026 13016 16082 13025
rect 16132 12986 16160 13262
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16026 12951 16082 12960
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16132 12866 16160 12922
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 16040 12838 16160 12866
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15948 11914 15976 12242
rect 16040 12102 16068 12838
rect 16224 12730 16252 13194
rect 16132 12702 16252 12730
rect 16316 12730 16344 17462
rect 16408 15502 16436 18924
rect 16500 18834 16528 22714
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16500 16096 16528 18158
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17338 16620 17478
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17202 16712 24006
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 16108 16632 16114
rect 16500 16068 16580 16096
rect 16580 16050 16632 16056
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 14958 16436 15438
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16592 14498 16620 16050
rect 16776 15434 16804 24024
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16868 21894 16896 22034
rect 17052 22030 17080 23598
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 17144 21146 17172 24822
rect 17328 24818 17356 29786
rect 17420 29102 17448 29974
rect 17604 29782 17632 29990
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17500 29504 17552 29510
rect 17500 29446 17552 29452
rect 17512 29306 17540 29446
rect 17604 29306 17632 29514
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17592 29028 17644 29034
rect 17592 28970 17644 28976
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17512 27878 17540 28018
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17328 24274 17356 24754
rect 17316 24268 17368 24274
rect 17316 24210 17368 24216
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17144 21010 17172 21082
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16408 14482 16620 14498
rect 16396 14476 16620 14482
rect 16448 14470 16620 14476
rect 16396 14418 16448 14424
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16408 12866 16436 14214
rect 16500 13258 16528 14214
rect 16592 13938 16620 14470
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16500 12986 16528 13194
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16408 12838 16528 12866
rect 16316 12702 16436 12730
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 15948 11886 16068 11914
rect 16132 11898 16160 12702
rect 16304 12640 16356 12646
rect 16210 12608 16266 12617
rect 16304 12582 16356 12588
rect 16210 12543 16266 12552
rect 16224 12306 16252 12543
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 15580 11614 15792 11642
rect 15580 3534 15608 11614
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 10674 15792 11494
rect 16040 11218 16068 11886
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 11014 15976 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15948 10538 15976 10950
rect 16040 10742 16068 11154
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15948 3942 15976 10474
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15304 800 15332 2450
rect 15672 800 15700 2926
rect 16040 800 16068 3538
rect 16316 3534 16344 12582
rect 16408 9654 16436 12702
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16500 6914 16528 12838
rect 16408 6886 16528 6914
rect 16408 6798 16436 6886
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16684 4146 16712 14826
rect 16868 12170 16896 16934
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16960 14550 16988 16390
rect 17144 16182 17172 17682
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17052 15094 17080 15302
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17144 14618 17172 16118
rect 17236 15094 17264 21626
rect 17420 21554 17448 26794
rect 17500 26512 17552 26518
rect 17500 26454 17552 26460
rect 17512 24750 17540 26454
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17512 24070 17540 24686
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17512 23526 17540 24006
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17314 20632 17370 20641
rect 17314 20567 17316 20576
rect 17368 20567 17370 20576
rect 17316 20538 17368 20544
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17328 15910 17356 19450
rect 17512 18358 17540 22714
rect 17604 22094 17632 28970
rect 17696 24954 17724 31622
rect 17788 30598 17816 32302
rect 17960 32224 18012 32230
rect 18012 32184 18092 32212
rect 17960 32166 18012 32172
rect 17960 32020 18012 32026
rect 17960 31962 18012 31968
rect 17972 31754 18000 31962
rect 18064 31822 18092 32184
rect 18340 31906 18368 33079
rect 18432 32026 18460 34002
rect 18420 32020 18472 32026
rect 18420 31962 18472 31968
rect 18248 31890 18368 31906
rect 18236 31884 18368 31890
rect 18288 31878 18368 31884
rect 18236 31826 18288 31832
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17880 31726 18000 31754
rect 17880 31278 17908 31726
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18340 31346 18368 31878
rect 18420 31408 18472 31414
rect 18420 31350 18472 31356
rect 18328 31340 18380 31346
rect 18328 31282 18380 31288
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 26586 17816 28562
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17880 26518 17908 31214
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18340 30394 18368 31282
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18052 30184 18104 30190
rect 18052 30126 18104 30132
rect 18064 30054 18092 30126
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 18340 29034 18368 29446
rect 18052 29028 18104 29034
rect 18052 28970 18104 28976
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 18064 28665 18092 28970
rect 18432 28966 18460 31350
rect 18524 30938 18552 35686
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18616 32366 18644 32710
rect 18708 32450 18736 37266
rect 18800 36854 18828 39306
rect 18788 36848 18840 36854
rect 18788 36790 18840 36796
rect 18788 36712 18840 36718
rect 18788 36654 18840 36660
rect 18800 34678 18828 36654
rect 18892 35578 18920 45222
rect 18984 44334 19012 46650
rect 18972 44328 19024 44334
rect 18972 44270 19024 44276
rect 18984 41682 19012 44270
rect 19076 42702 19104 49030
rect 19352 47274 19380 53926
rect 19616 53440 19668 53446
rect 19616 53382 19668 53388
rect 19260 47246 19380 47274
rect 19260 46986 19288 47246
rect 19340 47116 19392 47122
rect 19340 47058 19392 47064
rect 19248 46980 19300 46986
rect 19248 46922 19300 46928
rect 19248 46640 19300 46646
rect 19168 46600 19248 46628
rect 19168 46170 19196 46600
rect 19248 46582 19300 46588
rect 19352 46510 19380 47058
rect 19340 46504 19392 46510
rect 19340 46446 19392 46452
rect 19156 46164 19208 46170
rect 19156 46106 19208 46112
rect 19168 45558 19196 46106
rect 19352 45626 19380 46446
rect 19524 46368 19576 46374
rect 19524 46310 19576 46316
rect 19340 45620 19392 45626
rect 19340 45562 19392 45568
rect 19156 45552 19208 45558
rect 19156 45494 19208 45500
rect 19536 44878 19564 46310
rect 19628 45898 19656 53382
rect 19720 53242 19748 54062
rect 19904 53582 19932 56200
rect 19892 53576 19944 53582
rect 19892 53518 19944 53524
rect 19708 53236 19760 53242
rect 19708 53178 19760 53184
rect 20272 53106 20300 56200
rect 20640 55214 20668 56200
rect 20640 55186 20760 55214
rect 20732 54194 20760 55186
rect 20720 54188 20772 54194
rect 20720 54130 20772 54136
rect 20628 53508 20680 53514
rect 20628 53450 20680 53456
rect 20260 53100 20312 53106
rect 20260 53042 20312 53048
rect 20168 52896 20220 52902
rect 20168 52838 20220 52844
rect 20180 46034 20208 52838
rect 20536 48000 20588 48006
rect 20536 47942 20588 47948
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 20444 46028 20496 46034
rect 20444 45970 20496 45976
rect 19616 45892 19668 45898
rect 19616 45834 19668 45840
rect 19892 45824 19944 45830
rect 20076 45824 20128 45830
rect 19892 45766 19944 45772
rect 20074 45792 20076 45801
rect 20128 45792 20130 45801
rect 19524 44872 19576 44878
rect 19524 44814 19576 44820
rect 19536 44334 19564 44814
rect 19800 44804 19852 44810
rect 19800 44746 19852 44752
rect 19812 44538 19840 44746
rect 19800 44532 19852 44538
rect 19800 44474 19852 44480
rect 19524 44328 19576 44334
rect 19524 44270 19576 44276
rect 19340 43648 19392 43654
rect 19340 43590 19392 43596
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 19064 42696 19116 42702
rect 19064 42638 19116 42644
rect 19260 42158 19288 43046
rect 19064 42152 19116 42158
rect 19064 42094 19116 42100
rect 19248 42152 19300 42158
rect 19248 42094 19300 42100
rect 18972 41676 19024 41682
rect 18972 41618 19024 41624
rect 18972 40996 19024 41002
rect 18972 40938 19024 40944
rect 18984 38758 19012 40938
rect 19076 40066 19104 42094
rect 19260 41614 19288 42094
rect 19248 41608 19300 41614
rect 19246 41576 19248 41585
rect 19300 41576 19302 41585
rect 19156 41540 19208 41546
rect 19246 41511 19302 41520
rect 19156 41482 19208 41488
rect 19168 40934 19196 41482
rect 19156 40928 19208 40934
rect 19156 40870 19208 40876
rect 19168 40526 19196 40870
rect 19156 40520 19208 40526
rect 19156 40462 19208 40468
rect 19076 40038 19288 40066
rect 19064 39908 19116 39914
rect 19064 39850 19116 39856
rect 19076 39642 19104 39850
rect 19064 39636 19116 39642
rect 19064 39578 19116 39584
rect 18972 38752 19024 38758
rect 18972 38694 19024 38700
rect 18972 38344 19024 38350
rect 18972 38286 19024 38292
rect 18984 36310 19012 38286
rect 19076 38214 19104 39578
rect 19156 38888 19208 38894
rect 19156 38830 19208 38836
rect 19064 38208 19116 38214
rect 19064 38150 19116 38156
rect 18972 36304 19024 36310
rect 18972 36246 19024 36252
rect 18892 35550 19012 35578
rect 18788 34672 18840 34678
rect 18788 34614 18840 34620
rect 18708 32434 18920 32450
rect 18708 32428 18932 32434
rect 18708 32422 18880 32428
rect 18880 32370 18932 32376
rect 18604 32360 18656 32366
rect 18656 32320 18828 32348
rect 18604 32302 18656 32308
rect 18696 32224 18748 32230
rect 18696 32166 18748 32172
rect 18604 31476 18656 31482
rect 18604 31418 18656 31424
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18616 30818 18644 31418
rect 18524 30790 18644 30818
rect 18524 30054 18552 30790
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18512 30048 18564 30054
rect 18512 29990 18564 29996
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18420 28688 18472 28694
rect 18050 28656 18106 28665
rect 18420 28630 18472 28636
rect 18050 28591 18106 28600
rect 18064 28490 18092 28591
rect 18326 28520 18382 28529
rect 18052 28484 18104 28490
rect 18326 28455 18382 28464
rect 18052 28426 18104 28432
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 18340 28218 18368 28455
rect 18432 28422 18460 28630
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18328 28212 18380 28218
rect 18328 28154 18380 28160
rect 18340 27674 18368 28154
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 18234 27568 18290 27577
rect 18234 27503 18290 27512
rect 18248 27402 18276 27503
rect 18236 27396 18288 27402
rect 18236 27338 18288 27344
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18156 26926 18184 26998
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18340 26874 18368 27610
rect 18432 27062 18460 28358
rect 18420 27056 18472 27062
rect 18420 26998 18472 27004
rect 18340 26846 18460 26874
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 17868 26512 17920 26518
rect 17868 26454 17920 26460
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17788 25498 17816 26250
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17788 25226 17816 25434
rect 17776 25220 17828 25226
rect 17776 25162 17828 25168
rect 17880 25158 17908 25774
rect 18248 25498 18276 25774
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18340 25158 18368 26726
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17684 24948 17736 24954
rect 17684 24890 17736 24896
rect 18340 24818 18368 25094
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17788 22098 17816 24686
rect 17880 22506 17908 24754
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 17604 22066 17724 22094
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17604 20942 17632 21422
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19446 17632 19722
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17696 19310 17724 22066
rect 17776 22092 17828 22098
rect 18432 22094 18460 26846
rect 18524 25158 18552 29990
rect 18616 28014 18644 30534
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18616 27441 18644 27950
rect 18602 27432 18658 27441
rect 18602 27367 18658 27376
rect 18604 27328 18656 27334
rect 18604 27270 18656 27276
rect 18616 26081 18644 27270
rect 18602 26072 18658 26081
rect 18708 26042 18736 32166
rect 18800 31414 18828 32320
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18788 31408 18840 31414
rect 18788 31350 18840 31356
rect 18892 31278 18920 31758
rect 18984 31482 19012 35550
rect 19076 35290 19104 38150
rect 19168 35816 19196 38830
rect 19260 38418 19288 40038
rect 19352 39982 19380 43590
rect 19616 43240 19668 43246
rect 19616 43182 19668 43188
rect 19628 41070 19656 43182
rect 19708 42084 19760 42090
rect 19708 42026 19760 42032
rect 19720 41682 19748 42026
rect 19708 41676 19760 41682
rect 19708 41618 19760 41624
rect 19904 41274 19932 45766
rect 20074 45727 20130 45736
rect 20076 45416 20128 45422
rect 20076 45358 20128 45364
rect 20260 45416 20312 45422
rect 20260 45358 20312 45364
rect 20088 43450 20116 45358
rect 20272 44810 20300 45358
rect 20260 44804 20312 44810
rect 20260 44746 20312 44752
rect 20272 44470 20300 44746
rect 20456 44538 20484 45970
rect 20444 44532 20496 44538
rect 20444 44474 20496 44480
rect 20260 44464 20312 44470
rect 20260 44406 20312 44412
rect 20076 43444 20128 43450
rect 20076 43386 20128 43392
rect 19984 41472 20036 41478
rect 19984 41414 20036 41420
rect 19892 41268 19944 41274
rect 19892 41210 19944 41216
rect 19800 41132 19852 41138
rect 19800 41074 19852 41080
rect 19616 41064 19668 41070
rect 19616 41006 19668 41012
rect 19432 40928 19484 40934
rect 19432 40870 19484 40876
rect 19524 40928 19576 40934
rect 19524 40870 19576 40876
rect 19340 39976 19392 39982
rect 19340 39918 19392 39924
rect 19444 39506 19472 40870
rect 19536 40730 19564 40870
rect 19628 40730 19656 41006
rect 19524 40724 19576 40730
rect 19524 40666 19576 40672
rect 19616 40724 19668 40730
rect 19616 40666 19668 40672
rect 19616 40588 19668 40594
rect 19616 40530 19668 40536
rect 19432 39500 19484 39506
rect 19432 39442 19484 39448
rect 19248 38412 19300 38418
rect 19248 38354 19300 38360
rect 19260 37942 19288 38354
rect 19524 38276 19576 38282
rect 19524 38218 19576 38224
rect 19248 37936 19300 37942
rect 19248 37878 19300 37884
rect 19294 37664 19346 37670
rect 19260 37612 19294 37618
rect 19260 37606 19346 37612
rect 19260 37590 19334 37606
rect 19260 37505 19288 37590
rect 19246 37496 19302 37505
rect 19246 37431 19302 37440
rect 19248 37324 19300 37330
rect 19248 37266 19300 37272
rect 19260 36718 19288 37266
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 19248 35828 19300 35834
rect 19168 35788 19248 35816
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 19168 35222 19196 35788
rect 19248 35770 19300 35776
rect 19246 35728 19302 35737
rect 19246 35663 19248 35672
rect 19300 35663 19302 35672
rect 19248 35634 19300 35640
rect 19156 35216 19208 35222
rect 19156 35158 19208 35164
rect 19156 35012 19208 35018
rect 19156 34954 19208 34960
rect 19064 33856 19116 33862
rect 19064 33798 19116 33804
rect 18972 31476 19024 31482
rect 18972 31418 19024 31424
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 18788 31272 18840 31278
rect 18788 31214 18840 31220
rect 18880 31272 18932 31278
rect 18880 31214 18932 31220
rect 18800 30666 18828 31214
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18892 30546 18920 30738
rect 18800 30518 18920 30546
rect 18800 29714 18828 30518
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18788 29708 18840 29714
rect 18788 29650 18840 29656
rect 18800 27946 18828 29650
rect 18892 29238 18920 29990
rect 18880 29232 18932 29238
rect 18880 29174 18932 29180
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18892 28150 18920 28902
rect 18880 28144 18932 28150
rect 18880 28086 18932 28092
rect 18984 27962 19012 31282
rect 19076 28558 19104 33798
rect 19168 33658 19196 34954
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19260 32434 19288 32846
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19168 30598 19196 31826
rect 19352 31754 19380 36722
rect 19444 36650 19472 37130
rect 19432 36644 19484 36650
rect 19432 36586 19484 36592
rect 19536 36378 19564 38218
rect 19628 37806 19656 40530
rect 19812 40390 19840 41074
rect 19996 41002 20024 41414
rect 19984 40996 20036 41002
rect 19984 40938 20036 40944
rect 19800 40384 19852 40390
rect 19800 40326 19852 40332
rect 19984 40044 20036 40050
rect 19984 39986 20036 39992
rect 19708 39976 19760 39982
rect 19708 39918 19760 39924
rect 19616 37800 19668 37806
rect 19616 37742 19668 37748
rect 19524 36372 19576 36378
rect 19524 36314 19576 36320
rect 19720 35680 19748 39918
rect 19996 39846 20024 39986
rect 19984 39840 20036 39846
rect 19984 39782 20036 39788
rect 20088 39506 20116 43386
rect 20352 42900 20404 42906
rect 20352 42842 20404 42848
rect 20260 42016 20312 42022
rect 20260 41958 20312 41964
rect 20168 41268 20220 41274
rect 20168 41210 20220 41216
rect 20180 40662 20208 41210
rect 20168 40656 20220 40662
rect 20168 40598 20220 40604
rect 20076 39500 20128 39506
rect 20076 39442 20128 39448
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 19904 38282 19932 38898
rect 19984 38820 20036 38826
rect 19984 38762 20036 38768
rect 19892 38276 19944 38282
rect 19892 38218 19944 38224
rect 19798 37768 19854 37777
rect 19798 37703 19800 37712
rect 19852 37703 19854 37712
rect 19800 37674 19852 37680
rect 19800 37188 19852 37194
rect 19800 37130 19852 37136
rect 19536 35652 19748 35680
rect 19432 31952 19484 31958
rect 19430 31920 19432 31929
rect 19484 31920 19486 31929
rect 19430 31855 19486 31864
rect 19352 31726 19472 31754
rect 19340 31272 19392 31278
rect 19260 31232 19340 31260
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19156 30388 19208 30394
rect 19156 30330 19208 30336
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 18788 27940 18840 27946
rect 18788 27882 18840 27888
rect 18892 27934 19012 27962
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 18800 27577 18828 27610
rect 18786 27568 18842 27577
rect 18786 27503 18842 27512
rect 18786 27432 18842 27441
rect 18786 27367 18842 27376
rect 18602 26007 18658 26016
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18602 25800 18658 25809
rect 18602 25735 18658 25744
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18512 24948 18564 24954
rect 18512 24890 18564 24896
rect 18524 24721 18552 24890
rect 18510 24712 18566 24721
rect 18510 24647 18566 24656
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 22098 18552 24550
rect 18616 23746 18644 25735
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18708 23866 18736 25094
rect 18800 24750 18828 27367
rect 18892 24818 18920 27934
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18984 26450 19012 27814
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18788 24744 18840 24750
rect 18788 24686 18840 24692
rect 18800 24138 18828 24686
rect 18880 24676 18932 24682
rect 18880 24618 18932 24624
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18696 23860 18748 23866
rect 18748 23820 18828 23848
rect 18696 23802 18748 23808
rect 18616 23718 18736 23746
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18616 23186 18644 23598
rect 18604 23180 18656 23186
rect 18604 23122 18656 23128
rect 18616 22710 18644 23122
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 17776 22034 17828 22040
rect 18340 22066 18460 22094
rect 18512 22092 18564 22098
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17696 18970 17724 19246
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 12306 17172 13874
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17236 12986 17264 13126
rect 17328 12986 17356 15098
rect 17420 14006 17448 15506
rect 17408 14000 17460 14006
rect 17460 13948 17540 13954
rect 17408 13942 17540 13948
rect 17420 13926 17540 13942
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17512 12442 17540 13926
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16408 800 16436 4014
rect 16868 3058 16896 11494
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 800 16804 2790
rect 16960 2446 16988 9930
rect 17328 7478 17356 12106
rect 17420 12102 17448 12378
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17498 11928 17554 11937
rect 17498 11863 17500 11872
rect 17552 11863 17554 11872
rect 17500 11834 17552 11840
rect 17788 9654 17816 20198
rect 18340 19990 18368 22066
rect 18512 22034 18564 22040
rect 18708 21690 18736 23718
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18510 20632 18566 20641
rect 18510 20567 18566 20576
rect 18524 20466 18552 20567
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18800 20346 18828 23820
rect 18892 20942 18920 24618
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18524 20318 18828 20346
rect 18328 19984 18380 19990
rect 17866 19952 17922 19961
rect 18328 19926 18380 19932
rect 17866 19887 17922 19896
rect 17880 19854 17908 19887
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18340 14074 18368 18566
rect 18432 17270 18460 18634
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 18432 14278 18460 16118
rect 18524 14414 18552 20318
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18616 19417 18644 19722
rect 18602 19408 18658 19417
rect 18602 19343 18658 19352
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16250 18644 17070
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18616 15026 18644 16186
rect 18708 15502 18736 18362
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 15162 18736 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18432 13938 18460 14214
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18524 13818 18552 14214
rect 18432 13790 18552 13818
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18340 11898 18368 12718
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10130 18276 10406
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 18432 9586 18460 13790
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 11830 18552 13330
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17144 800 17172 2858
rect 17512 800 17540 4014
rect 17604 2582 17632 9386
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 5710 17724 9318
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4826 17816 5170
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18524 4622 18552 6598
rect 18616 4622 18644 12582
rect 18800 9926 18828 20198
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18892 18426 18920 19994
rect 18984 19854 19012 25706
rect 19076 25362 19104 27814
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19168 25242 19196 30330
rect 19076 25214 19196 25242
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18984 18902 19012 19654
rect 19076 18970 19104 25214
rect 19260 25106 19288 31232
rect 19340 31214 19392 31220
rect 19444 30734 19472 31726
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19340 30388 19392 30394
rect 19340 30330 19392 30336
rect 19352 30054 19380 30330
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19352 27674 19380 28018
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19352 26042 19380 26862
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19444 25294 19472 30534
rect 19536 29102 19564 35652
rect 19812 35578 19840 37130
rect 19904 36922 19932 38218
rect 19892 36916 19944 36922
rect 19892 36858 19944 36864
rect 19720 35550 19840 35578
rect 19720 35494 19748 35550
rect 19708 35488 19760 35494
rect 19708 35430 19760 35436
rect 19800 35488 19852 35494
rect 19800 35430 19852 35436
rect 19720 35154 19748 35430
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19708 35012 19760 35018
rect 19708 34954 19760 34960
rect 19616 34604 19668 34610
rect 19616 34546 19668 34552
rect 19628 33998 19656 34546
rect 19720 34202 19748 34954
rect 19812 34746 19840 35430
rect 19996 35018 20024 38762
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 20088 37670 20116 37878
rect 20076 37664 20128 37670
rect 20076 37606 20128 37612
rect 20180 37244 20208 40598
rect 20272 38418 20300 41958
rect 20364 39982 20392 42842
rect 20444 42560 20496 42566
rect 20444 42502 20496 42508
rect 20456 41274 20484 42502
rect 20548 42362 20576 47942
rect 20640 47025 20668 53450
rect 20732 53174 20760 54130
rect 20904 53984 20956 53990
rect 20904 53926 20956 53932
rect 20720 53168 20772 53174
rect 20720 53110 20772 53116
rect 20812 49972 20864 49978
rect 20812 49914 20864 49920
rect 20626 47016 20682 47025
rect 20626 46951 20682 46960
rect 20536 42356 20588 42362
rect 20536 42298 20588 42304
rect 20444 41268 20496 41274
rect 20444 41210 20496 41216
rect 20444 40384 20496 40390
rect 20444 40326 20496 40332
rect 20456 40118 20484 40326
rect 20444 40112 20496 40118
rect 20444 40054 20496 40060
rect 20352 39976 20404 39982
rect 20352 39918 20404 39924
rect 20352 39296 20404 39302
rect 20352 39238 20404 39244
rect 20444 39296 20496 39302
rect 20444 39238 20496 39244
rect 20260 38412 20312 38418
rect 20260 38354 20312 38360
rect 20180 37216 20300 37244
rect 20076 37120 20128 37126
rect 20076 37062 20128 37068
rect 20088 36582 20116 37062
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19800 34740 19852 34746
rect 19800 34682 19852 34688
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19892 34468 19944 34474
rect 19892 34410 19944 34416
rect 19708 34196 19760 34202
rect 19708 34138 19760 34144
rect 19800 34128 19852 34134
rect 19800 34070 19852 34076
rect 19616 33992 19668 33998
rect 19668 33952 19748 33980
rect 19616 33934 19668 33940
rect 19720 30734 19748 33952
rect 19812 31754 19840 34070
rect 19800 31748 19852 31754
rect 19800 31690 19852 31696
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 19904 30190 19932 34410
rect 19996 33930 20024 34614
rect 20088 33998 20116 36518
rect 20272 35630 20300 37216
rect 20260 35624 20312 35630
rect 20260 35566 20312 35572
rect 20260 35148 20312 35154
rect 20260 35090 20312 35096
rect 20168 34196 20220 34202
rect 20168 34138 20220 34144
rect 20076 33992 20128 33998
rect 20076 33934 20128 33940
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 20180 33862 20208 34138
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 19996 31890 20024 33594
rect 20180 33590 20208 33798
rect 20168 33584 20220 33590
rect 20168 33526 20220 33532
rect 20272 33436 20300 35090
rect 20180 33408 20300 33436
rect 20076 33040 20128 33046
rect 20076 32982 20128 32988
rect 20088 32774 20116 32982
rect 20076 32768 20128 32774
rect 20076 32710 20128 32716
rect 20076 32224 20128 32230
rect 20076 32166 20128 32172
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 20088 31686 20116 32166
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 20074 31512 20130 31521
rect 20074 31447 20076 31456
rect 20128 31447 20130 31456
rect 20076 31418 20128 31424
rect 20180 31362 20208 33408
rect 20364 33318 20392 39238
rect 20456 38894 20484 39238
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20456 38729 20484 38830
rect 20442 38720 20498 38729
rect 20442 38655 20498 38664
rect 20444 38208 20496 38214
rect 20444 38150 20496 38156
rect 20352 33312 20404 33318
rect 20352 33254 20404 33260
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20088 31334 20208 31362
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19892 30184 19944 30190
rect 19892 30126 19944 30132
rect 19524 29096 19576 29102
rect 19524 29038 19576 29044
rect 19536 28994 19564 29038
rect 19536 28966 19748 28994
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19720 26738 19748 28966
rect 19800 28484 19852 28490
rect 19904 28472 19932 30126
rect 19852 28444 19932 28472
rect 19800 28426 19852 28432
rect 19812 26926 19840 28426
rect 19996 28014 20024 30738
rect 20088 29238 20116 31334
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 20180 29578 20208 30194
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 20166 28248 20222 28257
rect 20166 28183 20168 28192
rect 20220 28183 20222 28192
rect 20168 28154 20220 28160
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19536 26042 19564 26726
rect 19720 26710 19840 26738
rect 19708 26512 19760 26518
rect 19708 26454 19760 26460
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19168 25078 19288 25106
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19168 20058 19196 25078
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19352 23050 19380 23190
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18892 15162 18920 17750
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18984 14278 19012 18838
rect 19076 18766 19104 18906
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19168 17134 19196 19858
rect 19260 19446 19288 22374
rect 19352 22098 19380 22578
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19444 21978 19472 25094
rect 19522 24984 19578 24993
rect 19522 24919 19578 24928
rect 19352 21950 19472 21978
rect 19352 20602 19380 21950
rect 19536 21894 19564 24919
rect 19720 22710 19748 26454
rect 19812 23746 19840 26710
rect 19890 24984 19946 24993
rect 19890 24919 19892 24928
rect 19944 24919 19946 24928
rect 19892 24890 19944 24896
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19904 23866 19932 24074
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19812 23718 19932 23746
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19812 22574 19840 23598
rect 19904 22930 19932 23718
rect 19996 23050 20024 27950
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20088 23322 20116 25298
rect 20180 24052 20208 26386
rect 20272 26382 20300 31894
rect 20456 31754 20484 38150
rect 20548 36922 20576 42298
rect 20720 42288 20772 42294
rect 20720 42230 20772 42236
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20640 40186 20668 42162
rect 20628 40180 20680 40186
rect 20628 40122 20680 40128
rect 20628 39840 20680 39846
rect 20628 39782 20680 39788
rect 20640 39302 20668 39782
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20628 39092 20680 39098
rect 20628 39034 20680 39040
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 20536 36032 20588 36038
rect 20536 35974 20588 35980
rect 20364 31726 20484 31754
rect 20364 30258 20392 31726
rect 20442 30968 20498 30977
rect 20548 30938 20576 35974
rect 20640 33998 20668 39034
rect 20732 37262 20760 42230
rect 20824 41274 20852 49914
rect 20916 45354 20944 53926
rect 21008 53582 21036 56200
rect 21376 54194 21404 56200
rect 21364 54188 21416 54194
rect 21364 54130 21416 54136
rect 21640 53984 21692 53990
rect 21640 53926 21692 53932
rect 21548 53712 21600 53718
rect 21548 53654 21600 53660
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 21008 53242 21036 53518
rect 21364 53440 21416 53446
rect 21364 53382 21416 53388
rect 20996 53236 21048 53242
rect 20996 53178 21048 53184
rect 21088 46368 21140 46374
rect 21088 46310 21140 46316
rect 20996 45824 21048 45830
rect 20996 45766 21048 45772
rect 20904 45348 20956 45354
rect 20904 45290 20956 45296
rect 20904 43444 20956 43450
rect 20904 43386 20956 43392
rect 20916 42702 20944 43386
rect 20904 42696 20956 42702
rect 20904 42638 20956 42644
rect 20916 42362 20944 42638
rect 20904 42356 20956 42362
rect 20904 42298 20956 42304
rect 20916 41682 20944 42298
rect 21008 42226 21036 45766
rect 21100 45422 21128 46310
rect 21376 46034 21404 53382
rect 21456 47252 21508 47258
rect 21456 47194 21508 47200
rect 21468 47025 21496 47194
rect 21454 47016 21510 47025
rect 21454 46951 21456 46960
rect 21508 46951 21510 46960
rect 21456 46922 21508 46928
rect 21364 46028 21416 46034
rect 21364 45970 21416 45976
rect 21456 46028 21508 46034
rect 21456 45970 21508 45976
rect 21272 45824 21324 45830
rect 21272 45766 21324 45772
rect 21088 45416 21140 45422
rect 21088 45358 21140 45364
rect 21100 44878 21128 45358
rect 21284 45354 21312 45766
rect 21468 45558 21496 45970
rect 21456 45552 21508 45558
rect 21456 45494 21508 45500
rect 21272 45348 21324 45354
rect 21272 45290 21324 45296
rect 21088 44872 21140 44878
rect 21088 44814 21140 44820
rect 21100 44470 21128 44814
rect 21272 44736 21324 44742
rect 21272 44678 21324 44684
rect 21088 44464 21140 44470
rect 21088 44406 21140 44412
rect 21100 43450 21128 44406
rect 21180 44328 21232 44334
rect 21180 44270 21232 44276
rect 21088 43444 21140 43450
rect 21088 43386 21140 43392
rect 21088 42628 21140 42634
rect 21088 42570 21140 42576
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 20904 41676 20956 41682
rect 20904 41618 20956 41624
rect 20996 41540 21048 41546
rect 20996 41482 21048 41488
rect 21008 41414 21036 41482
rect 20916 41386 21036 41414
rect 20812 41268 20864 41274
rect 20812 41210 20864 41216
rect 20812 40928 20864 40934
rect 20812 40870 20864 40876
rect 20824 39030 20852 40870
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20824 37194 20852 38422
rect 20916 38010 20944 41386
rect 20996 41268 21048 41274
rect 20996 41210 21048 41216
rect 21008 41070 21036 41210
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 21008 39098 21036 41006
rect 21100 40730 21128 42570
rect 21192 41750 21220 44270
rect 21284 43246 21312 44678
rect 21272 43240 21324 43246
rect 21272 43182 21324 43188
rect 21468 42906 21496 45494
rect 21560 43994 21588 53654
rect 21548 43988 21600 43994
rect 21548 43930 21600 43936
rect 21560 43722 21588 43930
rect 21548 43716 21600 43722
rect 21548 43658 21600 43664
rect 21456 42900 21508 42906
rect 21456 42842 21508 42848
rect 21272 42560 21324 42566
rect 21272 42502 21324 42508
rect 21284 42158 21312 42502
rect 21272 42152 21324 42158
rect 21272 42094 21324 42100
rect 21180 41744 21232 41750
rect 21180 41686 21232 41692
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 21088 39296 21140 39302
rect 21088 39238 21140 39244
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21100 38865 21128 39238
rect 21086 38856 21142 38865
rect 21086 38791 21142 38800
rect 21192 38418 21220 41686
rect 21560 41414 21588 43658
rect 21652 43450 21680 53926
rect 21744 53582 21772 56200
rect 22112 53582 22140 56200
rect 22480 54194 22508 56200
rect 22468 54188 22520 54194
rect 22468 54130 22520 54136
rect 22480 54074 22508 54130
rect 22480 54046 22600 54074
rect 22192 53984 22244 53990
rect 22284 53984 22336 53990
rect 22192 53926 22244 53932
rect 22282 53952 22284 53961
rect 22336 53952 22338 53961
rect 21732 53576 21784 53582
rect 21732 53518 21784 53524
rect 22100 53576 22152 53582
rect 22100 53518 22152 53524
rect 21744 53242 21772 53518
rect 22112 53242 22140 53518
rect 21732 53236 21784 53242
rect 21732 53178 21784 53184
rect 22100 53236 22152 53242
rect 22100 53178 22152 53184
rect 22204 52986 22232 53926
rect 22282 53887 22338 53896
rect 22376 53712 22428 53718
rect 22376 53654 22428 53660
rect 22112 52958 22232 52986
rect 22008 46912 22060 46918
rect 22008 46854 22060 46860
rect 21916 46708 21968 46714
rect 21916 46650 21968 46656
rect 21928 46374 21956 46650
rect 21916 46368 21968 46374
rect 21914 46336 21916 46345
rect 21968 46336 21970 46345
rect 21914 46271 21970 46280
rect 21916 43648 21968 43654
rect 21916 43590 21968 43596
rect 21640 43444 21692 43450
rect 21640 43386 21692 43392
rect 21652 43353 21680 43386
rect 21638 43344 21694 43353
rect 21638 43279 21694 43288
rect 21640 42832 21692 42838
rect 21640 42774 21692 42780
rect 21652 41478 21680 42774
rect 21640 41472 21692 41478
rect 21640 41414 21692 41420
rect 21376 41386 21588 41414
rect 21272 41200 21324 41206
rect 21272 41142 21324 41148
rect 21284 41070 21312 41142
rect 21272 41064 21324 41070
rect 21272 41006 21324 41012
rect 21272 40384 21324 40390
rect 21272 40326 21324 40332
rect 21284 39438 21312 40326
rect 21272 39432 21324 39438
rect 21272 39374 21324 39380
rect 21272 38752 21324 38758
rect 21272 38694 21324 38700
rect 21180 38412 21232 38418
rect 21180 38354 21232 38360
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 20904 38004 20956 38010
rect 20904 37946 20956 37952
rect 21100 37874 21128 38150
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20996 37188 21048 37194
rect 20996 37130 21048 37136
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20732 35154 20760 37062
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20720 35148 20772 35154
rect 20720 35090 20772 35096
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20640 33522 20668 33798
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20640 33114 20668 33458
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 20628 32360 20680 32366
rect 20626 32328 20628 32337
rect 20680 32328 20682 32337
rect 20626 32263 20682 32272
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 20442 30903 20444 30912
rect 20496 30903 20498 30912
rect 20536 30932 20588 30938
rect 20444 30874 20496 30880
rect 20536 30874 20588 30880
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20364 26042 20392 29446
rect 20456 29034 20484 30738
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20456 24682 20484 28970
rect 20548 27538 20576 30874
rect 20640 27538 20668 31214
rect 20732 29646 20760 34342
rect 20824 31822 20852 35974
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 20916 35154 20944 35430
rect 20904 35148 20956 35154
rect 20904 35090 20956 35096
rect 20916 34202 20944 35090
rect 21008 34746 21036 37130
rect 21100 37126 21128 37810
rect 21088 37120 21140 37126
rect 21088 37062 21140 37068
rect 21284 36242 21312 38694
rect 21272 36236 21324 36242
rect 21272 36178 21324 36184
rect 21376 36122 21404 41386
rect 21456 41268 21508 41274
rect 21456 41210 21508 41216
rect 21468 40934 21496 41210
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21100 36094 21404 36122
rect 20996 34740 21048 34746
rect 20996 34682 21048 34688
rect 20904 34196 20956 34202
rect 20904 34138 20956 34144
rect 20996 33448 21048 33454
rect 20996 33390 21048 33396
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 20916 32774 20944 33050
rect 21008 32910 21036 33390
rect 20996 32904 21048 32910
rect 20996 32846 21048 32852
rect 20904 32768 20956 32774
rect 20904 32710 20956 32716
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20916 32026 20944 32370
rect 20904 32020 20956 32026
rect 20904 31962 20956 31968
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20916 30394 20944 31962
rect 20904 30388 20956 30394
rect 20904 30330 20956 30336
rect 20720 29640 20772 29646
rect 21008 29594 21036 32506
rect 20720 29582 20772 29588
rect 20824 29566 21036 29594
rect 20824 28150 20852 29566
rect 20904 29504 20956 29510
rect 20904 29446 20956 29452
rect 20916 29306 20944 29446
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 21100 29186 21128 36094
rect 21468 36038 21496 40870
rect 21732 40452 21784 40458
rect 21732 40394 21784 40400
rect 21744 40050 21772 40394
rect 21732 40044 21784 40050
rect 21732 39986 21784 39992
rect 21744 39506 21772 39986
rect 21732 39500 21784 39506
rect 21732 39442 21784 39448
rect 21824 39296 21876 39302
rect 21824 39238 21876 39244
rect 21836 38010 21864 39238
rect 21928 38418 21956 43590
rect 22020 42770 22048 46854
rect 22112 46714 22140 52958
rect 22192 52896 22244 52902
rect 22192 52838 22244 52844
rect 22100 46708 22152 46714
rect 22100 46650 22152 46656
rect 22204 43858 22232 52838
rect 22284 45280 22336 45286
rect 22284 45222 22336 45228
rect 22296 44878 22324 45222
rect 22284 44872 22336 44878
rect 22284 44814 22336 44820
rect 22296 44334 22324 44814
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22192 43852 22244 43858
rect 22192 43794 22244 43800
rect 22388 43450 22416 53654
rect 22468 53440 22520 53446
rect 22468 53382 22520 53388
rect 22480 47122 22508 53382
rect 22572 53242 22600 54046
rect 22848 53582 22876 56200
rect 23216 55214 23244 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 23216 55186 23336 55214
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23308 53242 23336 55186
rect 23400 53582 23428 56063
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 22560 53236 22612 53242
rect 22560 53178 22612 53184
rect 23296 53236 23348 53242
rect 23296 53178 23348 53184
rect 23584 53106 23612 56200
rect 24490 55448 24546 55457
rect 24490 55383 24546 55392
rect 24504 54330 24532 55383
rect 24766 54632 24822 54641
rect 24766 54567 24822 54576
rect 24492 54324 24544 54330
rect 24492 54266 24544 54272
rect 23940 53984 23992 53990
rect 23940 53926 23992 53932
rect 23572 53100 23624 53106
rect 23572 53042 23624 53048
rect 23388 52896 23440 52902
rect 23388 52838 23440 52844
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22744 47592 22796 47598
rect 22744 47534 22796 47540
rect 22468 47116 22520 47122
rect 22468 47058 22520 47064
rect 22468 46504 22520 46510
rect 22468 46446 22520 46452
rect 22376 43444 22428 43450
rect 22376 43386 22428 43392
rect 22192 43376 22244 43382
rect 22192 43318 22244 43324
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22100 42560 22152 42566
rect 22100 42502 22152 42508
rect 22008 41472 22060 41478
rect 22008 41414 22060 41420
rect 22020 41274 22048 41414
rect 22008 41268 22060 41274
rect 22008 41210 22060 41216
rect 22006 40760 22062 40769
rect 22006 40695 22062 40704
rect 22020 40458 22048 40695
rect 22112 40594 22140 42502
rect 22204 41721 22232 43318
rect 22480 42514 22508 46446
rect 22652 46368 22704 46374
rect 22652 46310 22704 46316
rect 22560 44804 22612 44810
rect 22560 44746 22612 44752
rect 22572 44538 22600 44746
rect 22560 44532 22612 44538
rect 22560 44474 22612 44480
rect 22572 42770 22600 44474
rect 22560 42764 22612 42770
rect 22560 42706 22612 42712
rect 22296 42486 22508 42514
rect 22190 41712 22246 41721
rect 22190 41647 22246 41656
rect 22192 41540 22244 41546
rect 22192 41482 22244 41488
rect 22100 40588 22152 40594
rect 22100 40530 22152 40536
rect 22008 40452 22060 40458
rect 22008 40394 22060 40400
rect 22204 39642 22232 41482
rect 22296 41206 22324 42486
rect 22376 42356 22428 42362
rect 22376 42298 22428 42304
rect 22284 41200 22336 41206
rect 22284 41142 22336 41148
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22008 39432 22060 39438
rect 22008 39374 22060 39380
rect 21916 38412 21968 38418
rect 21916 38354 21968 38360
rect 21824 38004 21876 38010
rect 21824 37946 21876 37952
rect 21836 37466 21864 37946
rect 22020 37738 22048 39374
rect 22296 39302 22324 41142
rect 22284 39296 22336 39302
rect 22284 39238 22336 39244
rect 22388 39030 22416 42298
rect 22572 41834 22600 42706
rect 22480 41806 22600 41834
rect 22480 41682 22508 41806
rect 22560 41744 22612 41750
rect 22560 41686 22612 41692
rect 22468 41676 22520 41682
rect 22468 41618 22520 41624
rect 22466 41576 22522 41585
rect 22466 41511 22522 41520
rect 22480 41070 22508 41511
rect 22468 41064 22520 41070
rect 22468 41006 22520 41012
rect 22480 40610 22508 41006
rect 22572 40730 22600 41686
rect 22664 41682 22692 46310
rect 22756 43382 22784 47534
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22836 47116 22888 47122
rect 22836 47058 22888 47064
rect 22848 44282 22876 47058
rect 23400 46714 23428 52838
rect 23388 46708 23440 46714
rect 23388 46650 23440 46656
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 23664 45960 23716 45966
rect 23664 45902 23716 45908
rect 23572 45484 23624 45490
rect 23572 45426 23624 45432
rect 23388 45348 23440 45354
rect 23388 45290 23440 45296
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23020 44940 23072 44946
rect 23020 44882 23072 44888
rect 23032 44810 23060 44882
rect 23020 44804 23072 44810
rect 23020 44746 23072 44752
rect 23032 44470 23060 44746
rect 23400 44742 23428 45290
rect 23584 44946 23612 45426
rect 23572 44940 23624 44946
rect 23572 44882 23624 44888
rect 23388 44736 23440 44742
rect 23388 44678 23440 44684
rect 23020 44464 23072 44470
rect 23020 44406 23072 44412
rect 22928 44328 22980 44334
rect 22848 44276 22928 44282
rect 22848 44270 22980 44276
rect 22848 44254 22968 44270
rect 22744 43376 22796 43382
rect 22744 43318 22796 43324
rect 22744 43240 22796 43246
rect 22744 43182 22796 43188
rect 22652 41676 22704 41682
rect 22652 41618 22704 41624
rect 22560 40724 22612 40730
rect 22560 40666 22612 40672
rect 22480 40582 22600 40610
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22480 40186 22508 40462
rect 22468 40180 22520 40186
rect 22468 40122 22520 40128
rect 22376 39024 22428 39030
rect 22376 38966 22428 38972
rect 22100 38888 22152 38894
rect 22100 38830 22152 38836
rect 22112 37738 22140 38830
rect 22388 38554 22416 38966
rect 22572 38842 22600 40582
rect 22652 40384 22704 40390
rect 22652 40326 22704 40332
rect 22480 38814 22600 38842
rect 22192 38548 22244 38554
rect 22192 38490 22244 38496
rect 22376 38548 22428 38554
rect 22376 38490 22428 38496
rect 22008 37732 22060 37738
rect 22008 37674 22060 37680
rect 22100 37732 22152 37738
rect 22100 37674 22152 37680
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 22112 37262 22140 37674
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22112 36786 22140 37198
rect 22100 36780 22152 36786
rect 22100 36722 22152 36728
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 21640 36236 21692 36242
rect 21640 36178 21692 36184
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21548 35828 21600 35834
rect 21548 35770 21600 35776
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 21192 34746 21220 35226
rect 21180 34740 21232 34746
rect 21180 34682 21232 34688
rect 21456 33856 21508 33862
rect 21456 33798 21508 33804
rect 21468 33658 21496 33798
rect 21180 33652 21232 33658
rect 21180 33594 21232 33600
rect 21456 33652 21508 33658
rect 21456 33594 21508 33600
rect 21192 32910 21220 33594
rect 21560 32994 21588 35770
rect 21652 35154 21680 36178
rect 21640 35148 21692 35154
rect 21640 35090 21692 35096
rect 21652 34066 21680 35090
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21652 33386 21680 34002
rect 21640 33380 21692 33386
rect 21640 33322 21692 33328
rect 21376 32966 21588 32994
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21272 32768 21324 32774
rect 21272 32710 21324 32716
rect 21178 32328 21234 32337
rect 21178 32263 21234 32272
rect 21192 31754 21220 32263
rect 21284 31754 21312 32710
rect 21376 32366 21404 32966
rect 21560 32960 21588 32966
rect 21640 32972 21692 32978
rect 21560 32932 21640 32960
rect 21640 32914 21692 32920
rect 21456 32904 21508 32910
rect 21508 32864 21588 32892
rect 21456 32846 21508 32852
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21376 31890 21404 32166
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21560 31754 21588 32864
rect 21640 32768 21692 32774
rect 21638 32736 21640 32745
rect 21692 32736 21694 32745
rect 21638 32671 21694 32680
rect 21652 31958 21680 32671
rect 21744 32337 21772 36314
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 21822 32600 21878 32609
rect 21822 32535 21824 32544
rect 21876 32535 21878 32544
rect 21824 32506 21876 32512
rect 21730 32328 21786 32337
rect 21730 32263 21786 32272
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21640 31952 21692 31958
rect 21640 31894 21692 31900
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21180 31748 21232 31754
rect 21180 31690 21232 31696
rect 21272 31748 21324 31754
rect 21272 31690 21324 31696
rect 21376 31726 21588 31754
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21008 29158 21128 29186
rect 21008 29102 21036 29158
rect 20996 29096 21048 29102
rect 20996 29038 21048 29044
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20640 26858 20668 27474
rect 20628 26852 20680 26858
rect 20628 26794 20680 26800
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20640 24818 20668 26386
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20260 24064 20312 24070
rect 20180 24024 20260 24052
rect 20260 24006 20312 24012
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19904 22902 20024 22930
rect 19800 22568 19852 22574
rect 19852 22516 19932 22522
rect 19800 22510 19932 22516
rect 19812 22494 19932 22510
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 19812 21962 19840 22034
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19524 21888 19576 21894
rect 19524 21830 19576 21836
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19536 21350 19564 21422
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19812 21010 19840 21898
rect 19904 21894 19932 22494
rect 19996 22094 20024 22902
rect 20272 22234 20300 24006
rect 20548 23866 20576 24686
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20640 23798 20668 24618
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 19996 22066 20300 22094
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19444 20466 19472 20810
rect 20180 20777 20208 21082
rect 20166 20768 20222 20777
rect 20166 20703 20222 20712
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19536 19378 19564 19654
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19064 16992 19116 16998
rect 19260 16946 19288 19178
rect 19352 18426 19380 19246
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19352 17134 19380 18362
rect 19444 18358 19472 18634
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19444 17542 19472 18294
rect 19536 17882 19564 19314
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17270 19472 17478
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19116 16940 19288 16946
rect 19064 16934 19288 16940
rect 19076 16918 19288 16934
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18892 13530 18920 14010
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12850 18920 13126
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18984 12238 19012 13806
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18984 12102 19012 12174
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17880 800 17908 3538
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18708 3058 18736 9590
rect 19076 8566 19104 16918
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19352 16182 19380 16662
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 12238 19196 14758
rect 19260 12986 19288 15438
rect 19352 13190 19380 15574
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19432 13456 19484 13462
rect 19430 13424 19432 13433
rect 19484 13424 19486 13433
rect 19430 13359 19486 13368
rect 19536 13274 19564 14826
rect 19444 13246 19564 13274
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11898 19288 12038
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19444 10554 19472 13246
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19536 10674 19564 12786
rect 19628 12374 19656 15302
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10810 19656 10950
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19352 10526 19472 10554
rect 19064 8560 19116 8566
rect 19064 8502 19116 8508
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18800 4049 18828 4082
rect 18786 4040 18842 4049
rect 18786 3975 18842 3984
rect 18800 3738 18828 3975
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 19352 3534 19380 10526
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17972 2514 18000 2790
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18340 1170 18368 2314
rect 18248 1142 18368 1170
rect 18248 800 18276 1142
rect 18616 800 18644 2790
rect 18708 2650 18736 2994
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18984 800 19012 3402
rect 19444 2446 19472 9998
rect 19720 6914 19748 18566
rect 19812 15026 19840 20198
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19904 16250 19932 19314
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19904 14822 19932 15438
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19812 12170 19840 14758
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19812 7886 19840 12106
rect 19904 11150 19932 14758
rect 19996 14278 20024 19926
rect 20180 18222 20208 20703
rect 20272 20058 20300 22066
rect 20364 21434 20392 22714
rect 20456 22094 20484 23258
rect 20456 22066 20576 22094
rect 20364 21406 20484 21434
rect 20456 21350 20484 21406
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20272 19514 20300 19994
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20456 18766 20484 21286
rect 20548 21010 20576 22066
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20536 21004 20588 21010
rect 20536 20946 20588 20952
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17610 20208 18022
rect 20168 17604 20220 17610
rect 20168 17546 20220 17552
rect 20180 16658 20208 17546
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20456 16590 20484 17070
rect 20548 16590 20576 19382
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20640 16436 20668 21422
rect 20732 19854 20760 24346
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23526 20852 23598
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 21008 21486 21036 29038
rect 21192 28694 21220 29650
rect 21272 28756 21324 28762
rect 21272 28698 21324 28704
rect 21180 28688 21232 28694
rect 21180 28630 21232 28636
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 21100 25362 21128 27542
rect 21192 26926 21220 28630
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21192 26314 21220 26862
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20456 16408 20668 16436
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19996 13938 20024 14214
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20088 13258 20116 14350
rect 20456 13938 20484 16408
rect 20732 16250 20760 19110
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20824 15502 20852 21286
rect 20996 20324 21048 20330
rect 20996 20266 21048 20272
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 17746 20944 18634
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20916 17338 20944 17682
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20916 16658 20944 17274
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19996 11898 20024 12242
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19996 10538 20024 11834
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19536 6886 19748 6914
rect 19536 5234 19564 6886
rect 20364 5710 20392 13806
rect 20456 13530 20484 13874
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 10674 20576 12582
rect 20640 11082 20668 15302
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20824 11830 20852 14486
rect 20916 14414 20944 16594
rect 21008 16182 21036 20266
rect 21100 18358 21128 21558
rect 21192 19514 21220 25638
rect 21284 22094 21312 28698
rect 21376 27062 21404 31726
rect 21456 31680 21508 31686
rect 21456 31622 21508 31628
rect 21468 28914 21496 31622
rect 21652 31482 21680 31758
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21836 31346 21864 32166
rect 21928 31822 21956 36110
rect 22204 35816 22232 38490
rect 22480 38434 22508 38814
rect 22560 38752 22612 38758
rect 22560 38694 22612 38700
rect 22112 35788 22232 35816
rect 22296 38406 22508 38434
rect 22572 38418 22600 38694
rect 22560 38412 22612 38418
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21548 30116 21600 30122
rect 21548 30058 21600 30064
rect 21560 29238 21588 30058
rect 21732 30048 21784 30054
rect 21732 29990 21784 29996
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 21640 29028 21692 29034
rect 21640 28970 21692 28976
rect 21468 28886 21588 28914
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21468 28150 21496 28426
rect 21456 28144 21508 28150
rect 21456 28086 21508 28092
rect 21364 27056 21416 27062
rect 21364 26998 21416 27004
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21468 26450 21496 26862
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 21376 24138 21404 25978
rect 21560 25974 21588 28886
rect 21652 26450 21680 28970
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 25968 21600 25974
rect 21548 25910 21600 25916
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25294 21680 25774
rect 21640 25288 21692 25294
rect 21640 25230 21692 25236
rect 21744 24206 21772 29990
rect 21836 26246 21864 30534
rect 21928 29510 21956 31146
rect 22020 29646 22048 34342
rect 22112 32434 22140 35788
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22204 35086 22232 35634
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22204 33522 22232 35022
rect 22296 34610 22324 38406
rect 22560 38354 22612 38360
rect 22468 37392 22520 37398
rect 22468 37334 22520 37340
rect 22376 36712 22428 36718
rect 22480 36689 22508 37334
rect 22376 36654 22428 36660
rect 22466 36680 22522 36689
rect 22388 36038 22416 36654
rect 22466 36615 22522 36624
rect 22480 36281 22508 36615
rect 22466 36272 22522 36281
rect 22466 36207 22522 36216
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22388 34746 22416 35974
rect 22468 35624 22520 35630
rect 22468 35566 22520 35572
rect 22480 34746 22508 35566
rect 22572 35018 22600 38354
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22296 34202 22324 34546
rect 22374 34368 22430 34377
rect 22374 34303 22430 34312
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22100 32224 22152 32230
rect 22100 32166 22152 32172
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 22020 28082 22048 28562
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 22020 27554 22048 28018
rect 21928 27538 22048 27554
rect 21916 27532 22048 27538
rect 21968 27526 22048 27532
rect 21916 27474 21968 27480
rect 22020 26926 22048 27526
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 21824 26240 21876 26246
rect 21824 26182 21876 26188
rect 22112 25770 22140 32166
rect 22204 31278 22232 33458
rect 22192 31272 22244 31278
rect 22192 31214 22244 31220
rect 22204 30258 22232 31214
rect 22296 30734 22324 33798
rect 22388 32910 22416 34303
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22376 32904 22428 32910
rect 22376 32846 22428 32852
rect 22480 32842 22508 33798
rect 22572 33046 22600 34954
rect 22664 34610 22692 40326
rect 22756 38570 22784 43182
rect 22848 42786 22876 44254
rect 23296 44192 23348 44198
rect 23296 44134 23348 44140
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23308 43994 23336 44134
rect 23296 43988 23348 43994
rect 23296 43930 23348 43936
rect 23296 43852 23348 43858
rect 23296 43794 23348 43800
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22848 42758 22968 42786
rect 22836 42696 22888 42702
rect 22836 42638 22888 42644
rect 22848 42158 22876 42638
rect 22940 42242 22968 42758
rect 23112 42764 23164 42770
rect 23112 42706 23164 42712
rect 23124 42401 23152 42706
rect 23110 42392 23166 42401
rect 23308 42362 23336 43794
rect 23110 42327 23166 42336
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 22940 42214 23336 42242
rect 22836 42152 22888 42158
rect 22836 42094 22888 42100
rect 22848 41070 22876 42094
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22928 41812 22980 41818
rect 22928 41754 22980 41760
rect 22940 41721 22968 41754
rect 22926 41712 22982 41721
rect 22926 41647 22982 41656
rect 23204 41200 23256 41206
rect 23204 41142 23256 41148
rect 23216 41070 23244 41142
rect 22836 41064 22888 41070
rect 22836 41006 22888 41012
rect 23204 41064 23256 41070
rect 23204 41006 23256 41012
rect 22848 40118 22876 41006
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 23032 40526 23060 40666
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 22928 40384 22980 40390
rect 22928 40326 22980 40332
rect 22836 40112 22888 40118
rect 22836 40054 22888 40060
rect 22940 40050 22968 40326
rect 23308 40186 23336 42214
rect 23400 40594 23428 44678
rect 23584 43994 23612 44882
rect 23480 43988 23532 43994
rect 23480 43930 23532 43936
rect 23572 43988 23624 43994
rect 23572 43930 23624 43936
rect 23492 43246 23520 43930
rect 23572 43376 23624 43382
rect 23572 43318 23624 43324
rect 23480 43240 23532 43246
rect 23480 43182 23532 43188
rect 23492 42158 23520 43182
rect 23480 42152 23532 42158
rect 23480 42094 23532 42100
rect 23584 41970 23612 43318
rect 23492 41942 23612 41970
rect 23492 41682 23520 41942
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23492 41274 23520 41618
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23388 40588 23440 40594
rect 23388 40530 23440 40536
rect 23296 40180 23348 40186
rect 23296 40122 23348 40128
rect 22928 40044 22980 40050
rect 22928 39986 22980 39992
rect 23388 39976 23440 39982
rect 23388 39918 23440 39924
rect 22836 39908 22888 39914
rect 22836 39850 22888 39856
rect 22848 38894 22876 39850
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22836 38888 22888 38894
rect 22836 38830 22888 38836
rect 23400 38826 23428 39918
rect 23492 39506 23520 41210
rect 23480 39500 23532 39506
rect 23480 39442 23532 39448
rect 23388 38820 23440 38826
rect 23388 38762 23440 38768
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22756 38542 22876 38570
rect 22744 38480 22796 38486
rect 22744 38422 22796 38428
rect 22652 34604 22704 34610
rect 22652 34546 22704 34552
rect 22652 34468 22704 34474
rect 22652 34410 22704 34416
rect 22560 33040 22612 33046
rect 22560 32982 22612 32988
rect 22468 32836 22520 32842
rect 22468 32778 22520 32784
rect 22376 32768 22428 32774
rect 22560 32768 22612 32774
rect 22376 32710 22428 32716
rect 22558 32736 22560 32745
rect 22612 32736 22614 32745
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22284 27396 22336 27402
rect 22284 27338 22336 27344
rect 22204 26586 22232 27338
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22204 25906 22232 26522
rect 22296 26382 22324 27338
rect 22284 26376 22336 26382
rect 22284 26318 22336 26324
rect 22296 26042 22324 26318
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22100 25764 22152 25770
rect 22100 25706 22152 25712
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21376 23730 21404 24074
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21376 23594 21404 23666
rect 21364 23588 21416 23594
rect 21364 23530 21416 23536
rect 21376 23322 21404 23530
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21376 23050 21404 23258
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21376 22234 21404 22986
rect 22020 22642 22048 23666
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21364 22228 21416 22234
rect 21416 22188 21496 22216
rect 21364 22170 21416 22176
rect 21284 22066 21404 22094
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21284 21690 21312 21830
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 12986 20944 14350
rect 21100 14074 21128 18158
rect 21284 17882 21312 19246
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 15570 21220 16390
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 14482 21220 15506
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13938 21128 14010
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20628 11076 20680 11082
rect 20628 11018 20680 11024
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20640 10554 20668 11018
rect 20824 10606 20852 11018
rect 20548 10526 20668 10554
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20548 7886 20576 10526
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 8974 20668 10406
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19616 5160 19668 5166
rect 19616 5102 19668 5108
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19352 870 19472 898
rect 19352 800 19380 870
rect 13188 734 13400 762
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19444 762 19472 870
rect 19628 762 19656 5102
rect 19720 4010 19748 5238
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19720 800 19748 2858
rect 19904 2854 19932 4626
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 20088 800 20116 4014
rect 20456 800 20484 5714
rect 20640 5710 20668 7210
rect 20824 6798 20852 7686
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20640 2990 20668 4490
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20732 2922 20760 4626
rect 20824 3670 20852 6190
rect 20916 5914 20944 7346
rect 21100 6322 21128 7686
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20812 2916 20864 2922
rect 20812 2858 20864 2864
rect 20824 800 20852 2858
rect 21100 2802 21128 5578
rect 21192 3534 21220 14282
rect 21376 13870 21404 22066
rect 21468 21962 21496 22188
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21468 21146 21496 21898
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21468 20942 21496 21082
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21652 20806 21680 22510
rect 22020 22098 22048 22578
rect 22008 22092 22060 22098
rect 22008 22034 22060 22040
rect 22020 21622 22048 22034
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 20398 21680 20742
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 21468 13938 21496 19382
rect 21928 19310 21956 19450
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 21928 16640 21956 19246
rect 22020 18766 22048 19246
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22112 18290 22140 24006
rect 22296 22094 22324 25774
rect 22388 25226 22416 32710
rect 22558 32671 22614 32680
rect 22572 31226 22600 32671
rect 22664 31482 22692 34410
rect 22756 34066 22784 38422
rect 22848 37806 22876 38542
rect 23400 37942 23428 38762
rect 23570 38584 23626 38593
rect 23570 38519 23626 38528
rect 23584 38282 23612 38519
rect 23572 38276 23624 38282
rect 23572 38218 23624 38224
rect 23388 37936 23440 37942
rect 23202 37904 23258 37913
rect 23388 37878 23440 37884
rect 23202 37839 23204 37848
rect 23256 37839 23258 37848
rect 23204 37810 23256 37816
rect 22836 37800 22888 37806
rect 22836 37742 22888 37748
rect 22848 36922 22876 37742
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22836 36916 22888 36922
rect 22836 36858 22888 36864
rect 23296 36916 23348 36922
rect 23296 36858 23348 36864
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22848 35698 22876 36722
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22926 36272 22982 36281
rect 22926 36207 22982 36216
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22940 35578 22968 36207
rect 23308 35834 23336 36858
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 22848 35550 22968 35578
rect 22744 34060 22796 34066
rect 22744 34002 22796 34008
rect 22744 33312 22796 33318
rect 22744 33254 22796 33260
rect 22756 32434 22784 33254
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22652 31476 22704 31482
rect 22652 31418 22704 31424
rect 22480 31198 22600 31226
rect 22480 26042 22508 31198
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 22572 27282 22600 29650
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22664 27402 22692 28154
rect 22756 27538 22784 32166
rect 22848 30938 22876 35550
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23308 33454 23336 35770
rect 23400 35714 23428 37878
rect 23584 37670 23612 38218
rect 23572 37664 23624 37670
rect 23572 37606 23624 37612
rect 23676 37330 23704 45902
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 23664 37324 23716 37330
rect 23664 37266 23716 37272
rect 23768 36242 23796 38150
rect 23860 37942 23888 38354
rect 23848 37936 23900 37942
rect 23848 37878 23900 37884
rect 23860 36922 23888 37878
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23756 36236 23808 36242
rect 23756 36178 23808 36184
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35894 23704 35974
rect 23584 35866 23704 35894
rect 23400 35686 23520 35714
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23400 34950 23428 35566
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23400 34066 23428 34886
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23492 33946 23520 35686
rect 23584 34542 23612 35866
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23400 33918 23520 33946
rect 23296 33448 23348 33454
rect 23296 33390 23348 33396
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 23400 32450 23428 33918
rect 23676 33590 23704 34478
rect 23860 34474 23888 36858
rect 23952 35578 23980 53926
rect 24780 53582 24808 54567
rect 24952 54188 25004 54194
rect 24952 54130 25004 54136
rect 24964 53825 24992 54130
rect 25780 53984 25832 53990
rect 25780 53926 25832 53932
rect 24950 53816 25006 53825
rect 24950 53751 25006 53760
rect 25318 53816 25374 53825
rect 25318 53751 25374 53760
rect 24768 53576 24820 53582
rect 24768 53518 24820 53524
rect 24032 53508 24084 53514
rect 24032 53450 24084 53456
rect 24044 38350 24072 53450
rect 24780 52698 24808 53518
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 25056 53009 25084 53042
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24952 52896 25004 52902
rect 24952 52838 25004 52844
rect 24768 52692 24820 52698
rect 24768 52634 24820 52640
rect 24768 52488 24820 52494
rect 24768 52430 24820 52436
rect 24780 52193 24808 52430
rect 24766 52184 24822 52193
rect 24766 52119 24822 52128
rect 24768 46980 24820 46986
rect 24768 46922 24820 46928
rect 24492 46504 24544 46510
rect 24492 46446 24544 46452
rect 24584 46504 24636 46510
rect 24780 46481 24808 46922
rect 24584 46446 24636 46452
rect 24766 46472 24822 46481
rect 24504 46170 24532 46446
rect 24492 46164 24544 46170
rect 24492 46106 24544 46112
rect 24124 45484 24176 45490
rect 24124 45426 24176 45432
rect 24032 38344 24084 38350
rect 24032 38286 24084 38292
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 24044 37330 24072 37606
rect 24136 37398 24164 45426
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24504 44742 24532 45358
rect 24492 44736 24544 44742
rect 24492 44678 24544 44684
rect 24216 43988 24268 43994
rect 24216 43930 24268 43936
rect 24228 43450 24256 43930
rect 24216 43444 24268 43450
rect 24216 43386 24268 43392
rect 24228 42906 24256 43386
rect 24216 42900 24268 42906
rect 24216 42842 24268 42848
rect 24228 42294 24256 42842
rect 24216 42288 24268 42294
rect 24216 42230 24268 42236
rect 24228 41818 24256 42230
rect 24216 41812 24268 41818
rect 24216 41754 24268 41760
rect 24228 41206 24256 41754
rect 24216 41200 24268 41206
rect 24216 41142 24268 41148
rect 24228 40730 24256 41142
rect 24216 40724 24268 40730
rect 24216 40666 24268 40672
rect 24228 40118 24256 40666
rect 24216 40112 24268 40118
rect 24216 40054 24268 40060
rect 24228 39030 24256 40054
rect 24492 39976 24544 39982
rect 24492 39918 24544 39924
rect 24308 39296 24360 39302
rect 24308 39238 24360 39244
rect 24216 39024 24268 39030
rect 24216 38966 24268 38972
rect 24216 38888 24268 38894
rect 24216 38830 24268 38836
rect 24228 38282 24256 38830
rect 24216 38276 24268 38282
rect 24216 38218 24268 38224
rect 24124 37392 24176 37398
rect 24124 37334 24176 37340
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 23952 35550 24072 35578
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23664 33584 23716 33590
rect 23664 33526 23716 33532
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23308 32422 23428 32450
rect 23308 32230 23336 32422
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 32026 23336 32166
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22848 30598 22876 30874
rect 22836 30592 22888 30598
rect 22836 30534 22888 30540
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23400 29714 23428 31894
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23492 31226 23520 31826
rect 23492 31198 23612 31226
rect 23584 31142 23612 31198
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30326 23612 31078
rect 23572 30320 23624 30326
rect 23572 30262 23624 30268
rect 23388 29708 23440 29714
rect 23388 29650 23440 29656
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 22848 28626 22876 29446
rect 23308 29034 23336 29446
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23296 29028 23348 29034
rect 23296 28970 23348 28976
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 23400 28200 23428 28970
rect 23308 28172 23428 28200
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22744 27532 22796 27538
rect 22744 27474 22796 27480
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22756 27390 23152 27418
rect 22572 27254 22692 27282
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 22572 26858 22600 27066
rect 22560 26852 22612 26858
rect 22560 26794 22612 26800
rect 22664 26586 22692 27254
rect 22756 27130 22784 27390
rect 23124 27334 23152 27390
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 23032 27062 23060 27270
rect 23020 27056 23072 27062
rect 23020 26998 23072 27004
rect 23204 26920 23256 26926
rect 22756 26868 23204 26874
rect 22756 26862 23256 26868
rect 22756 26846 23244 26862
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22480 25498 22508 25978
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22376 25220 22428 25226
rect 22376 25162 22428 25168
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22204 22066 22324 22094
rect 22204 19292 22232 22066
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21486 22324 21898
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22284 19304 22336 19310
rect 22204 19264 22284 19292
rect 22284 19246 22336 19252
rect 22296 18970 22324 19246
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22008 16652 22060 16658
rect 21928 16612 22008 16640
rect 22008 16594 22060 16600
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21270 13424 21326 13433
rect 21270 13359 21326 13368
rect 21284 10062 21312 13359
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21468 12986 21496 13262
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21284 4622 21312 8298
rect 21376 6322 21404 11630
rect 21560 9654 21588 15302
rect 21548 9648 21600 9654
rect 21548 9590 21600 9596
rect 21652 8566 21680 16118
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21836 15434 21864 15846
rect 21824 15428 21876 15434
rect 21824 15370 21876 15376
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21100 2774 21220 2802
rect 21192 800 21220 2774
rect 21560 800 21588 5714
rect 21652 2417 21680 7278
rect 21744 6914 21772 13942
rect 21836 12782 21864 14214
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21836 12306 21864 12718
rect 21928 12306 21956 15846
rect 22112 12850 22140 16458
rect 22296 16046 22324 18906
rect 22388 16402 22416 24006
rect 22572 21690 22600 26454
rect 22664 25362 22692 26522
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22756 23118 22784 26846
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22836 25764 22888 25770
rect 22836 25706 22888 25712
rect 22848 25294 22876 25706
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23204 25356 23256 25362
rect 23204 25298 23256 25304
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 23216 24886 23244 25298
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22848 24274 22876 24754
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22848 23730 22876 24210
rect 23308 24206 23336 28172
rect 23492 28132 23520 29106
rect 23584 29102 23612 30262
rect 23768 30190 23796 33390
rect 23952 31482 23980 35430
rect 24044 33046 24072 35550
rect 24320 33998 24348 39238
rect 24504 37806 24532 39918
rect 24492 37800 24544 37806
rect 24492 37742 24544 37748
rect 24400 37324 24452 37330
rect 24400 37266 24452 37272
rect 24412 36786 24440 37266
rect 24400 36780 24452 36786
rect 24400 36722 24452 36728
rect 24400 36304 24452 36310
rect 24400 36246 24452 36252
rect 24216 33992 24268 33998
rect 24216 33934 24268 33940
rect 24308 33992 24360 33998
rect 24308 33934 24360 33940
rect 24032 33040 24084 33046
rect 24032 32982 24084 32988
rect 24228 32026 24256 33934
rect 24308 33856 24360 33862
rect 24308 33798 24360 33804
rect 24320 33590 24348 33798
rect 24308 33584 24360 33590
rect 24308 33526 24360 33532
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 24320 31822 24348 33526
rect 24308 31816 24360 31822
rect 24308 31758 24360 31764
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 24320 31414 24348 31758
rect 24308 31408 24360 31414
rect 24308 31350 24360 31356
rect 24320 30394 24348 31350
rect 24412 31346 24440 36246
rect 24504 36242 24532 37742
rect 24492 36236 24544 36242
rect 24492 36178 24544 36184
rect 24596 36174 24624 46446
rect 24766 46407 24822 46416
rect 24860 45824 24912 45830
rect 24860 45766 24912 45772
rect 24872 45665 24900 45766
rect 24858 45656 24914 45665
rect 24858 45591 24914 45600
rect 24964 45554 24992 52838
rect 25332 52154 25360 53751
rect 25688 53440 25740 53446
rect 25688 53382 25740 53388
rect 25320 52148 25372 52154
rect 25320 52090 25372 52096
rect 25504 51808 25556 51814
rect 25504 51750 25556 51756
rect 25516 51406 25544 51750
rect 25504 51400 25556 51406
rect 25502 51368 25504 51377
rect 25556 51368 25558 51377
rect 25502 51303 25558 51312
rect 25228 51264 25280 51270
rect 25228 51206 25280 51212
rect 25240 51105 25268 51206
rect 25226 51096 25282 51105
rect 25226 51031 25282 51040
rect 25044 50924 25096 50930
rect 25044 50866 25096 50872
rect 25056 50561 25084 50866
rect 25042 50552 25098 50561
rect 25042 50487 25098 50496
rect 25320 50176 25372 50182
rect 25320 50118 25372 50124
rect 25332 49842 25360 50118
rect 25320 49836 25372 49842
rect 25320 49778 25372 49784
rect 25332 49745 25360 49778
rect 25318 49736 25374 49745
rect 25318 49671 25374 49680
rect 25320 49224 25372 49230
rect 25320 49166 25372 49172
rect 25332 48929 25360 49166
rect 25318 48920 25374 48929
rect 25318 48855 25374 48864
rect 25504 48544 25556 48550
rect 25504 48486 25556 48492
rect 25320 48136 25372 48142
rect 25318 48104 25320 48113
rect 25372 48104 25374 48113
rect 25318 48039 25374 48048
rect 25516 47666 25544 48486
rect 25504 47660 25556 47666
rect 25504 47602 25556 47608
rect 25516 47297 25544 47602
rect 25502 47288 25558 47297
rect 25502 47223 25558 47232
rect 25596 47184 25648 47190
rect 25596 47126 25648 47132
rect 25504 46164 25556 46170
rect 25504 46106 25556 46112
rect 24872 45526 24992 45554
rect 24768 44328 24820 44334
rect 24766 44296 24768 44305
rect 24820 44296 24822 44305
rect 24766 44231 24822 44240
rect 24872 42770 24900 45526
rect 25516 44849 25544 46106
rect 25502 44840 25558 44849
rect 25502 44775 25558 44784
rect 25504 44736 25556 44742
rect 25504 44678 25556 44684
rect 25320 44396 25372 44402
rect 25320 44338 25372 44344
rect 25332 43654 25360 44338
rect 25516 44033 25544 44678
rect 25502 44024 25558 44033
rect 25502 43959 25558 43968
rect 25320 43648 25372 43654
rect 25320 43590 25372 43596
rect 25332 43217 25360 43590
rect 25318 43208 25374 43217
rect 25318 43143 25374 43152
rect 24952 43104 25004 43110
rect 24952 43046 25004 43052
rect 25136 43104 25188 43110
rect 25136 43046 25188 43052
rect 24860 42764 24912 42770
rect 24860 42706 24912 42712
rect 24860 42560 24912 42566
rect 24860 42502 24912 42508
rect 24872 42401 24900 42502
rect 24858 42392 24914 42401
rect 24858 42327 24914 42336
rect 24860 41472 24912 41478
rect 24860 41414 24912 41420
rect 24872 41070 24900 41414
rect 24860 41064 24912 41070
rect 24860 41006 24912 41012
rect 24768 40452 24820 40458
rect 24768 40394 24820 40400
rect 24780 39114 24808 40394
rect 24858 39128 24914 39137
rect 24780 39086 24858 39114
rect 24858 39063 24914 39072
rect 24872 38962 24900 39063
rect 24860 38956 24912 38962
rect 24860 38898 24912 38904
rect 24964 38350 24992 43046
rect 25148 42158 25176 43046
rect 25136 42152 25188 42158
rect 25136 42094 25188 42100
rect 25044 41744 25096 41750
rect 25044 41686 25096 41692
rect 25056 39506 25084 41686
rect 25148 39506 25176 42094
rect 25412 41744 25464 41750
rect 25412 41686 25464 41692
rect 25320 41608 25372 41614
rect 25318 41576 25320 41585
rect 25372 41576 25374 41585
rect 25318 41511 25374 41520
rect 25320 41472 25372 41478
rect 25320 41414 25372 41420
rect 25332 41138 25360 41414
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25320 40520 25372 40526
rect 25320 40462 25372 40468
rect 25228 40452 25280 40458
rect 25228 40394 25280 40400
rect 25240 39794 25268 40394
rect 25332 39953 25360 40462
rect 25318 39944 25374 39953
rect 25318 39879 25374 39888
rect 25240 39766 25360 39794
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 25136 39500 25188 39506
rect 25136 39442 25188 39448
rect 25332 38962 25360 39766
rect 25424 39642 25452 41686
rect 25608 39846 25636 47126
rect 25596 39840 25648 39846
rect 25596 39782 25648 39788
rect 25412 39636 25464 39642
rect 25412 39578 25464 39584
rect 25320 38956 25372 38962
rect 25320 38898 25372 38904
rect 25136 38752 25188 38758
rect 25136 38694 25188 38700
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24688 38010 24716 38150
rect 24676 38004 24728 38010
rect 24676 37946 24728 37952
rect 24860 37936 24912 37942
rect 24780 37884 24860 37890
rect 24780 37878 24912 37884
rect 24780 37862 24900 37878
rect 24780 37126 24808 37862
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 24780 36854 24808 37062
rect 24768 36848 24820 36854
rect 24768 36790 24820 36796
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24504 35494 24532 35634
rect 24780 35494 24808 36790
rect 25148 36718 25176 38694
rect 25332 38321 25360 38898
rect 25700 38729 25728 53382
rect 25792 40390 25820 53926
rect 25964 52624 26016 52630
rect 25964 52566 26016 52572
rect 25872 50720 25924 50726
rect 25872 50662 25924 50668
rect 25780 40384 25832 40390
rect 25780 40326 25832 40332
rect 25884 38826 25912 50662
rect 25976 38894 26004 52566
rect 25964 38888 26016 38894
rect 25964 38830 26016 38836
rect 25872 38820 25924 38826
rect 25872 38762 25924 38768
rect 25686 38720 25742 38729
rect 25686 38655 25742 38664
rect 25318 38312 25374 38321
rect 25318 38247 25374 38256
rect 25318 37496 25374 37505
rect 25228 37460 25280 37466
rect 25318 37431 25374 37440
rect 25228 37402 25280 37408
rect 25136 36712 25188 36718
rect 25136 36654 25188 36660
rect 24492 35488 24544 35494
rect 24492 35430 24544 35436
rect 24768 35488 24820 35494
rect 24768 35430 24820 35436
rect 24504 34950 24532 35430
rect 24492 34944 24544 34950
rect 24492 34886 24544 34892
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24504 33930 24532 34886
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24492 33924 24544 33930
rect 24492 33866 24544 33872
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24492 31136 24544 31142
rect 24492 31078 24544 31084
rect 24308 30388 24360 30394
rect 24308 30330 24360 30336
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 29714 23796 30126
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 23756 29708 23808 29714
rect 23756 29650 23808 29656
rect 23952 29306 23980 29786
rect 24400 29776 24452 29782
rect 24400 29718 24452 29724
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 23572 29096 23624 29102
rect 23572 29038 23624 29044
rect 23400 28104 23520 28132
rect 23400 25906 23428 28104
rect 24136 27713 24164 29106
rect 24216 28484 24268 28490
rect 24216 28426 24268 28432
rect 24122 27704 24178 27713
rect 24228 27674 24256 28426
rect 24122 27639 24178 27648
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 23572 27056 23624 27062
rect 23572 26998 23624 27004
rect 23584 26518 23612 26998
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23860 25906 23888 26726
rect 24216 26376 24268 26382
rect 24216 26318 24268 26324
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23400 25498 23428 25842
rect 23756 25764 23808 25770
rect 23756 25706 23808 25712
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 23400 23050 23428 24550
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23492 23066 23520 23734
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23388 23044 23440 23050
rect 23492 23038 23612 23066
rect 23388 22986 23440 22992
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23294 22808 23350 22817
rect 23294 22743 23350 22752
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22094 23336 22743
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23216 22066 23336 22094
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 23216 21434 23244 22066
rect 23400 22030 23428 22578
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21690 23428 21966
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23492 21570 23520 22918
rect 23584 22778 23612 23038
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23308 21554 23520 21570
rect 23296 21548 23520 21554
rect 23348 21542 23520 21548
rect 23296 21490 23348 21496
rect 22468 21412 22520 21418
rect 23216 21406 23336 21434
rect 22468 21354 22520 21360
rect 22480 17270 22508 21354
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20398 23336 21406
rect 23386 21176 23442 21185
rect 23386 21111 23442 21120
rect 23400 20534 23428 21111
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23584 19446 23612 21626
rect 23676 21622 23704 23462
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22572 17882 22600 18634
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 22744 18148 22796 18154
rect 22744 18090 22796 18096
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22388 16374 22508 16402
rect 22480 16114 22508 16374
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22388 15162 22416 16050
rect 22572 16046 22600 17818
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22020 12238 22048 12718
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22020 7410 22048 8366
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22204 6914 22232 13738
rect 22296 13190 22324 14350
rect 22664 13326 22692 17002
rect 22756 14006 22784 18090
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23400 17921 23428 18158
rect 23386 17912 23442 17921
rect 23386 17847 23442 17856
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12918 22324 13126
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 7426 22324 9318
rect 22388 8090 22416 11698
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 22296 7398 22416 7426
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 21744 6886 21864 6914
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21744 2854 21772 6190
rect 21836 5234 21864 6886
rect 22112 6886 22232 6914
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21638 2408 21694 2417
rect 21638 2343 21694 2352
rect 21928 800 21956 6190
rect 22020 3398 22048 6666
rect 22112 4146 22140 6886
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22098 4040 22154 4049
rect 22098 3975 22100 3984
rect 22152 3975 22154 3984
rect 22100 3946 22152 3952
rect 22204 3942 22232 6258
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22296 800 22324 7278
rect 22388 6934 22416 7398
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22480 5710 22508 10134
rect 22572 9042 22600 12582
rect 22664 11898 22692 12854
rect 23308 12850 23336 17002
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23400 14618 23428 16594
rect 23676 15026 23704 19722
rect 23768 17202 23796 25706
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23846 23624 23902 23633
rect 23846 23559 23902 23568
rect 23860 23118 23888 23559
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23952 18290 23980 25094
rect 24044 20466 24072 25094
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23860 17338 23888 17614
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23860 16794 23888 17274
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 24136 16114 24164 21966
rect 24228 20466 24256 26318
rect 24412 24206 24440 29718
rect 24504 26314 24532 31078
rect 24596 29238 24624 33798
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24596 27130 24624 28358
rect 24688 28150 24716 34682
rect 24780 30666 24808 34886
rect 25240 33658 25268 37402
rect 25332 37262 25360 37431
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25332 36689 25360 36722
rect 25318 36680 25374 36689
rect 25318 36615 25374 36624
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25332 35873 25360 36110
rect 25318 35864 25374 35873
rect 25318 35799 25374 35808
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 35086 25360 35430
rect 25320 35080 25372 35086
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25320 34176
rect 25372 34167 25374 34176
rect 25320 34138 25372 34144
rect 25228 33652 25280 33658
rect 25228 33594 25280 33600
rect 25410 33416 25466 33425
rect 25410 33351 25466 33360
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 32609 25360 32846
rect 25318 32600 25374 32609
rect 25318 32535 25374 32544
rect 25424 32434 25452 33351
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25320 31340 25372 31346
rect 25320 31282 25372 31288
rect 25332 30977 25360 31282
rect 25318 30968 25374 30977
rect 25318 30903 25320 30912
rect 25372 30903 25374 30912
rect 25320 30874 25372 30880
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 24768 30660 24820 30666
rect 24768 30602 24820 30608
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24858 28520 24914 28529
rect 24858 28455 24860 28464
rect 24912 28455 24914 28464
rect 24860 28426 24912 28432
rect 24676 28144 24728 28150
rect 24676 28086 24728 28092
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24584 27124 24636 27130
rect 24584 27066 24636 27072
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24596 26586 24624 26726
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24584 26444 24636 26450
rect 24584 26386 24636 26392
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24504 23798 24532 24822
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 24320 22098 24348 23530
rect 24504 22778 24532 23734
rect 24596 23610 24624 26386
rect 24688 24750 24716 27950
rect 24964 27062 24992 30534
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25332 29306 25360 29582
rect 25516 29345 25544 30670
rect 25502 29336 25558 29345
rect 25320 29300 25372 29306
rect 25502 29271 25504 29280
rect 25320 29242 25372 29248
rect 25556 29271 25558 29280
rect 25504 29242 25556 29248
rect 25136 27940 25188 27946
rect 25136 27882 25188 27888
rect 25044 27396 25096 27402
rect 25044 27338 25096 27344
rect 24952 27056 25004 27062
rect 24952 26998 25004 27004
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 24688 24342 24716 24686
rect 24858 24440 24914 24449
rect 24858 24375 24914 24384
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24872 24274 24900 24375
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24964 24138 24992 25366
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24596 23582 24716 23610
rect 24688 23526 24716 23582
rect 24676 23520 24728 23526
rect 24676 23462 24728 23468
rect 24688 23254 24716 23462
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24858 21992 24914 22001
rect 24858 21927 24914 21936
rect 24872 21010 24900 21927
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24766 19544 24822 19553
rect 24766 19479 24822 19488
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18970 24440 19110
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24412 18698 24440 18906
rect 24674 18728 24730 18737
rect 24400 18692 24452 18698
rect 24674 18663 24730 18672
rect 24400 18634 24452 18640
rect 24412 17882 24440 18634
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22756 9994 22784 12106
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22848 9586 22876 12310
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23296 10464 23348 10470
rect 23296 10406 23348 10412
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22468 5704 22520 5710
rect 22468 5646 22520 5652
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22480 2922 22508 5102
rect 22572 3233 22600 8366
rect 22664 7018 22692 9046
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22848 7290 22876 8774
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23308 7410 23336 10406
rect 23400 8974 23428 14010
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 22848 7262 23336 7290
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22664 6990 22876 7018
rect 22744 6928 22796 6934
rect 22744 6870 22796 6876
rect 22756 4622 22784 6870
rect 22848 6798 22876 6990
rect 22836 6792 22888 6798
rect 22836 6734 22888 6740
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 23308 4554 23336 7262
rect 23400 4865 23428 7890
rect 23492 7886 23520 8774
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23386 4856 23442 4865
rect 23386 4791 23442 4800
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22558 3224 22614 3233
rect 22558 3159 22614 3168
rect 22468 2916 22520 2922
rect 22468 2858 22520 2864
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 22664 800 22692 2790
rect 22848 2530 22876 3334
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22848 2502 23060 2530
rect 23032 800 23060 2502
rect 23400 800 23428 2926
rect 23768 800 23796 13806
rect 23860 10674 23888 15914
rect 24228 15502 24256 17478
rect 24688 17134 24716 18663
rect 24780 18222 24808 19479
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24872 17678 24900 20810
rect 24950 20360 25006 20369
rect 24950 20295 25006 20304
rect 24964 19922 24992 20295
rect 24952 19916 25004 19922
rect 24952 19858 25004 19864
rect 25056 19854 25084 27338
rect 25148 25974 25176 27882
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25240 26518 25268 27270
rect 25502 26888 25558 26897
rect 25502 26823 25558 26832
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25136 25968 25188 25974
rect 25136 25910 25188 25916
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25240 25498 25268 26454
rect 25318 26072 25374 26081
rect 25318 26007 25374 26016
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25240 24886 25268 25434
rect 25228 24880 25280 24886
rect 25228 24822 25280 24828
rect 25134 24712 25190 24721
rect 25134 24647 25136 24656
rect 25188 24647 25190 24656
rect 25136 24618 25188 24624
rect 25332 23730 25360 26007
rect 25412 25968 25464 25974
rect 25412 25910 25464 25916
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25332 22778 25360 23666
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25424 20942 25452 25910
rect 25516 25498 25544 26823
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25516 24818 25544 25434
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24766 17096 24822 17105
rect 24766 17031 24822 17040
rect 24674 16280 24730 16289
rect 24674 16215 24730 16224
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24688 14958 24716 16215
rect 24780 16046 24808 17031
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 26054 15464 26110 15473
rect 26054 15399 26056 15408
rect 26108 15399 26110 15408
rect 26056 15370 26108 15376
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 25134 14648 25190 14657
rect 25134 14583 25190 14592
rect 25148 14006 25176 14583
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24780 12782 24808 13767
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25148 13025 25176 13194
rect 25134 13016 25190 13025
rect 25134 12951 25190 12960
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24766 12200 24822 12209
rect 24766 12135 24822 12144
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23952 8498 23980 11018
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 24044 5234 24072 9862
rect 24136 6798 24164 12038
rect 24674 11384 24730 11393
rect 24674 11319 24730 11328
rect 24582 10568 24638 10577
rect 24582 10503 24638 10512
rect 24596 8430 24624 10503
rect 24688 9518 24716 11319
rect 24780 10606 24808 12135
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9761 24992 9998
rect 24950 9752 25006 9761
rect 24950 9687 25006 9696
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24582 8120 24638 8129
rect 24582 8055 24638 8064
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 24596 6254 24624 8055
rect 24688 7342 24716 8871
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24766 7304 24822 7313
rect 24766 7239 24822 7248
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24688 4146 24716 6598
rect 24780 5166 24808 7239
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24872 4758 24900 8298
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6497 24992 6666
rect 24950 6488 25006 6497
rect 24950 6423 25006 6432
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24136 2854 24164 3402
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 24136 800 24164 2790
rect 24596 2446 24624 3334
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24872 1601 24900 2450
rect 24858 1592 24914 1601
rect 24858 1527 24914 1536
rect 19444 734 19656 762
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 24964 785 24992 3606
rect 25056 3194 25084 7822
rect 25134 5672 25190 5681
rect 25134 5607 25190 5616
rect 25148 4214 25176 5607
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 25332 2650 25360 2994
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 24950 776 25006 785
rect 24950 711 25006 720
<< via2 >>
rect 1306 52944 1362 53000
rect 1306 50496 1362 50552
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 3974 55392 4030 55448
rect 1306 48068 1362 48104
rect 1306 48048 1308 48068
rect 1308 48048 1360 48068
rect 1360 48048 1362 48068
rect 1306 45620 1362 45656
rect 1306 45600 1308 45620
rect 1308 45600 1360 45620
rect 1360 45600 1362 45620
rect 1306 43152 1362 43208
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 1306 40704 1362 40760
rect 1306 38292 1308 38312
rect 1308 38292 1360 38312
rect 1360 38292 1362 38312
rect 1306 38256 1362 38292
rect 1306 33360 1362 33416
rect 1306 30912 1362 30968
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 1766 35808 1822 35864
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 1306 28464 1362 28520
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 1306 23604 1308 23624
rect 1308 23604 1360 23624
rect 1360 23604 1362 23624
rect 1306 23568 1362 23604
rect 2778 26016 2834 26072
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 1306 21120 1362 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 1306 18672 1362 18728
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 1306 16224 1362 16280
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 1306 13812 1308 13832
rect 1308 13812 1360 13832
rect 1360 13812 1362 13832
rect 1306 13776 1362 13812
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 1950 8336 2006 8392
rect 1306 1536 1362 1592
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3514 11192 3570 11248
rect 4066 8880 4122 8936
rect 4066 6432 4122 6488
rect 4066 4020 4068 4040
rect 4068 4020 4120 4040
rect 4120 4020 4122 4040
rect 4066 3984 4122 4020
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 8206 38256 8262 38312
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 9494 44260 9550 44296
rect 9494 44240 9496 44260
rect 9496 44240 9548 44260
rect 9548 44240 9550 44260
rect 8758 36216 8814 36272
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 9770 44684 9772 44704
rect 9772 44684 9824 44704
rect 9824 44684 9826 44704
rect 9770 44648 9826 44684
rect 9678 37848 9734 37904
rect 9402 35808 9458 35864
rect 10322 42508 10324 42528
rect 10324 42508 10376 42528
rect 10376 42508 10378 42528
rect 10322 42472 10378 42508
rect 10138 38936 10194 38992
rect 9954 36760 10010 36816
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 11242 38256 11298 38312
rect 9862 24268 9918 24304
rect 9862 24248 9864 24268
rect 9864 24248 9916 24268
rect 9916 24248 9918 24268
rect 8666 19660 8668 19680
rect 8668 19660 8720 19680
rect 8720 19660 8722 19680
rect 8666 19624 8722 19660
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 8942 16088 8998 16144
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 8206 4120 8262 4176
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 10414 22888 10470 22944
rect 11518 38700 11520 38720
rect 11520 38700 11572 38720
rect 11572 38700 11574 38720
rect 11518 38664 11574 38700
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 14002 52536 14058 52592
rect 14462 52536 14518 52592
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 11886 37304 11942 37360
rect 12254 39092 12310 39128
rect 12254 39072 12256 39092
rect 12256 39072 12308 39092
rect 12308 39072 12310 39092
rect 12346 38664 12402 38720
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12346 37168 12402 37224
rect 11426 30676 11428 30696
rect 11428 30676 11480 30696
rect 11480 30676 11482 30696
rect 11426 30640 11482 30676
rect 12438 36080 12494 36136
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12990 39092 13046 39128
rect 12990 39072 12992 39092
rect 12992 39072 13044 39092
rect 13044 39072 13046 39092
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 13266 38004 13322 38040
rect 13266 37984 13268 38004
rect 13268 37984 13320 38004
rect 13320 37984 13322 38004
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12438 33360 12494 33416
rect 12254 32308 12256 32328
rect 12256 32308 12308 32328
rect 12308 32308 12310 32328
rect 12254 32272 12310 32308
rect 10782 22888 10838 22944
rect 9586 5616 9642 5672
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 9862 5480 9918 5536
rect 12530 26288 12586 26344
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 13818 38256 13874 38312
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 11978 19488 12034 19544
rect 12162 19352 12218 19408
rect 12990 24692 12992 24712
rect 12992 24692 13044 24712
rect 13044 24692 13046 24712
rect 12990 24656 13046 24692
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 14278 38412 14334 38448
rect 14278 38392 14280 38412
rect 14280 38392 14332 38412
rect 14332 38392 14334 38412
rect 14278 37304 14334 37360
rect 14186 35808 14242 35864
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12898 19896 12954 19952
rect 12898 19216 12954 19272
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 14370 32544 14426 32600
rect 14738 33224 14794 33280
rect 14370 30252 14426 30288
rect 14370 30232 14372 30252
rect 14372 30232 14424 30252
rect 14424 30232 14426 30252
rect 13910 24656 13966 24712
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12806 13912 12862 13968
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 17038 53932 17040 53952
rect 17040 53932 17092 53952
rect 17092 53932 17094 53952
rect 17038 53896 17094 53932
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 16394 52536 16450 52592
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 15566 35672 15622 35728
rect 15290 30640 15346 30696
rect 13726 18128 13782 18184
rect 15290 28364 15292 28384
rect 15292 28364 15344 28384
rect 15344 28364 15346 28384
rect 15290 28328 15346 28364
rect 14646 21664 14702 21720
rect 14830 19660 14832 19680
rect 14832 19660 14884 19680
rect 14884 19660 14886 19680
rect 14830 19624 14886 19660
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14738 16244 14794 16280
rect 14738 16224 14740 16244
rect 14740 16224 14792 16244
rect 14792 16224 14794 16244
rect 15934 40024 15990 40080
rect 15842 36660 15844 36680
rect 15844 36660 15896 36680
rect 15896 36660 15898 36680
rect 15842 36624 15898 36660
rect 15750 36236 15806 36272
rect 15750 36216 15752 36236
rect 15752 36216 15804 36236
rect 15804 36216 15806 36236
rect 15290 19352 15346 19408
rect 15842 28212 15898 28248
rect 15842 28192 15844 28212
rect 15844 28192 15896 28212
rect 15896 28192 15898 28212
rect 16670 41520 16726 41576
rect 16394 37732 16450 37768
rect 16394 37712 16396 37732
rect 16396 37712 16448 37732
rect 16448 37712 16450 37732
rect 16118 33260 16120 33280
rect 16120 33260 16172 33280
rect 16172 33260 16174 33280
rect 16118 33224 16174 33260
rect 16670 36780 16726 36816
rect 16670 36760 16672 36780
rect 16672 36760 16724 36780
rect 16724 36760 16726 36780
rect 17038 37848 17094 37904
rect 17406 37984 17462 38040
rect 17130 33224 17186 33280
rect 16026 27956 16028 27976
rect 16028 27956 16080 27976
rect 16080 27956 16082 27976
rect 16026 27920 16082 27956
rect 16394 29688 16450 29744
rect 16394 29044 16396 29064
rect 16396 29044 16448 29064
rect 16448 29044 16450 29064
rect 16394 29008 16450 29044
rect 16394 24248 16450 24304
rect 16854 24656 16910 24712
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17590 38664 17646 38720
rect 17590 38392 17646 38448
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 18234 40024 18290 40080
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17866 38936 17922 38992
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 18418 38836 18420 38856
rect 18420 38836 18472 38856
rect 18472 38836 18474 38856
rect 18418 38800 18474 38836
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 18326 33088 18382 33144
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 15750 16768 15806 16824
rect 15934 16224 15990 16280
rect 16026 12960 16082 13016
rect 16210 12552 16266 12608
rect 17314 20596 17370 20632
rect 17314 20576 17316 20596
rect 17316 20576 17368 20596
rect 17368 20576 17370 20596
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 20074 45772 20076 45792
rect 20076 45772 20128 45792
rect 20128 45772 20130 45792
rect 19246 41556 19248 41576
rect 19248 41556 19300 41576
rect 19300 41556 19302 41576
rect 19246 41520 19302 41556
rect 18050 28600 18106 28656
rect 18326 28464 18382 28520
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 18234 27512 18290 27568
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 18602 27376 18658 27432
rect 18602 26016 18658 26072
rect 20074 45736 20130 45772
rect 19246 37440 19302 37496
rect 19246 35692 19302 35728
rect 19246 35672 19248 35692
rect 19248 35672 19300 35692
rect 19300 35672 19302 35692
rect 19798 37732 19854 37768
rect 19798 37712 19800 37732
rect 19800 37712 19852 37732
rect 19852 37712 19854 37732
rect 19430 31900 19432 31920
rect 19432 31900 19484 31920
rect 19484 31900 19486 31920
rect 19430 31864 19486 31900
rect 18786 27512 18842 27568
rect 18786 27376 18842 27432
rect 18602 25744 18658 25800
rect 18510 24656 18566 24712
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17498 11892 17554 11928
rect 17498 11872 17500 11892
rect 17500 11872 17552 11892
rect 17552 11872 17554 11892
rect 18510 20576 18566 20632
rect 17866 19896 17922 19952
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18602 19352 18658 19408
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 20626 46960 20682 47016
rect 20074 31476 20130 31512
rect 20074 31456 20076 31476
rect 20076 31456 20128 31476
rect 20128 31456 20130 31476
rect 20442 38664 20498 38720
rect 20166 28212 20222 28248
rect 20166 28192 20168 28212
rect 20168 28192 20220 28212
rect 20220 28192 20222 28212
rect 19522 24928 19578 24984
rect 19890 24948 19946 24984
rect 19890 24928 19892 24948
rect 19892 24928 19944 24948
rect 19944 24928 19946 24948
rect 20442 30932 20498 30968
rect 21454 46980 21510 47016
rect 21454 46960 21456 46980
rect 21456 46960 21508 46980
rect 21508 46960 21510 46980
rect 21086 38800 21142 38856
rect 22282 53932 22284 53952
rect 22284 53932 22336 53952
rect 22336 53932 22338 53952
rect 22282 53896 22338 53932
rect 21914 46316 21916 46336
rect 21916 46316 21968 46336
rect 21968 46316 21970 46336
rect 21914 46280 21970 46316
rect 21638 43288 21694 43344
rect 20626 32308 20628 32328
rect 20628 32308 20680 32328
rect 20680 32308 20682 32328
rect 20626 32272 20682 32308
rect 20442 30912 20444 30932
rect 20444 30912 20496 30932
rect 20496 30912 20498 30932
rect 23386 56072 23442 56128
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 24490 55392 24546 55448
rect 24766 54576 24822 54632
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22006 40704 22062 40760
rect 22190 41656 22246 41712
rect 22466 41520 22522 41576
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 21178 32272 21234 32328
rect 21638 32716 21640 32736
rect 21640 32716 21692 32736
rect 21692 32716 21694 32736
rect 21638 32680 21694 32716
rect 21822 32564 21878 32600
rect 21822 32544 21824 32564
rect 21824 32544 21876 32564
rect 21876 32544 21878 32564
rect 21730 32272 21786 32328
rect 20166 20712 20222 20768
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19430 13404 19432 13424
rect 19432 13404 19484 13424
rect 19484 13404 19486 13424
rect 19430 13368 19486 13404
rect 18786 3984 18842 4040
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22466 36624 22522 36680
rect 22466 36216 22522 36272
rect 22374 34312 22430 34368
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 23110 42336 23166 42392
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22926 41656 22982 41712
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22558 32716 22560 32736
rect 22560 32716 22612 32736
rect 22612 32716 22614 32736
rect 22558 32680 22614 32716
rect 23570 38528 23626 38584
rect 23202 37868 23258 37904
rect 23202 37848 23204 37868
rect 23204 37848 23256 37868
rect 23256 37848 23258 37868
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22926 36216 22982 36272
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 24950 53760 25006 53816
rect 25318 53760 25374 53816
rect 25042 52944 25098 53000
rect 24766 52128 24822 52184
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 21270 13368 21326 13424
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 24766 46416 24822 46472
rect 24858 45600 24914 45656
rect 25502 51348 25504 51368
rect 25504 51348 25556 51368
rect 25556 51348 25558 51368
rect 25502 51312 25558 51348
rect 25226 51040 25282 51096
rect 25042 50496 25098 50552
rect 25318 49680 25374 49736
rect 25318 48864 25374 48920
rect 25318 48084 25320 48104
rect 25320 48084 25372 48104
rect 25372 48084 25374 48104
rect 25318 48048 25374 48084
rect 25502 47232 25558 47288
rect 24766 44276 24768 44296
rect 24768 44276 24820 44296
rect 24820 44276 24822 44296
rect 24766 44240 24822 44276
rect 25502 44784 25558 44840
rect 25502 43968 25558 44024
rect 25318 43152 25374 43208
rect 24858 42336 24914 42392
rect 24858 39072 24914 39128
rect 25318 41556 25320 41576
rect 25320 41556 25372 41576
rect 25372 41556 25374 41576
rect 25318 41520 25374 41556
rect 25318 40704 25374 40760
rect 25318 39888 25374 39944
rect 25686 38664 25742 38720
rect 25318 38256 25374 38312
rect 25318 37440 25374 37496
rect 24122 27648 24178 27704
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 23294 22752 23350 22808
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23386 21120 23442 21176
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23386 17856 23442 17912
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 21638 2352 21694 2408
rect 22098 4004 22154 4040
rect 22098 3984 22100 4004
rect 22100 3984 22152 4004
rect 22152 3984 22154 4004
rect 23846 23568 23902 23624
rect 25318 36624 25374 36680
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34196 25374 34232
rect 25318 34176 25320 34196
rect 25320 34176 25372 34196
rect 25372 34176 25374 34196
rect 25410 33360 25466 33416
rect 25318 32544 25374 32600
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30932 25374 30968
rect 25318 30912 25320 30932
rect 25320 30912 25372 30932
rect 25372 30912 25374 30932
rect 24858 28484 24914 28520
rect 24858 28464 24860 28484
rect 24860 28464 24912 28484
rect 24912 28464 24914 28484
rect 25318 30096 25374 30152
rect 25502 29300 25558 29336
rect 25502 29280 25504 29300
rect 25504 29280 25556 29300
rect 25556 29280 25558 29300
rect 24858 24384 24914 24440
rect 24858 21936 24914 21992
rect 24766 19488 24822 19544
rect 24674 18672 24730 18728
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 23386 4800 23442 4856
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22558 3168 22614 3224
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 24950 20304 25006 20360
rect 25502 26832 25558 26888
rect 25318 26016 25374 26072
rect 25134 25200 25190 25256
rect 25134 24676 25190 24712
rect 25134 24656 25136 24676
rect 25136 24656 25188 24676
rect 25188 24656 25190 24676
rect 24766 17040 24822 17096
rect 24674 16224 24730 16280
rect 26054 15428 26110 15464
rect 26054 15408 26056 15428
rect 26056 15408 26108 15428
rect 26108 15408 26110 15428
rect 25134 14592 25190 14648
rect 24766 13776 24822 13832
rect 25134 12960 25190 13016
rect 24766 12144 24822 12200
rect 24674 11328 24730 11384
rect 24582 10512 24638 10568
rect 24950 9696 25006 9752
rect 24674 8880 24730 8936
rect 24582 8064 24638 8120
rect 24766 7248 24822 7304
rect 24950 6432 25006 6488
rect 24858 1536 24914 1592
rect 25134 5616 25190 5672
rect 24950 720 25006 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 0 55450 800 55480
rect 3969 55450 4035 55453
rect 0 55448 4035 55450
rect 0 55392 3974 55448
rect 4030 55392 4035 55448
rect 0 55390 4035 55392
rect 0 55360 800 55390
rect 3969 55387 4035 55390
rect 24485 55450 24551 55453
rect 26200 55450 27000 55480
rect 24485 55448 27000 55450
rect 24485 55392 24490 55448
rect 24546 55392 27000 55448
rect 24485 55390 27000 55392
rect 24485 55387 24551 55390
rect 26200 55360 27000 55390
rect 24761 54634 24827 54637
rect 26200 54634 27000 54664
rect 24761 54632 27000 54634
rect 24761 54576 24766 54632
rect 24822 54576 27000 54632
rect 24761 54574 27000 54576
rect 24761 54571 24827 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 17033 53954 17099 53957
rect 17166 53954 17172 53956
rect 17033 53952 17172 53954
rect 17033 53896 17038 53952
rect 17094 53896 17172 53952
rect 17033 53894 17172 53896
rect 17033 53891 17099 53894
rect 17166 53892 17172 53894
rect 17236 53892 17242 53956
rect 21950 53892 21956 53956
rect 22020 53954 22026 53956
rect 22277 53954 22343 53957
rect 22020 53952 22343 53954
rect 22020 53896 22282 53952
rect 22338 53896 22343 53952
rect 22020 53894 22343 53896
rect 22020 53892 22026 53894
rect 22277 53891 22343 53894
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 24945 53818 25011 53821
rect 25313 53818 25379 53821
rect 26200 53818 27000 53848
rect 24945 53816 27000 53818
rect 24945 53760 24950 53816
rect 25006 53760 25318 53816
rect 25374 53760 27000 53816
rect 24945 53758 27000 53760
rect 24945 53755 25011 53758
rect 25313 53755 25379 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 0 53002 800 53032
rect 1301 53002 1367 53005
rect 0 53000 1367 53002
rect 0 52944 1306 53000
rect 1362 52944 1367 53000
rect 0 52942 1367 52944
rect 0 52912 800 52942
rect 1301 52939 1367 52942
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 13997 52596 14063 52597
rect 13997 52592 14044 52596
rect 14108 52594 14114 52596
rect 14457 52594 14523 52597
rect 16389 52596 16455 52597
rect 14590 52594 14596 52596
rect 13997 52536 14002 52592
rect 13997 52532 14044 52536
rect 14108 52534 14154 52594
rect 14457 52592 14596 52594
rect 14457 52536 14462 52592
rect 14518 52536 14596 52592
rect 14457 52534 14596 52536
rect 14108 52532 14114 52534
rect 13997 52531 14063 52532
rect 14457 52531 14523 52534
rect 14590 52532 14596 52534
rect 14660 52532 14666 52596
rect 16389 52592 16436 52596
rect 16500 52594 16506 52596
rect 16389 52536 16394 52592
rect 16389 52532 16436 52536
rect 16500 52534 16546 52594
rect 16500 52532 16506 52534
rect 16389 52531 16455 52532
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24761 52186 24827 52189
rect 26200 52186 27000 52216
rect 24761 52184 27000 52186
rect 24761 52128 24766 52184
rect 24822 52128 27000 52184
rect 24761 52126 27000 52128
rect 24761 52123 24827 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 25497 51370 25563 51373
rect 26200 51370 27000 51400
rect 25497 51368 27000 51370
rect 25497 51312 25502 51368
rect 25558 51312 27000 51368
rect 25497 51310 27000 51312
rect 25497 51307 25563 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 22318 51036 22324 51100
rect 22388 51098 22394 51100
rect 25221 51098 25287 51101
rect 22388 51096 25287 51098
rect 22388 51040 25226 51096
rect 25282 51040 25287 51096
rect 22388 51038 25287 51040
rect 22388 51036 22394 51038
rect 25221 51035 25287 51038
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 1301 50554 1367 50557
rect 0 50552 1367 50554
rect 0 50496 1306 50552
rect 1362 50496 1367 50552
rect 0 50494 1367 50496
rect 0 50464 800 50494
rect 1301 50491 1367 50494
rect 25037 50554 25103 50557
rect 26200 50554 27000 50584
rect 25037 50552 27000 50554
rect 25037 50496 25042 50552
rect 25098 50496 27000 50552
rect 25037 50494 27000 50496
rect 25037 50491 25103 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25313 49738 25379 49741
rect 26200 49738 27000 49768
rect 25313 49736 27000 49738
rect 25313 49680 25318 49736
rect 25374 49680 27000 49736
rect 25313 49678 27000 49680
rect 25313 49675 25379 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25313 48922 25379 48925
rect 26200 48922 27000 48952
rect 25313 48920 27000 48922
rect 25313 48864 25318 48920
rect 25374 48864 27000 48920
rect 25313 48862 27000 48864
rect 25313 48859 25379 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 25313 48106 25379 48109
rect 26200 48106 27000 48136
rect 25313 48104 27000 48106
rect 25313 48048 25318 48104
rect 25374 48048 27000 48104
rect 25313 48046 27000 48048
rect 25313 48043 25379 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25497 47290 25563 47293
rect 26200 47290 27000 47320
rect 25497 47288 27000 47290
rect 25497 47232 25502 47288
rect 25558 47232 27000 47288
rect 25497 47230 27000 47232
rect 25497 47227 25563 47230
rect 26200 47200 27000 47230
rect 20294 46956 20300 47020
rect 20364 47018 20370 47020
rect 20621 47018 20687 47021
rect 21449 47018 21515 47021
rect 20364 47016 21515 47018
rect 20364 46960 20626 47016
rect 20682 46960 21454 47016
rect 21510 46960 21515 47016
rect 20364 46958 21515 46960
rect 20364 46956 20370 46958
rect 20621 46955 20687 46958
rect 21449 46955 21515 46958
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 24761 46474 24827 46477
rect 26200 46474 27000 46504
rect 24761 46472 27000 46474
rect 24761 46416 24766 46472
rect 24822 46416 27000 46472
rect 24761 46414 27000 46416
rect 24761 46411 24827 46414
rect 26200 46384 27000 46414
rect 21766 46276 21772 46340
rect 21836 46338 21842 46340
rect 21909 46338 21975 46341
rect 21836 46336 21975 46338
rect 21836 46280 21914 46336
rect 21970 46280 21975 46336
rect 21836 46278 21975 46280
rect 21836 46276 21842 46278
rect 21909 46275 21975 46278
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 20069 45796 20135 45797
rect 20069 45794 20116 45796
rect 20024 45792 20116 45794
rect 20024 45736 20074 45792
rect 20024 45734 20116 45736
rect 20069 45732 20116 45734
rect 20180 45732 20186 45796
rect 20069 45731 20135 45732
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 24853 45658 24919 45661
rect 26200 45658 27000 45688
rect 24853 45656 27000 45658
rect 24853 45600 24858 45656
rect 24914 45600 27000 45656
rect 24853 45598 27000 45600
rect 24853 45595 24919 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25497 44842 25563 44845
rect 26200 44842 27000 44872
rect 25497 44840 27000 44842
rect 25497 44784 25502 44840
rect 25558 44784 27000 44840
rect 25497 44782 27000 44784
rect 25497 44779 25563 44782
rect 26200 44752 27000 44782
rect 9765 44708 9831 44709
rect 9765 44706 9812 44708
rect 9720 44704 9812 44706
rect 9720 44648 9770 44704
rect 9720 44646 9812 44648
rect 9765 44644 9812 44646
rect 9876 44644 9882 44708
rect 9765 44643 9831 44644
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 9489 44298 9555 44301
rect 12198 44298 12204 44300
rect 9489 44296 12204 44298
rect 9489 44240 9494 44296
rect 9550 44240 12204 44296
rect 9489 44238 12204 44240
rect 9489 44235 9555 44238
rect 12198 44236 12204 44238
rect 12268 44236 12274 44300
rect 23422 44236 23428 44300
rect 23492 44298 23498 44300
rect 24761 44298 24827 44301
rect 23492 44296 24827 44298
rect 23492 44240 24766 44296
rect 24822 44240 24827 44296
rect 23492 44238 24827 44240
rect 23492 44236 23498 44238
rect 24761 44235 24827 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 25497 44026 25563 44029
rect 26200 44026 27000 44056
rect 25497 44024 27000 44026
rect 25497 43968 25502 44024
rect 25558 43968 27000 44024
rect 25497 43966 27000 43968
rect 25497 43963 25563 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 21633 43348 21699 43349
rect 21582 43346 21588 43348
rect 21542 43286 21588 43346
rect 21652 43344 21699 43348
rect 21694 43288 21699 43344
rect 21582 43284 21588 43286
rect 21652 43284 21699 43288
rect 21633 43283 21699 43284
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 25313 43210 25379 43213
rect 26200 43210 27000 43240
rect 25313 43208 27000 43210
rect 25313 43152 25318 43208
rect 25374 43152 27000 43208
rect 25313 43150 27000 43152
rect 25313 43147 25379 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 10317 42530 10383 42533
rect 10910 42530 10916 42532
rect 10317 42528 10916 42530
rect 10317 42472 10322 42528
rect 10378 42472 10916 42528
rect 10317 42470 10916 42472
rect 10317 42467 10383 42470
rect 10910 42468 10916 42470
rect 10980 42468 10986 42532
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 22686 42332 22692 42396
rect 22756 42394 22762 42396
rect 23105 42394 23171 42397
rect 22756 42392 23171 42394
rect 22756 42336 23110 42392
rect 23166 42336 23171 42392
rect 22756 42334 23171 42336
rect 22756 42332 22762 42334
rect 23105 42331 23171 42334
rect 24853 42394 24919 42397
rect 26200 42394 27000 42424
rect 24853 42392 27000 42394
rect 24853 42336 24858 42392
rect 24914 42336 27000 42392
rect 24853 42334 27000 42336
rect 24853 42331 24919 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 22185 41714 22251 41717
rect 22185 41712 22386 41714
rect 22185 41656 22190 41712
rect 22246 41656 22386 41712
rect 22185 41654 22386 41656
rect 22185 41651 22251 41654
rect 16665 41578 16731 41581
rect 19241 41578 19307 41581
rect 16665 41576 19307 41578
rect 16665 41520 16670 41576
rect 16726 41520 19246 41576
rect 19302 41520 19307 41576
rect 16665 41518 19307 41520
rect 22326 41578 22386 41654
rect 22686 41652 22692 41716
rect 22756 41714 22762 41716
rect 22921 41714 22987 41717
rect 22756 41712 22987 41714
rect 22756 41656 22926 41712
rect 22982 41656 22987 41712
rect 22756 41654 22987 41656
rect 22756 41652 22762 41654
rect 22921 41651 22987 41654
rect 22461 41578 22527 41581
rect 22326 41576 22527 41578
rect 22326 41520 22466 41576
rect 22522 41520 22527 41576
rect 22326 41518 22527 41520
rect 16665 41515 16731 41518
rect 19241 41515 19307 41518
rect 22461 41515 22527 41518
rect 25313 41578 25379 41581
rect 26200 41578 27000 41608
rect 25313 41576 27000 41578
rect 25313 41520 25318 41576
rect 25374 41520 27000 41576
rect 25313 41518 27000 41520
rect 25313 41515 25379 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 22001 40762 22067 40765
rect 22318 40762 22324 40764
rect 22001 40760 22324 40762
rect 22001 40704 22006 40760
rect 22062 40704 22324 40760
rect 22001 40702 22324 40704
rect 22001 40699 22067 40702
rect 22318 40700 22324 40702
rect 22388 40700 22394 40764
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 15929 40084 15995 40085
rect 15878 40020 15884 40084
rect 15948 40082 15995 40084
rect 18229 40082 18295 40085
rect 20662 40082 20668 40084
rect 15948 40080 16040 40082
rect 15990 40024 16040 40080
rect 15948 40022 16040 40024
rect 18229 40080 20668 40082
rect 18229 40024 18234 40080
rect 18290 40024 20668 40080
rect 18229 40022 20668 40024
rect 15948 40020 15995 40022
rect 15929 40019 15995 40020
rect 18229 40019 18295 40022
rect 20662 40020 20668 40022
rect 20732 40020 20738 40084
rect 25313 39946 25379 39949
rect 26200 39946 27000 39976
rect 25313 39944 27000 39946
rect 25313 39888 25318 39944
rect 25374 39888 27000 39944
rect 25313 39886 27000 39888
rect 25313 39883 25379 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 12249 39130 12315 39133
rect 12985 39130 13051 39133
rect 12249 39128 13051 39130
rect 12249 39072 12254 39128
rect 12310 39072 12990 39128
rect 13046 39072 13051 39128
rect 12249 39070 13051 39072
rect 12249 39067 12315 39070
rect 12985 39067 13051 39070
rect 24853 39130 24919 39133
rect 26200 39130 27000 39160
rect 24853 39128 27000 39130
rect 24853 39072 24858 39128
rect 24914 39072 27000 39128
rect 24853 39070 27000 39072
rect 24853 39067 24919 39070
rect 26200 39040 27000 39070
rect 10133 38994 10199 38997
rect 17861 38994 17927 38997
rect 10133 38992 17927 38994
rect 10133 38936 10138 38992
rect 10194 38936 17866 38992
rect 17922 38936 17927 38992
rect 10133 38934 17927 38936
rect 10133 38931 10199 38934
rect 17861 38931 17927 38934
rect 18413 38858 18479 38861
rect 18638 38858 18644 38860
rect 18413 38856 18644 38858
rect 18413 38800 18418 38856
rect 18474 38800 18644 38856
rect 18413 38798 18644 38800
rect 18413 38795 18479 38798
rect 18638 38796 18644 38798
rect 18708 38796 18714 38860
rect 21081 38858 21147 38861
rect 21081 38856 23674 38858
rect 21081 38800 21086 38856
rect 21142 38800 23674 38856
rect 21081 38798 23674 38800
rect 21081 38795 21147 38798
rect 11513 38722 11579 38725
rect 12341 38722 12407 38725
rect 11513 38720 12407 38722
rect 11513 38664 11518 38720
rect 11574 38664 12346 38720
rect 12402 38664 12407 38720
rect 11513 38662 12407 38664
rect 11513 38659 11579 38662
rect 12341 38659 12407 38662
rect 17350 38660 17356 38724
rect 17420 38722 17426 38724
rect 17585 38722 17651 38725
rect 20437 38722 20503 38725
rect 17420 38720 20503 38722
rect 17420 38664 17590 38720
rect 17646 38664 20442 38720
rect 20498 38664 20503 38720
rect 17420 38662 20503 38664
rect 17420 38660 17426 38662
rect 17585 38659 17651 38662
rect 20437 38659 20503 38662
rect 23614 38722 23674 38798
rect 25681 38722 25747 38725
rect 23614 38720 25747 38722
rect 23614 38664 25686 38720
rect 25742 38664 25747 38720
rect 23614 38662 25747 38664
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 23614 38589 23674 38662
rect 25681 38659 25747 38662
rect 23565 38584 23674 38589
rect 23565 38528 23570 38584
rect 23626 38528 23674 38584
rect 23565 38526 23674 38528
rect 23565 38523 23631 38526
rect 14273 38450 14339 38453
rect 17585 38450 17651 38453
rect 14273 38448 17651 38450
rect 14273 38392 14278 38448
rect 14334 38392 17590 38448
rect 17646 38392 17651 38448
rect 14273 38390 17651 38392
rect 14273 38387 14339 38390
rect 17585 38387 17651 38390
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 8201 38314 8267 38317
rect 11237 38314 11303 38317
rect 13813 38314 13879 38317
rect 8201 38312 13879 38314
rect 8201 38256 8206 38312
rect 8262 38256 11242 38312
rect 11298 38256 13818 38312
rect 13874 38256 13879 38312
rect 8201 38254 13879 38256
rect 8201 38251 8267 38254
rect 11237 38251 11303 38254
rect 13813 38251 13879 38254
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 13261 38042 13327 38045
rect 17401 38042 17467 38045
rect 13261 38040 17467 38042
rect 13261 37984 13266 38040
rect 13322 37984 17406 38040
rect 17462 37984 17467 38040
rect 13261 37982 17467 37984
rect 13261 37979 13327 37982
rect 17401 37979 17467 37982
rect 9673 37906 9739 37909
rect 17033 37906 17099 37909
rect 9673 37904 17099 37906
rect 9673 37848 9678 37904
rect 9734 37848 17038 37904
rect 17094 37848 17099 37904
rect 9673 37846 17099 37848
rect 9673 37843 9739 37846
rect 17033 37843 17099 37846
rect 22686 37844 22692 37908
rect 22756 37906 22762 37908
rect 23197 37906 23263 37909
rect 22756 37904 23263 37906
rect 22756 37848 23202 37904
rect 23258 37848 23263 37904
rect 22756 37846 23263 37848
rect 22756 37844 22762 37846
rect 23197 37843 23263 37846
rect 12198 37708 12204 37772
rect 12268 37770 12274 37772
rect 16389 37770 16455 37773
rect 12268 37768 16455 37770
rect 12268 37712 16394 37768
rect 16450 37712 16455 37768
rect 12268 37710 16455 37712
rect 12268 37708 12274 37710
rect 16389 37707 16455 37710
rect 19793 37770 19859 37773
rect 20478 37770 20484 37772
rect 19793 37768 20484 37770
rect 19793 37712 19798 37768
rect 19854 37712 20484 37768
rect 19793 37710 20484 37712
rect 19793 37707 19859 37710
rect 20478 37708 20484 37710
rect 20548 37770 20554 37772
rect 23422 37770 23428 37772
rect 20548 37710 23428 37770
rect 20548 37708 20554 37710
rect 23422 37708 23428 37710
rect 23492 37708 23498 37772
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 19241 37498 19307 37501
rect 19198 37496 19307 37498
rect 19198 37440 19246 37496
rect 19302 37440 19307 37496
rect 19198 37435 19307 37440
rect 25313 37498 25379 37501
rect 26200 37498 27000 37528
rect 25313 37496 27000 37498
rect 25313 37440 25318 37496
rect 25374 37440 27000 37496
rect 25313 37438 27000 37440
rect 25313 37435 25379 37438
rect 11881 37362 11947 37365
rect 14273 37362 14339 37365
rect 11881 37360 14339 37362
rect 11881 37304 11886 37360
rect 11942 37304 14278 37360
rect 14334 37304 14339 37360
rect 11881 37302 14339 37304
rect 11881 37299 11947 37302
rect 14273 37299 14339 37302
rect 12341 37226 12407 37229
rect 19198 37226 19258 37435
rect 26200 37408 27000 37438
rect 12341 37224 19258 37226
rect 12341 37168 12346 37224
rect 12402 37168 19258 37224
rect 12341 37166 19258 37168
rect 12341 37163 12407 37166
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 9806 36756 9812 36820
rect 9876 36818 9882 36820
rect 9949 36818 10015 36821
rect 16665 36818 16731 36821
rect 9876 36816 16731 36818
rect 9876 36760 9954 36816
rect 10010 36760 16670 36816
rect 16726 36760 16731 36816
rect 9876 36758 16731 36760
rect 9876 36756 9882 36758
rect 9949 36755 10015 36758
rect 16665 36755 16731 36758
rect 15837 36682 15903 36685
rect 22461 36682 22527 36685
rect 15837 36680 22527 36682
rect 15837 36624 15842 36680
rect 15898 36624 22466 36680
rect 22522 36624 22527 36680
rect 15837 36622 22527 36624
rect 15837 36619 15903 36622
rect 22461 36619 22527 36622
rect 25313 36682 25379 36685
rect 26200 36682 27000 36712
rect 25313 36680 27000 36682
rect 25313 36624 25318 36680
rect 25374 36624 27000 36680
rect 25313 36622 27000 36624
rect 25313 36619 25379 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 8753 36274 8819 36277
rect 15745 36274 15811 36277
rect 8753 36272 15811 36274
rect 8753 36216 8758 36272
rect 8814 36216 15750 36272
rect 15806 36216 15811 36272
rect 8753 36214 15811 36216
rect 8753 36211 8819 36214
rect 15745 36211 15811 36214
rect 22461 36274 22527 36277
rect 22921 36274 22987 36277
rect 22461 36272 22987 36274
rect 22461 36216 22466 36272
rect 22522 36216 22926 36272
rect 22982 36216 22987 36272
rect 22461 36214 22987 36216
rect 22461 36211 22527 36214
rect 22921 36211 22987 36214
rect 12433 36138 12499 36141
rect 12750 36138 12756 36140
rect 12433 36136 12756 36138
rect 12433 36080 12438 36136
rect 12494 36080 12756 36136
rect 12433 36078 12756 36080
rect 12433 36075 12499 36078
rect 12750 36076 12756 36078
rect 12820 36076 12826 36140
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 1761 35866 1827 35869
rect 0 35864 1827 35866
rect 0 35808 1766 35864
rect 1822 35808 1827 35864
rect 0 35806 1827 35808
rect 0 35776 800 35806
rect 1761 35803 1827 35806
rect 9397 35866 9463 35869
rect 14181 35866 14247 35869
rect 9397 35864 14247 35866
rect 9397 35808 9402 35864
rect 9458 35808 14186 35864
rect 14242 35808 14247 35864
rect 9397 35806 14247 35808
rect 9397 35803 9463 35806
rect 14181 35803 14247 35806
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 15561 35730 15627 35733
rect 19241 35730 19307 35733
rect 15561 35728 19307 35730
rect 15561 35672 15566 35728
rect 15622 35672 19246 35728
rect 19302 35672 19307 35728
rect 15561 35670 19307 35672
rect 15561 35667 15627 35670
rect 19241 35667 19307 35670
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 20662 34308 20668 34372
rect 20732 34370 20738 34372
rect 22369 34370 22435 34373
rect 20732 34368 22435 34370
rect 20732 34312 22374 34368
rect 22430 34312 22435 34368
rect 20732 34310 22435 34312
rect 20732 34308 20738 34310
rect 22369 34307 22435 34310
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 0 33418 800 33448
rect 1301 33418 1367 33421
rect 0 33416 1367 33418
rect 0 33360 1306 33416
rect 1362 33360 1367 33416
rect 0 33358 1367 33360
rect 0 33328 800 33358
rect 1301 33355 1367 33358
rect 12198 33356 12204 33420
rect 12268 33418 12274 33420
rect 12433 33418 12499 33421
rect 12268 33416 12499 33418
rect 12268 33360 12438 33416
rect 12494 33360 12499 33416
rect 12268 33358 12499 33360
rect 12268 33356 12274 33358
rect 12433 33355 12499 33358
rect 25405 33418 25471 33421
rect 26200 33418 27000 33448
rect 25405 33416 27000 33418
rect 25405 33360 25410 33416
rect 25466 33360 27000 33416
rect 25405 33358 27000 33360
rect 25405 33355 25471 33358
rect 26200 33328 27000 33358
rect 14733 33282 14799 33285
rect 16113 33282 16179 33285
rect 17125 33282 17191 33285
rect 14733 33280 17191 33282
rect 14733 33224 14738 33280
rect 14794 33224 16118 33280
rect 16174 33224 17130 33280
rect 17186 33224 17191 33280
rect 14733 33222 17191 33224
rect 14733 33219 14799 33222
rect 16113 33219 16179 33222
rect 17125 33219 17191 33222
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 18321 33146 18387 33149
rect 20294 33146 20300 33148
rect 18321 33144 20300 33146
rect 18321 33088 18326 33144
rect 18382 33088 20300 33144
rect 18321 33086 20300 33088
rect 18321 33083 18387 33086
rect 20294 33084 20300 33086
rect 20364 33084 20370 33148
rect 21633 32738 21699 32741
rect 22553 32738 22619 32741
rect 22686 32738 22692 32740
rect 21633 32736 22692 32738
rect 21633 32680 21638 32736
rect 21694 32680 22558 32736
rect 22614 32680 22692 32736
rect 21633 32678 22692 32680
rect 21633 32675 21699 32678
rect 22553 32675 22619 32678
rect 22686 32676 22692 32678
rect 22756 32676 22762 32740
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 14365 32604 14431 32605
rect 14365 32600 14412 32604
rect 14476 32602 14482 32604
rect 21817 32602 21883 32605
rect 21950 32602 21956 32604
rect 14365 32544 14370 32600
rect 14365 32540 14412 32544
rect 14476 32542 14522 32602
rect 21817 32600 21956 32602
rect 21817 32544 21822 32600
rect 21878 32544 21956 32600
rect 21817 32542 21956 32544
rect 14476 32540 14482 32542
rect 14365 32539 14431 32540
rect 21817 32539 21883 32542
rect 21950 32540 21956 32542
rect 22020 32540 22026 32604
rect 25313 32602 25379 32605
rect 26200 32602 27000 32632
rect 25313 32600 27000 32602
rect 25313 32544 25318 32600
rect 25374 32544 27000 32600
rect 25313 32542 27000 32544
rect 25313 32539 25379 32542
rect 26200 32512 27000 32542
rect 12249 32332 12315 32333
rect 12198 32330 12204 32332
rect 12158 32270 12204 32330
rect 12268 32328 12315 32332
rect 12310 32272 12315 32328
rect 12198 32268 12204 32270
rect 12268 32268 12315 32272
rect 12249 32267 12315 32268
rect 20621 32330 20687 32333
rect 21173 32330 21239 32333
rect 21725 32330 21791 32333
rect 20621 32328 21791 32330
rect 20621 32272 20626 32328
rect 20682 32272 21178 32328
rect 21234 32272 21730 32328
rect 21786 32272 21791 32328
rect 20621 32270 21791 32272
rect 20621 32267 20687 32270
rect 21173 32267 21239 32270
rect 21725 32267 21791 32270
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 19425 31922 19491 31925
rect 19558 31922 19564 31924
rect 19425 31920 19564 31922
rect 19425 31864 19430 31920
rect 19486 31864 19564 31920
rect 19425 31862 19564 31864
rect 19425 31859 19491 31862
rect 19558 31860 19564 31862
rect 19628 31860 19634 31924
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 20069 31516 20135 31517
rect 20069 31512 20116 31516
rect 20180 31514 20186 31516
rect 20069 31456 20074 31512
rect 20069 31452 20116 31456
rect 20180 31454 20226 31514
rect 20180 31452 20186 31454
rect 20069 31451 20135 31452
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 1301 30970 1367 30973
rect 20437 30972 20503 30973
rect 20437 30970 20484 30972
rect 0 30968 1367 30970
rect 0 30912 1306 30968
rect 1362 30912 1367 30968
rect 0 30910 1367 30912
rect 20392 30968 20484 30970
rect 20392 30912 20442 30968
rect 20392 30910 20484 30912
rect 0 30880 800 30910
rect 1301 30907 1367 30910
rect 20437 30908 20484 30910
rect 20548 30908 20554 30972
rect 25313 30970 25379 30973
rect 26200 30970 27000 31000
rect 25313 30968 27000 30970
rect 25313 30912 25318 30968
rect 25374 30912 27000 30968
rect 25313 30910 27000 30912
rect 20437 30907 20503 30908
rect 25313 30907 25379 30910
rect 26200 30880 27000 30910
rect 10174 30636 10180 30700
rect 10244 30698 10250 30700
rect 11421 30698 11487 30701
rect 10244 30696 11487 30698
rect 10244 30640 11426 30696
rect 11482 30640 11487 30696
rect 10244 30638 11487 30640
rect 10244 30636 10250 30638
rect 11421 30635 11487 30638
rect 14038 30636 14044 30700
rect 14108 30698 14114 30700
rect 15285 30698 15351 30701
rect 14108 30696 15351 30698
rect 14108 30640 15290 30696
rect 15346 30640 15351 30696
rect 14108 30638 15351 30640
rect 14108 30636 14114 30638
rect 15285 30635 15351 30638
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 14365 30290 14431 30293
rect 14590 30290 14596 30292
rect 14365 30288 14596 30290
rect 14365 30232 14370 30288
rect 14426 30232 14596 30288
rect 14365 30230 14596 30232
rect 14365 30227 14431 30230
rect 14590 30228 14596 30230
rect 14660 30228 14666 30292
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 16389 29748 16455 29749
rect 16389 29744 16436 29748
rect 16500 29746 16506 29748
rect 16389 29688 16394 29744
rect 16389 29684 16436 29688
rect 16500 29686 16546 29746
rect 16500 29684 16506 29686
rect 16389 29683 16455 29684
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 25497 29338 25563 29341
rect 26200 29338 27000 29368
rect 25497 29336 27000 29338
rect 25497 29280 25502 29336
rect 25558 29280 27000 29336
rect 25497 29278 27000 29280
rect 25497 29275 25563 29278
rect 26200 29248 27000 29278
rect 16062 29004 16068 29068
rect 16132 29066 16138 29068
rect 16389 29066 16455 29069
rect 16132 29064 16455 29066
rect 16132 29008 16394 29064
rect 16450 29008 16455 29064
rect 16132 29006 16455 29008
rect 16132 29004 16138 29006
rect 16389 29003 16455 29006
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 18045 28658 18111 28661
rect 19190 28658 19196 28660
rect 18045 28656 19196 28658
rect 18045 28600 18050 28656
rect 18106 28600 19196 28656
rect 18045 28598 19196 28600
rect 18045 28595 18111 28598
rect 19190 28596 19196 28598
rect 19260 28596 19266 28660
rect 0 28522 800 28552
rect 1301 28522 1367 28525
rect 0 28520 1367 28522
rect 0 28464 1306 28520
rect 1362 28464 1367 28520
rect 0 28462 1367 28464
rect 0 28432 800 28462
rect 1301 28459 1367 28462
rect 18321 28522 18387 28525
rect 21582 28522 21588 28524
rect 18321 28520 21588 28522
rect 18321 28464 18326 28520
rect 18382 28464 21588 28520
rect 18321 28462 21588 28464
rect 18321 28459 18387 28462
rect 21582 28460 21588 28462
rect 21652 28460 21658 28524
rect 24853 28522 24919 28525
rect 26200 28522 27000 28552
rect 24853 28520 27000 28522
rect 24853 28464 24858 28520
rect 24914 28464 27000 28520
rect 24853 28462 27000 28464
rect 24853 28459 24919 28462
rect 26200 28432 27000 28462
rect 14958 28324 14964 28388
rect 15028 28386 15034 28388
rect 15285 28386 15351 28389
rect 15028 28384 15351 28386
rect 15028 28328 15290 28384
rect 15346 28328 15351 28384
rect 15028 28326 15351 28328
rect 15028 28324 15034 28326
rect 15285 28323 15351 28326
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 15837 28252 15903 28253
rect 20161 28252 20227 28253
rect 15837 28250 15884 28252
rect 15792 28248 15884 28250
rect 15792 28192 15842 28248
rect 15792 28190 15884 28192
rect 15837 28188 15884 28190
rect 15948 28188 15954 28252
rect 20110 28250 20116 28252
rect 20034 28190 20116 28250
rect 20180 28250 20227 28252
rect 21766 28250 21772 28252
rect 20180 28248 21772 28250
rect 20222 28192 21772 28248
rect 20110 28188 20116 28190
rect 20180 28190 21772 28192
rect 20180 28188 20227 28190
rect 21766 28188 21772 28190
rect 21836 28188 21842 28252
rect 15837 28187 15903 28188
rect 20161 28187 20227 28188
rect 15694 27916 15700 27980
rect 15764 27978 15770 27980
rect 16021 27978 16087 27981
rect 15764 27976 16087 27978
rect 15764 27920 16026 27976
rect 16082 27920 16087 27976
rect 15764 27918 16087 27920
rect 15764 27916 15770 27918
rect 16021 27915 16087 27918
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24117 27706 24183 27709
rect 26200 27706 27000 27736
rect 24117 27704 27000 27706
rect 24117 27648 24122 27704
rect 24178 27648 27000 27704
rect 24117 27646 27000 27648
rect 24117 27643 24183 27646
rect 26200 27616 27000 27646
rect 17166 27508 17172 27572
rect 17236 27570 17242 27572
rect 18229 27570 18295 27573
rect 18781 27570 18847 27573
rect 17236 27568 18847 27570
rect 17236 27512 18234 27568
rect 18290 27512 18786 27568
rect 18842 27512 18847 27568
rect 17236 27510 18847 27512
rect 17236 27508 17242 27510
rect 18229 27507 18295 27510
rect 18781 27507 18847 27510
rect 18597 27434 18663 27437
rect 18781 27434 18847 27437
rect 18597 27432 18847 27434
rect 18597 27376 18602 27432
rect 18658 27376 18786 27432
rect 18842 27376 18847 27432
rect 18597 27374 18847 27376
rect 18597 27371 18663 27374
rect 18781 27371 18847 27374
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25497 26890 25563 26893
rect 26200 26890 27000 26920
rect 25497 26888 27000 26890
rect 25497 26832 25502 26888
rect 25558 26832 27000 26888
rect 25497 26830 27000 26832
rect 25497 26827 25563 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 12382 26284 12388 26348
rect 12452 26346 12458 26348
rect 12525 26346 12591 26349
rect 12452 26344 12591 26346
rect 12452 26288 12530 26344
rect 12586 26288 12591 26344
rect 12452 26286 12591 26288
rect 12452 26284 12458 26286
rect 12525 26283 12591 26286
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 2773 26074 2839 26077
rect 0 26072 2839 26074
rect 0 26016 2778 26072
rect 2834 26016 2839 26072
rect 0 26014 2839 26016
rect 0 25984 800 26014
rect 2773 26011 2839 26014
rect 18597 26072 18663 26077
rect 18597 26016 18602 26072
rect 18658 26016 18663 26072
rect 18597 26011 18663 26016
rect 25313 26074 25379 26077
rect 26200 26074 27000 26104
rect 25313 26072 27000 26074
rect 25313 26016 25318 26072
rect 25374 26016 27000 26072
rect 25313 26014 27000 26016
rect 25313 26011 25379 26014
rect 18600 25805 18660 26011
rect 26200 25984 27000 26014
rect 18597 25800 18663 25805
rect 18597 25744 18602 25800
rect 18658 25744 18663 25800
rect 18597 25739 18663 25744
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 19190 24924 19196 24988
rect 19260 24986 19266 24988
rect 19517 24986 19583 24989
rect 19885 24986 19951 24989
rect 19260 24984 19951 24986
rect 19260 24928 19522 24984
rect 19578 24928 19890 24984
rect 19946 24928 19951 24984
rect 19260 24926 19951 24928
rect 19260 24924 19266 24926
rect 19517 24923 19583 24926
rect 19885 24923 19951 24926
rect 12985 24714 13051 24717
rect 13905 24714 13971 24717
rect 16849 24714 16915 24717
rect 12985 24712 16915 24714
rect 12985 24656 12990 24712
rect 13046 24656 13910 24712
rect 13966 24656 16854 24712
rect 16910 24656 16915 24712
rect 12985 24654 16915 24656
rect 12985 24651 13051 24654
rect 13905 24651 13971 24654
rect 16849 24651 16915 24654
rect 18505 24714 18571 24717
rect 25129 24714 25195 24717
rect 18505 24712 25195 24714
rect 18505 24656 18510 24712
rect 18566 24656 25134 24712
rect 25190 24656 25195 24712
rect 18505 24654 25195 24656
rect 18505 24651 18571 24654
rect 25129 24651 25195 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 24853 24442 24919 24445
rect 26200 24442 27000 24472
rect 24853 24440 27000 24442
rect 24853 24384 24858 24440
rect 24914 24384 27000 24440
rect 24853 24382 27000 24384
rect 24853 24379 24919 24382
rect 26200 24352 27000 24382
rect 9857 24306 9923 24309
rect 16389 24306 16455 24309
rect 9857 24304 16455 24306
rect 9857 24248 9862 24304
rect 9918 24248 16394 24304
rect 16450 24248 16455 24304
rect 9857 24246 16455 24248
rect 9857 24243 9923 24246
rect 16389 24243 16455 24246
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 0 23626 800 23656
rect 1301 23626 1367 23629
rect 0 23624 1367 23626
rect 0 23568 1306 23624
rect 1362 23568 1367 23624
rect 0 23566 1367 23568
rect 0 23536 800 23566
rect 1301 23563 1367 23566
rect 23841 23626 23907 23629
rect 26200 23626 27000 23656
rect 23841 23624 27000 23626
rect 23841 23568 23846 23624
rect 23902 23568 27000 23624
rect 23841 23566 27000 23568
rect 23841 23563 23907 23566
rect 26200 23536 27000 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 9806 22884 9812 22948
rect 9876 22946 9882 22948
rect 10409 22946 10475 22949
rect 10777 22946 10843 22949
rect 9876 22944 10843 22946
rect 9876 22888 10414 22944
rect 10470 22888 10782 22944
rect 10838 22888 10843 22944
rect 9876 22886 10843 22888
rect 9876 22884 9882 22886
rect 10409 22883 10475 22886
rect 10777 22883 10843 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 23289 22810 23355 22813
rect 26200 22810 27000 22840
rect 23289 22808 27000 22810
rect 23289 22752 23294 22808
rect 23350 22752 27000 22808
rect 23289 22750 27000 22752
rect 23289 22747 23355 22750
rect 26200 22720 27000 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 24853 21994 24919 21997
rect 26200 21994 27000 22024
rect 24853 21992 27000 21994
rect 24853 21936 24858 21992
rect 24914 21936 27000 21992
rect 24853 21934 27000 21936
rect 24853 21931 24919 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 14406 21660 14412 21724
rect 14476 21722 14482 21724
rect 14641 21722 14707 21725
rect 14476 21720 14707 21722
rect 14476 21664 14646 21720
rect 14702 21664 14707 21720
rect 14476 21662 14707 21664
rect 14476 21660 14482 21662
rect 14641 21659 14707 21662
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 23381 21178 23447 21181
rect 26200 21178 27000 21208
rect 23381 21176 27000 21178
rect 23381 21120 23386 21176
rect 23442 21120 27000 21176
rect 23381 21118 27000 21120
rect 23381 21115 23447 21118
rect 26200 21088 27000 21118
rect 20161 20772 20227 20773
rect 20110 20770 20116 20772
rect 20070 20710 20116 20770
rect 20180 20768 20227 20772
rect 20222 20712 20227 20768
rect 20110 20708 20116 20710
rect 20180 20708 20227 20712
rect 20161 20707 20227 20708
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 17309 20636 17375 20637
rect 17309 20634 17356 20636
rect 17264 20632 17356 20634
rect 17264 20576 17314 20632
rect 17264 20574 17356 20576
rect 17309 20572 17356 20574
rect 17420 20572 17426 20636
rect 18505 20634 18571 20637
rect 19558 20634 19564 20636
rect 18505 20632 19564 20634
rect 18505 20576 18510 20632
rect 18566 20576 19564 20632
rect 18505 20574 19564 20576
rect 17309 20571 17375 20572
rect 18505 20571 18571 20574
rect 19558 20572 19564 20574
rect 19628 20572 19634 20636
rect 24945 20362 25011 20365
rect 26200 20362 27000 20392
rect 24945 20360 27000 20362
rect 24945 20304 24950 20360
rect 25006 20304 27000 20360
rect 24945 20302 27000 20304
rect 24945 20299 25011 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 12382 19892 12388 19956
rect 12452 19954 12458 19956
rect 12893 19954 12959 19957
rect 12452 19952 12959 19954
rect 12452 19896 12898 19952
rect 12954 19896 12959 19952
rect 12452 19894 12959 19896
rect 12452 19892 12458 19894
rect 12893 19891 12959 19894
rect 17861 19954 17927 19957
rect 18638 19954 18644 19956
rect 17861 19952 18644 19954
rect 17861 19896 17866 19952
rect 17922 19896 18644 19952
rect 17861 19894 18644 19896
rect 17861 19891 17927 19894
rect 18638 19892 18644 19894
rect 18708 19892 18714 19956
rect 8661 19682 8727 19685
rect 14825 19684 14891 19685
rect 9254 19682 9260 19684
rect 8661 19680 9260 19682
rect 8661 19624 8666 19680
rect 8722 19624 9260 19680
rect 8661 19622 9260 19624
rect 8661 19619 8727 19622
rect 9254 19620 9260 19622
rect 9324 19620 9330 19684
rect 14774 19620 14780 19684
rect 14844 19682 14891 19684
rect 14844 19680 14936 19682
rect 14886 19624 14936 19680
rect 14844 19622 14936 19624
rect 14844 19620 14891 19622
rect 14825 19619 14891 19620
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 11973 19546 12039 19549
rect 12198 19546 12204 19548
rect 11973 19544 12204 19546
rect 11973 19488 11978 19544
rect 12034 19488 12204 19544
rect 11973 19486 12204 19488
rect 11973 19483 12039 19486
rect 12198 19484 12204 19486
rect 12268 19484 12274 19548
rect 24761 19546 24827 19549
rect 26200 19546 27000 19576
rect 24761 19544 27000 19546
rect 24761 19488 24766 19544
rect 24822 19488 27000 19544
rect 24761 19486 27000 19488
rect 24761 19483 24827 19486
rect 26200 19456 27000 19486
rect 12157 19410 12223 19413
rect 15285 19410 15351 19413
rect 17534 19410 17540 19412
rect 12157 19408 17540 19410
rect 12157 19352 12162 19408
rect 12218 19352 15290 19408
rect 15346 19352 17540 19408
rect 12157 19350 17540 19352
rect 12157 19347 12223 19350
rect 15285 19347 15351 19350
rect 17534 19348 17540 19350
rect 17604 19348 17610 19412
rect 18597 19410 18663 19413
rect 18822 19410 18828 19412
rect 18597 19408 18828 19410
rect 18597 19352 18602 19408
rect 18658 19352 18828 19408
rect 18597 19350 18828 19352
rect 18597 19347 18663 19350
rect 18822 19348 18828 19350
rect 18892 19348 18898 19412
rect 12750 19212 12756 19276
rect 12820 19274 12826 19276
rect 12893 19274 12959 19277
rect 12820 19272 12959 19274
rect 12820 19216 12898 19272
rect 12954 19216 12959 19272
rect 12820 19214 12959 19216
rect 12820 19212 12826 19214
rect 12893 19211 12959 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 0 18730 800 18760
rect 1301 18730 1367 18733
rect 0 18728 1367 18730
rect 0 18672 1306 18728
rect 1362 18672 1367 18728
rect 0 18670 1367 18672
rect 0 18640 800 18670
rect 1301 18667 1367 18670
rect 24669 18730 24735 18733
rect 26200 18730 27000 18760
rect 24669 18728 27000 18730
rect 24669 18672 24674 18728
rect 24730 18672 27000 18728
rect 24669 18670 27000 18672
rect 24669 18667 24735 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 12566 18124 12572 18188
rect 12636 18186 12642 18188
rect 13721 18186 13787 18189
rect 12636 18184 13787 18186
rect 12636 18128 13726 18184
rect 13782 18128 13787 18184
rect 12636 18126 13787 18128
rect 12636 18124 12642 18126
rect 13721 18123 13787 18126
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 23381 17914 23447 17917
rect 26200 17914 27000 17944
rect 23381 17912 27000 17914
rect 23381 17856 23386 17912
rect 23442 17856 27000 17912
rect 23381 17854 27000 17856
rect 23381 17851 23447 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 24761 17098 24827 17101
rect 26200 17098 27000 17128
rect 24761 17096 27000 17098
rect 24761 17040 24766 17096
rect 24822 17040 27000 17096
rect 24761 17038 27000 17040
rect 24761 17035 24827 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 15745 16828 15811 16829
rect 15694 16826 15700 16828
rect 15654 16766 15700 16826
rect 15764 16824 15811 16828
rect 15806 16768 15811 16824
rect 15694 16764 15700 16766
rect 15764 16764 15811 16768
rect 15745 16763 15811 16764
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 14733 16282 14799 16285
rect 14958 16282 14964 16284
rect 14733 16280 14964 16282
rect 14733 16224 14738 16280
rect 14794 16224 14964 16280
rect 14733 16222 14964 16224
rect 14733 16219 14799 16222
rect 14958 16220 14964 16222
rect 15028 16220 15034 16284
rect 15929 16282 15995 16285
rect 16062 16282 16068 16284
rect 15929 16280 16068 16282
rect 15929 16224 15934 16280
rect 15990 16224 16068 16280
rect 15929 16222 16068 16224
rect 15929 16219 15995 16222
rect 16062 16220 16068 16222
rect 16132 16220 16138 16284
rect 24669 16282 24735 16285
rect 26200 16282 27000 16312
rect 24669 16280 27000 16282
rect 24669 16224 24674 16280
rect 24730 16224 27000 16280
rect 24669 16222 27000 16224
rect 24669 16219 24735 16222
rect 26200 16192 27000 16222
rect 8937 16146 9003 16149
rect 10174 16146 10180 16148
rect 8937 16144 10180 16146
rect 8937 16088 8942 16144
rect 8998 16088 10180 16144
rect 8937 16086 10180 16088
rect 8937 16083 9003 16086
rect 10174 16084 10180 16086
rect 10244 16084 10250 16148
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 26049 15466 26115 15469
rect 26200 15466 27000 15496
rect 26049 15464 27000 15466
rect 26049 15408 26054 15464
rect 26110 15408 27000 15464
rect 26049 15406 27000 15408
rect 26049 15403 26115 15406
rect 26200 15376 27000 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 25129 14650 25195 14653
rect 26200 14650 27000 14680
rect 25129 14648 27000 14650
rect 25129 14592 25134 14648
rect 25190 14592 27000 14648
rect 25129 14590 27000 14592
rect 25129 14587 25195 14590
rect 26200 14560 27000 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 12801 13972 12867 13973
rect 12750 13908 12756 13972
rect 12820 13970 12867 13972
rect 12820 13968 12912 13970
rect 12862 13912 12912 13968
rect 12820 13910 12912 13912
rect 12820 13908 12867 13910
rect 12801 13907 12867 13908
rect 0 13834 800 13864
rect 1301 13834 1367 13837
rect 0 13832 1367 13834
rect 0 13776 1306 13832
rect 1362 13776 1367 13832
rect 0 13774 1367 13776
rect 0 13744 800 13774
rect 1301 13771 1367 13774
rect 24761 13834 24827 13837
rect 26200 13834 27000 13864
rect 24761 13832 27000 13834
rect 24761 13776 24766 13832
rect 24822 13776 27000 13832
rect 24761 13774 27000 13776
rect 24761 13771 24827 13774
rect 26200 13744 27000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 19425 13426 19491 13429
rect 21265 13426 21331 13429
rect 19425 13424 21331 13426
rect 19425 13368 19430 13424
rect 19486 13368 21270 13424
rect 21326 13368 21331 13424
rect 19425 13366 21331 13368
rect 19425 13363 19491 13366
rect 21265 13363 21331 13366
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 16021 13018 16087 13021
rect 25129 13018 25195 13021
rect 26200 13018 27000 13048
rect 16021 13016 16130 13018
rect 16021 12960 16026 13016
rect 16082 12960 16130 13016
rect 16021 12955 16130 12960
rect 25129 13016 27000 13018
rect 25129 12960 25134 13016
rect 25190 12960 27000 13016
rect 25129 12958 27000 12960
rect 25129 12955 25195 12958
rect 16070 12610 16130 12955
rect 26200 12928 27000 12958
rect 16205 12610 16271 12613
rect 16070 12608 16271 12610
rect 16070 12552 16210 12608
rect 16266 12552 16271 12608
rect 16070 12550 16271 12552
rect 16205 12547 16271 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 24761 12202 24827 12205
rect 26200 12202 27000 12232
rect 24761 12200 27000 12202
rect 24761 12144 24766 12200
rect 24822 12144 27000 12200
rect 24761 12142 27000 12144
rect 24761 12139 24827 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 17493 11932 17559 11933
rect 17493 11930 17540 11932
rect 17448 11928 17540 11930
rect 17448 11872 17498 11928
rect 17448 11870 17540 11872
rect 17493 11868 17540 11870
rect 17604 11868 17610 11932
rect 17493 11867 17559 11868
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24669 11386 24735 11389
rect 26200 11386 27000 11416
rect 0 11326 1778 11386
rect 0 11296 800 11326
rect 1718 11250 1778 11326
rect 24669 11384 27000 11386
rect 24669 11328 24674 11384
rect 24730 11328 27000 11384
rect 24669 11326 27000 11328
rect 24669 11323 24735 11326
rect 26200 11296 27000 11326
rect 3509 11250 3575 11253
rect 1718 11248 3575 11250
rect 1718 11192 3514 11248
rect 3570 11192 3575 11248
rect 1718 11190 3575 11192
rect 3509 11187 3575 11190
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 24577 10570 24643 10573
rect 26200 10570 27000 10600
rect 24577 10568 27000 10570
rect 24577 10512 24582 10568
rect 24638 10512 27000 10568
rect 24577 10510 27000 10512
rect 24577 10507 24643 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 24945 9754 25011 9757
rect 26200 9754 27000 9784
rect 24945 9752 27000 9754
rect 24945 9696 24950 9752
rect 25006 9696 27000 9752
rect 24945 9694 27000 9696
rect 24945 9691 25011 9694
rect 26200 9664 27000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 0 8938 800 8968
rect 4061 8938 4127 8941
rect 0 8936 4127 8938
rect 0 8880 4066 8936
rect 4122 8880 4127 8936
rect 0 8878 4127 8880
rect 0 8848 800 8878
rect 4061 8875 4127 8878
rect 24669 8938 24735 8941
rect 26200 8938 27000 8968
rect 24669 8936 27000 8938
rect 24669 8880 24674 8936
rect 24730 8880 27000 8936
rect 24669 8878 27000 8880
rect 24669 8875 24735 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 1945 8394 2011 8397
rect 9254 8394 9260 8396
rect 1945 8392 9260 8394
rect 1945 8336 1950 8392
rect 2006 8336 9260 8392
rect 1945 8334 9260 8336
rect 1945 8331 2011 8334
rect 9254 8332 9260 8334
rect 9324 8332 9330 8396
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24577 8122 24643 8125
rect 26200 8122 27000 8152
rect 24577 8120 27000 8122
rect 24577 8064 24582 8120
rect 24638 8064 27000 8120
rect 24577 8062 27000 8064
rect 24577 8059 24643 8062
rect 26200 8032 27000 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 24761 7306 24827 7309
rect 26200 7306 27000 7336
rect 24761 7304 27000 7306
rect 24761 7248 24766 7304
rect 24822 7248 27000 7304
rect 24761 7246 27000 7248
rect 24761 7243 24827 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 4061 6490 4127 6493
rect 0 6488 4127 6490
rect 0 6432 4066 6488
rect 4122 6432 4127 6488
rect 0 6430 4127 6432
rect 0 6400 800 6430
rect 4061 6427 4127 6430
rect 24945 6490 25011 6493
rect 26200 6490 27000 6520
rect 24945 6488 27000 6490
rect 24945 6432 24950 6488
rect 25006 6432 27000 6488
rect 24945 6430 27000 6432
rect 24945 6427 25011 6430
rect 26200 6400 27000 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 9581 5674 9647 5677
rect 14774 5674 14780 5676
rect 9581 5672 14780 5674
rect 9581 5616 9586 5672
rect 9642 5616 14780 5672
rect 9581 5614 14780 5616
rect 9581 5611 9647 5614
rect 14774 5612 14780 5614
rect 14844 5612 14850 5676
rect 25129 5674 25195 5677
rect 26200 5674 27000 5704
rect 25129 5672 27000 5674
rect 25129 5616 25134 5672
rect 25190 5616 27000 5672
rect 25129 5614 27000 5616
rect 25129 5611 25195 5614
rect 26200 5584 27000 5614
rect 9857 5538 9923 5541
rect 12198 5538 12204 5540
rect 9857 5536 12204 5538
rect 9857 5480 9862 5536
rect 9918 5480 12204 5536
rect 9857 5478 12204 5480
rect 9857 5475 9923 5478
rect 12198 5476 12204 5478
rect 12268 5476 12274 5540
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23381 4858 23447 4861
rect 26200 4858 27000 4888
rect 23381 4856 27000 4858
rect 23381 4800 23386 4856
rect 23442 4800 27000 4856
rect 23381 4798 27000 4800
rect 23381 4795 23447 4798
rect 26200 4768 27000 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 8201 4178 8267 4181
rect 9806 4178 9812 4180
rect 8201 4176 9812 4178
rect 8201 4120 8206 4176
rect 8262 4120 9812 4176
rect 8201 4118 9812 4120
rect 8201 4115 8267 4118
rect 9806 4116 9812 4118
rect 9876 4116 9882 4180
rect 0 4042 800 4072
rect 4061 4042 4127 4045
rect 18781 4044 18847 4045
rect 18781 4042 18828 4044
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 18736 4040 18828 4042
rect 18736 3984 18786 4040
rect 18736 3982 18828 3984
rect 0 3952 800 3982
rect 4061 3979 4127 3982
rect 18781 3980 18828 3982
rect 18892 3980 18898 4044
rect 22093 4042 22159 4045
rect 26200 4042 27000 4072
rect 22093 4040 27000 4042
rect 22093 3984 22098 4040
rect 22154 3984 27000 4040
rect 22093 3982 27000 3984
rect 18781 3979 18847 3980
rect 22093 3979 22159 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 22553 3226 22619 3229
rect 26200 3226 27000 3256
rect 22553 3224 27000 3226
rect 22553 3168 22558 3224
rect 22614 3168 27000 3224
rect 22553 3166 27000 3168
rect 22553 3163 22619 3166
rect 26200 3136 27000 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 21633 2410 21699 2413
rect 26200 2410 27000 2440
rect 21633 2408 27000 2410
rect 21633 2352 21638 2408
rect 21694 2352 27000 2408
rect 21633 2350 27000 2352
rect 21633 2347 21699 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 24853 1594 24919 1597
rect 26200 1594 27000 1624
rect 24853 1592 27000 1594
rect 24853 1536 24858 1592
rect 24914 1536 27000 1592
rect 24853 1534 27000 1536
rect 24853 1531 24919 1534
rect 26200 1504 27000 1534
rect 24945 778 25011 781
rect 26200 778 27000 808
rect 24945 776 27000 778
rect 24945 720 24950 776
rect 25006 720 27000 776
rect 24945 718 27000 720
rect 24945 715 25011 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 17172 53892 17236 53956
rect 21956 53892 22020 53956
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 14044 52592 14108 52596
rect 14044 52536 14058 52592
rect 14058 52536 14108 52592
rect 14044 52532 14108 52536
rect 14596 52532 14660 52596
rect 16436 52592 16500 52596
rect 16436 52536 16450 52592
rect 16450 52536 16500 52592
rect 16436 52532 16500 52536
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 22324 51036 22388 51100
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 20300 46956 20364 47020
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 21772 46276 21836 46340
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 20116 45792 20180 45796
rect 20116 45736 20130 45792
rect 20130 45736 20180 45792
rect 20116 45732 20180 45736
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 9812 44704 9876 44708
rect 9812 44648 9826 44704
rect 9826 44648 9876 44704
rect 9812 44644 9876 44648
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 12204 44236 12268 44300
rect 23428 44236 23492 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 21588 43344 21652 43348
rect 21588 43288 21638 43344
rect 21638 43288 21652 43344
rect 21588 43284 21652 43288
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 10916 42468 10980 42532
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 22692 42332 22756 42396
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 22692 41652 22756 41716
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 22324 40700 22388 40764
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 15884 40080 15948 40084
rect 15884 40024 15934 40080
rect 15934 40024 15948 40080
rect 15884 40020 15948 40024
rect 20668 40020 20732 40084
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 18644 38796 18708 38860
rect 17356 38660 17420 38724
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 22692 37844 22756 37908
rect 12204 37708 12268 37772
rect 20484 37708 20548 37772
rect 23428 37708 23492 37772
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 9812 36756 9876 36820
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 12756 36076 12820 36140
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 20668 34308 20732 34372
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 12204 33356 12268 33420
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 20300 33084 20364 33148
rect 22692 32676 22756 32740
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 14412 32600 14476 32604
rect 14412 32544 14426 32600
rect 14426 32544 14476 32600
rect 14412 32540 14476 32544
rect 21956 32540 22020 32604
rect 12204 32328 12268 32332
rect 12204 32272 12254 32328
rect 12254 32272 12268 32328
rect 12204 32268 12268 32272
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 19564 31860 19628 31924
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 20116 31512 20180 31516
rect 20116 31456 20130 31512
rect 20130 31456 20180 31512
rect 20116 31452 20180 31456
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 20484 30968 20548 30972
rect 20484 30912 20498 30968
rect 20498 30912 20548 30968
rect 20484 30908 20548 30912
rect 10180 30636 10244 30700
rect 14044 30636 14108 30700
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 14596 30228 14660 30292
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 16436 29744 16500 29748
rect 16436 29688 16450 29744
rect 16450 29688 16500 29744
rect 16436 29684 16500 29688
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 16068 29004 16132 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 19196 28596 19260 28660
rect 21588 28460 21652 28524
rect 14964 28324 15028 28388
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 15884 28248 15948 28252
rect 15884 28192 15898 28248
rect 15898 28192 15948 28248
rect 15884 28188 15948 28192
rect 20116 28248 20180 28252
rect 20116 28192 20166 28248
rect 20166 28192 20180 28248
rect 20116 28188 20180 28192
rect 21772 28188 21836 28252
rect 15700 27916 15764 27980
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 17172 27508 17236 27572
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 12388 26284 12452 26348
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 19196 24924 19260 24988
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 9812 22884 9876 22948
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 14412 21660 14476 21724
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 20116 20768 20180 20772
rect 20116 20712 20166 20768
rect 20166 20712 20180 20768
rect 20116 20708 20180 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 17356 20632 17420 20636
rect 17356 20576 17370 20632
rect 17370 20576 17420 20632
rect 17356 20572 17420 20576
rect 19564 20572 19628 20636
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 12388 19892 12452 19956
rect 18644 19892 18708 19956
rect 9260 19620 9324 19684
rect 14780 19680 14844 19684
rect 14780 19624 14830 19680
rect 14830 19624 14844 19680
rect 14780 19620 14844 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 12204 19484 12268 19548
rect 17540 19348 17604 19412
rect 18828 19348 18892 19412
rect 12756 19212 12820 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 12572 18124 12636 18188
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 15700 16824 15764 16828
rect 15700 16768 15750 16824
rect 15750 16768 15764 16824
rect 15700 16764 15764 16768
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 14964 16220 15028 16284
rect 16068 16220 16132 16284
rect 10180 16084 10244 16148
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 12756 13968 12820 13972
rect 12756 13912 12806 13968
rect 12806 13912 12820 13968
rect 12756 13908 12820 13912
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 17540 11928 17604 11932
rect 17540 11872 17554 11928
rect 17554 11872 17604 11928
rect 17540 11868 17604 11872
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 9260 8332 9324 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 14780 5612 14844 5676
rect 12204 5476 12268 5540
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 9812 4116 9876 4180
rect 18828 4040 18892 4044
rect 18828 3984 18842 4040
rect 18842 3984 18892 4040
rect 18828 3980 18892 3984
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 12944 53888 13264 54448
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17171 53956 17237 53957
rect 17171 53892 17172 53956
rect 17236 53892 17237 53956
rect 17171 53891 17237 53892
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 14043 52596 14109 52597
rect 14043 52532 14044 52596
rect 14108 52532 14109 52596
rect 14043 52531 14109 52532
rect 14595 52596 14661 52597
rect 14595 52532 14596 52596
rect 14660 52532 14661 52596
rect 14595 52531 14661 52532
rect 16435 52596 16501 52597
rect 16435 52532 16436 52596
rect 16500 52532 16501 52596
rect 16435 52531 16501 52532
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 9811 44708 9877 44709
rect 9811 44644 9812 44708
rect 9876 44644 9877 44708
rect 9811 44643 9877 44644
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 9814 36821 9874 44643
rect 12203 44300 12269 44301
rect 12203 44236 12204 44300
rect 12268 44236 12269 44300
rect 12203 44235 12269 44236
rect 10915 42532 10981 42533
rect 10915 42468 10916 42532
rect 10980 42468 10981 42532
rect 10915 42467 10981 42468
rect 9811 36820 9877 36821
rect 9811 36756 9812 36820
rect 9876 36756 9877 36820
rect 9811 36755 9877 36756
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 10918 31770 10978 42467
rect 12206 37773 12266 44235
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12203 37772 12269 37773
rect 12203 37708 12204 37772
rect 12268 37708 12269 37772
rect 12203 37707 12269 37708
rect 12206 33421 12266 37707
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12755 36140 12821 36141
rect 12755 36076 12756 36140
rect 12820 36076 12821 36140
rect 12755 36075 12821 36076
rect 12203 33420 12269 33421
rect 12203 33356 12204 33420
rect 12268 33356 12269 33420
rect 12203 33355 12269 33356
rect 12203 32332 12269 32333
rect 12203 32268 12204 32332
rect 12268 32268 12269 32332
rect 12203 32267 12269 32268
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 10182 31710 10978 31770
rect 10182 30701 10242 31710
rect 10179 30700 10245 30701
rect 10179 30636 10180 30700
rect 10244 30636 10245 30700
rect 10179 30635 10245 30636
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 9811 22948 9877 22949
rect 9811 22884 9812 22948
rect 9876 22884 9877 22948
rect 9811 22883 9877 22884
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 9259 19684 9325 19685
rect 9259 19620 9260 19684
rect 9324 19620 9325 19684
rect 9259 19619 9325 19620
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 9262 8397 9322 19619
rect 9259 8396 9325 8397
rect 9259 8332 9260 8396
rect 9324 8332 9325 8396
rect 9259 8331 9325 8332
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 9814 4181 9874 22883
rect 10182 16149 10242 30635
rect 12206 19549 12266 32267
rect 12387 26348 12453 26349
rect 12387 26284 12388 26348
rect 12452 26284 12453 26348
rect 12387 26283 12453 26284
rect 12390 19957 12450 26283
rect 12758 22110 12818 36075
rect 12574 22050 12818 22110
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 14046 30701 14106 52531
rect 14411 32604 14477 32605
rect 14411 32540 14412 32604
rect 14476 32540 14477 32604
rect 14411 32539 14477 32540
rect 14043 30700 14109 30701
rect 14043 30636 14044 30700
rect 14108 30636 14109 30700
rect 14043 30635 14109 30636
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12387 19956 12453 19957
rect 12387 19892 12388 19956
rect 12452 19892 12453 19956
rect 12387 19891 12453 19892
rect 12203 19548 12269 19549
rect 12203 19484 12204 19548
rect 12268 19484 12269 19548
rect 12203 19483 12269 19484
rect 12574 18189 12634 22050
rect 12944 21248 13264 22272
rect 14414 21725 14474 32539
rect 14598 30293 14658 52531
rect 15883 40084 15949 40085
rect 15883 40020 15884 40084
rect 15948 40020 15949 40084
rect 15883 40019 15949 40020
rect 14595 30292 14661 30293
rect 14595 30228 14596 30292
rect 14660 30228 14661 30292
rect 14595 30227 14661 30228
rect 14963 28388 15029 28389
rect 14963 28324 14964 28388
rect 15028 28324 15029 28388
rect 14963 28323 15029 28324
rect 14411 21724 14477 21725
rect 14411 21660 14412 21724
rect 14476 21660 14477 21724
rect 14411 21659 14477 21660
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12755 19276 12821 19277
rect 12755 19212 12756 19276
rect 12820 19212 12821 19276
rect 12755 19211 12821 19212
rect 12571 18188 12637 18189
rect 12571 18124 12572 18188
rect 12636 18124 12637 18188
rect 12571 18123 12637 18124
rect 10179 16148 10245 16149
rect 10179 16084 10180 16148
rect 10244 16084 10245 16148
rect 10179 16083 10245 16084
rect 12574 12450 12634 18123
rect 12758 13973 12818 19211
rect 12944 19072 13264 20096
rect 14779 19684 14845 19685
rect 14779 19620 14780 19684
rect 14844 19620 14845 19684
rect 14779 19619 14845 19620
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12755 13972 12821 13973
rect 12755 13908 12756 13972
rect 12820 13908 12821 13972
rect 12755 13907 12821 13908
rect 12206 12390 12634 12450
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12206 5541 12266 12390
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12203 5540 12269 5541
rect 12203 5476 12204 5540
rect 12268 5476 12269 5540
rect 12203 5475 12269 5476
rect 12944 4928 13264 5952
rect 14782 5677 14842 19619
rect 14966 16285 15026 28323
rect 15886 28253 15946 40019
rect 16438 29749 16498 52531
rect 16435 29748 16501 29749
rect 16435 29684 16436 29748
rect 16500 29684 16501 29748
rect 16435 29683 16501 29684
rect 16067 29068 16133 29069
rect 16067 29004 16068 29068
rect 16132 29004 16133 29068
rect 16067 29003 16133 29004
rect 15883 28252 15949 28253
rect 15883 28188 15884 28252
rect 15948 28188 15949 28252
rect 15883 28187 15949 28188
rect 15699 27980 15765 27981
rect 15699 27916 15700 27980
rect 15764 27916 15765 27980
rect 15699 27915 15765 27916
rect 15702 16829 15762 27915
rect 15699 16828 15765 16829
rect 15699 16764 15700 16828
rect 15764 16764 15765 16828
rect 15699 16763 15765 16764
rect 16070 16285 16130 29003
rect 17174 27573 17234 53891
rect 17944 53344 18264 54368
rect 21955 53956 22021 53957
rect 21955 53892 21956 53956
rect 22020 53892 22021 53956
rect 21955 53891 22021 53892
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 20299 47020 20365 47021
rect 20299 46956 20300 47020
rect 20364 46956 20365 47020
rect 20299 46955 20365 46956
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 20115 45796 20181 45797
rect 20115 45732 20116 45796
rect 20180 45732 20181 45796
rect 20115 45731 20181 45732
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17355 38724 17421 38725
rect 17355 38660 17356 38724
rect 17420 38660 17421 38724
rect 17355 38659 17421 38660
rect 17171 27572 17237 27573
rect 17171 27508 17172 27572
rect 17236 27508 17237 27572
rect 17171 27507 17237 27508
rect 17358 20637 17418 38659
rect 17944 38112 18264 39136
rect 18643 38860 18709 38861
rect 18643 38796 18644 38860
rect 18708 38796 18709 38860
rect 18643 38795 18709 38796
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17355 20636 17421 20637
rect 17355 20572 17356 20636
rect 17420 20572 17421 20636
rect 17355 20571 17421 20572
rect 17944 19616 18264 20640
rect 18646 19957 18706 38795
rect 19563 31924 19629 31925
rect 19563 31860 19564 31924
rect 19628 31860 19629 31924
rect 19563 31859 19629 31860
rect 19195 28660 19261 28661
rect 19195 28596 19196 28660
rect 19260 28596 19261 28660
rect 19195 28595 19261 28596
rect 19198 24989 19258 28595
rect 19195 24988 19261 24989
rect 19195 24924 19196 24988
rect 19260 24924 19261 24988
rect 19195 24923 19261 24924
rect 19566 20637 19626 31859
rect 20118 31517 20178 45731
rect 20302 33149 20362 46955
rect 21771 46340 21837 46341
rect 21771 46276 21772 46340
rect 21836 46276 21837 46340
rect 21771 46275 21837 46276
rect 21587 43348 21653 43349
rect 21587 43284 21588 43348
rect 21652 43284 21653 43348
rect 21587 43283 21653 43284
rect 20667 40084 20733 40085
rect 20667 40020 20668 40084
rect 20732 40020 20733 40084
rect 20667 40019 20733 40020
rect 20483 37772 20549 37773
rect 20483 37708 20484 37772
rect 20548 37708 20549 37772
rect 20483 37707 20549 37708
rect 20299 33148 20365 33149
rect 20299 33084 20300 33148
rect 20364 33084 20365 33148
rect 20299 33083 20365 33084
rect 20115 31516 20181 31517
rect 20115 31452 20116 31516
rect 20180 31452 20181 31516
rect 20115 31451 20181 31452
rect 20486 30973 20546 37707
rect 20670 34373 20730 40019
rect 20667 34372 20733 34373
rect 20667 34308 20668 34372
rect 20732 34308 20733 34372
rect 20667 34307 20733 34308
rect 20483 30972 20549 30973
rect 20483 30908 20484 30972
rect 20548 30908 20549 30972
rect 20483 30907 20549 30908
rect 21590 28525 21650 43283
rect 21587 28524 21653 28525
rect 21587 28460 21588 28524
rect 21652 28460 21653 28524
rect 21587 28459 21653 28460
rect 21774 28253 21834 46275
rect 21958 32605 22018 53891
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22323 51100 22389 51101
rect 22323 51036 22324 51100
rect 22388 51036 22389 51100
rect 22323 51035 22389 51036
rect 22326 40765 22386 51035
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 23427 44300 23493 44301
rect 23427 44236 23428 44300
rect 23492 44236 23493 44300
rect 23427 44235 23493 44236
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22691 42396 22757 42397
rect 22691 42332 22692 42396
rect 22756 42332 22757 42396
rect 22691 42331 22757 42332
rect 22694 41717 22754 42331
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22691 41716 22757 41717
rect 22691 41652 22692 41716
rect 22756 41652 22757 41716
rect 22691 41651 22757 41652
rect 22323 40764 22389 40765
rect 22323 40700 22324 40764
rect 22388 40700 22389 40764
rect 22323 40699 22389 40700
rect 22694 37909 22754 41651
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22691 37908 22757 37909
rect 22691 37844 22692 37908
rect 22756 37844 22757 37908
rect 22691 37843 22757 37844
rect 22694 32741 22754 37843
rect 22944 37568 23264 38592
rect 23430 37773 23490 44235
rect 23427 37772 23493 37773
rect 23427 37708 23428 37772
rect 23492 37708 23493 37772
rect 23427 37707 23493 37708
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22691 32740 22757 32741
rect 22691 32676 22692 32740
rect 22756 32676 22757 32740
rect 22691 32675 22757 32676
rect 21955 32604 22021 32605
rect 21955 32540 21956 32604
rect 22020 32540 22021 32604
rect 21955 32539 22021 32540
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 20115 28252 20181 28253
rect 20115 28188 20116 28252
rect 20180 28188 20181 28252
rect 20115 28187 20181 28188
rect 21771 28252 21837 28253
rect 21771 28188 21772 28252
rect 21836 28188 21837 28252
rect 21771 28187 21837 28188
rect 20118 20773 20178 28187
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 20115 20772 20181 20773
rect 20115 20708 20116 20772
rect 20180 20708 20181 20772
rect 20115 20707 20181 20708
rect 19563 20636 19629 20637
rect 19563 20572 19564 20636
rect 19628 20572 19629 20636
rect 19563 20571 19629 20572
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 18643 19956 18709 19957
rect 18643 19892 18644 19956
rect 18708 19892 18709 19956
rect 18643 19891 18709 19892
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 14963 16284 15029 16285
rect 14963 16220 14964 16284
rect 15028 16220 15029 16284
rect 14963 16219 15029 16220
rect 16067 16284 16133 16285
rect 16067 16220 16068 16284
rect 16132 16220 16133 16284
rect 16067 16219 16133 16220
rect 17542 11933 17602 19347
rect 17944 18528 18264 19552
rect 18827 19412 18893 19413
rect 18827 19348 18828 19412
rect 18892 19348 18893 19412
rect 18827 19347 18893 19348
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17539 11932 17605 11933
rect 17539 11868 17540 11932
rect 17604 11868 17605 11932
rect 17539 11867 17605 11868
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 14779 5676 14845 5677
rect 14779 5612 14780 5676
rect 14844 5612 14845 5676
rect 14779 5611 14845 5612
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 9811 4180 9877 4181
rect 9811 4116 9812 4180
rect 9876 4116 9877 4180
rect 9811 4115 9877 4116
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 18830 4045 18890 19347
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 18827 4044 18893 4045
rect 18827 3980 18828 4044
rect 18892 3980 18893 4044
rect 18827 3979 18893 3980
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1676037725
transform 1 0 23736 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1676037725
transform 1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 23184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 24656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 23736 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 24564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 25024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 22172 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 14076 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 13616 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 17112 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 20608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 19044 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 21068 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 3128 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 6716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform 1 0 4692 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 4968 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 6532 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 6808 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 6624 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 6532 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 7268 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 7636 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 7912 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform 1 0 6808 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 10396 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1676037725
transform 1 0 9200 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 11408 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 10856 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 11408 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 9016 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 9292 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1676037725
transform 1 0 10212 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 11684 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 12604 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 12328 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1676037725
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _203_
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12696 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform -1 0 11408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 11960 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1676037725
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 18952 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1676037725
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1676037725
transform 1 0 19596 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1676037725
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1676037725
transform 1 0 3680 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1676037725
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1676037725
transform 1 0 3772 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1676037725
transform 1 0 5244 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1676037725
transform 1 0 5520 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1676037725
transform 1 0 7084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1676037725
transform 1 0 7176 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1676037725
transform 1 0 6348 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1676037725
transform 1 0 8464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1676037725
transform 1 0 9384 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1676037725
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1676037725
transform 1 0 10212 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1676037725
transform 1 0 11960 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1676037725
transform 1 0 11040 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1676037725
transform 1 0 12052 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 9384 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__CLK
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 12144 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16008 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15088 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13156 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10028 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13616 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 7452 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 10396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 3956 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 2576 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6624 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 4324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 10304 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 10672 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21068 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 18492 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 24104 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold10_A
timestamp 1676037725
transform 1 0 3956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold12_A
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 25208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 24472 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 24748 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 25208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 24748 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 24748 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 24748 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 24748 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 9016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 17204 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 18860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 18676 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 19688 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 19320 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 19504 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 20700 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 13156 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 20792 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 21160 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 20976 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 23276 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 22264 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform 1 0 22540 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform 1 0 24380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform 1 0 14812 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform 1 0 14444 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform 1 0 16100 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform 1 0 16100 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform 1 0 2024 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform 1 0 2024 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform 1 0 2024 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform 1 0 2024 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform 1 0 2116 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform 1 0 24656 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform 1 0 25208 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform 1 0 2116 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform 1 0 5060 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1676037725
transform 1 0 3220 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1676037725
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 16100 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21896 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17572 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17940 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18216 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 15824 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17112 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21712 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20792 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 24748 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24656 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 23736 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20424 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17664 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 17112 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11776 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9752 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 6532 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 8832 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 9844 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 15180 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14168 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14260 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 13156 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12972 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 10580 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 8648 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10488 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7268 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 7728 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 7544 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 9016 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10856 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8096 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 6900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1676037725
transform 1 0 8004 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__CLK
timestamp 1676037725
transform 1 0 8096 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 7912 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 9292 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12788 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18032 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17020 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 19228 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19044 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 17848 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 11592 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 12972 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18860 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20056 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20424 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18124 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18124 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 17940 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20240 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 18216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 13064 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21528 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 17204 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20516 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20700 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23276 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19688 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15732 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17296 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20976 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18768 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20424 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16008 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_bottom_track_53.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 10856 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 23276 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22816 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22632 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21896 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 23276 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22448 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 22264 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 22264 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 21252 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21620 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 23184 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 20608 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21252 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21620 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 22080 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21896 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18584 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 20608 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20700 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 20976 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 20792 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 15732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19320 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 20240 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 19044 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19044 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17664 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 12328 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15640 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 14168 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13616 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 10028 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16100 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11040 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16100 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15088 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12236 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 7268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 23276 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 8556 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9108 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18308 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18124 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 13984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 15548 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 8832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 9016 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 17848 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18400 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 12328 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14812 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 14628 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 10580 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 10764 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 12144 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 8464 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 10212 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18216 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 13616 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 8464 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 8096 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 8280 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 8464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 17848 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 12420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 8280 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11776 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 7268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 7452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15732 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 14352 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 8924 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 9108 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13156 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 12512 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 4600 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 12236 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11040 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1676037725
transform 1 0 12880 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 7452 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4048 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5704 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 8004 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6624 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 5336 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5796 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__256 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 8280 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7084 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14260 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11408 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10120 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__257
timestamp 1676037725
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10488 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14444 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12328 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__258
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8924 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 6256 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13524 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__259
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 6808 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3680 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 4232 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 2944 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 4232 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 4508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 3680 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9844 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8464 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 10488 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17480 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 20516 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 9108 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 10212 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 9292 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 11960 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1676037725
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1676037725
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1676037725
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_37
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_59
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_66
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1676037725
transform 1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1676037725
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1676037725
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1676037725
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1676037725
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_207 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_252
timestamp 1676037725
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_260
timestamp 1676037725
transform 1 0 25024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_31
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1676037725
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_63
timestamp 1676037725
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_73
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_79
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1676037725
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1676037725
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1676037725
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1676037725
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1676037725
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1676037725
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_235 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_241
timestamp 1676037725
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1676037725
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_59
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_71
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1676037725
transform 1 0 8740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_95
timestamp 1676037725
transform 1 0 9844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1676037725
transform 1 0 14996 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1676037725
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1676037725
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1676037725
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_235
timestamp 1676037725
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_8
timestamp 1676037725
transform 1 0 1840 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 1676037725
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_32
timestamp 1676037725
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_44
timestamp 1676037725
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1676037725
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_195
timestamp 1676037725
transform 1 0 19044 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1676037725
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_29
timestamp 1676037725
transform 1 0 3772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_41
timestamp 1676037725
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1676037725
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1676037725
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1676037725
transform 1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1676037725
transform 1 0 20148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1676037725
transform 1 0 19044 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_203
timestamp 1676037725
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1676037725
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_61
timestamp 1676037725
transform 1 0 6716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_73
timestamp 1676037725
transform 1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1676037725
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_205
timestamp 1676037725
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_211
timestamp 1676037725
transform 1 0 20516 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_220
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_263
timestamp 1676037725
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_203
timestamp 1676037725
transform 1 0 19780 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1676037725
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_225
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_237
timestamp 1676037725
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1676037725
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1676037725
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1676037725
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_80
timestamp 1676037725
transform 1 0 8464 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1676037725
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1676037725
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_175
timestamp 1676037725
transform 1 0 17204 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_198
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_210
timestamp 1676037725
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1676037725
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_238
timestamp 1676037725
transform 1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_246
timestamp 1676037725
transform 1 0 23736 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1676037725
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_150
timestamp 1676037725
transform 1 0 14904 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_162
timestamp 1676037725
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_168
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1676037725
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1676037725
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1676037725
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_222
timestamp 1676037725
transform 1 0 21528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_226
timestamp 1676037725
transform 1 0 21896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1676037725
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_259
timestamp 1676037725
transform 1 0 24932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1676037725
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_126
timestamp 1676037725
transform 1 0 12696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_138
timestamp 1676037725
transform 1 0 13800 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1676037725
transform 1 0 14536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1676037725
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_156
timestamp 1676037725
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1676037725
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1676037725
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_212
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_243
timestamp 1676037725
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_151
timestamp 1676037725
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_212
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1676037725
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1676037725
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1676037725
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1676037725
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_257
timestamp 1676037725
transform 1 0 24748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_265
timestamp 1676037725
transform 1 0 25484 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1676037725
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_199
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1676037725
transform 1 0 23000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1676037725
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_115
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_127
timestamp 1676037725
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_131
timestamp 1676037725
transform 1 0 13156 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_134
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1676037725
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1676037725
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1676037725
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1676037725
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_196
timestamp 1676037725
transform 1 0 19136 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1676037725
transform 1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1676037725
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1676037725
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1676037725
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_89
timestamp 1676037725
transform 1 0 9292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1676037725
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1676037725
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1676037725
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1676037725
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_170
timestamp 1676037725
transform 1 0 16744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1676037725
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1676037725
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_212
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_215
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1676037725
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_142
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_154
timestamp 1676037725
transform 1 0 15272 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1676037725
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_227
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_241
timestamp 1676037725
transform 1 0 23276 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1676037725
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_120
timestamp 1676037725
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1676037725
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_147
timestamp 1676037725
transform 1 0 14628 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_179
timestamp 1676037725
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1676037725
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_202
timestamp 1676037725
transform 1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_207
timestamp 1676037725
transform 1 0 20148 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_235
timestamp 1676037725
transform 1 0 22724 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1676037725
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_115
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1676037725
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1676037725
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1676037725
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1676037725
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1676037725
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1676037725
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1676037725
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_182
timestamp 1676037725
transform 1 0 17848 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1676037725
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1676037725
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_208
timestamp 1676037725
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_233
timestamp 1676037725
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_245
timestamp 1676037725
transform 1 0 23644 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_100
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1676037725
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_129
timestamp 1676037725
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_164
timestamp 1676037725
transform 1 0 16192 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_174
timestamp 1676037725
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1676037725
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1676037725
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1676037725
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1676037725
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_228
timestamp 1676037725
transform 1 0 22080 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_18
timestamp 1676037725
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1676037725
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1676037725
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1676037725
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1676037725
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_124
timestamp 1676037725
transform 1 0 12512 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_128
timestamp 1676037725
transform 1 0 12880 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_131
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1676037725
transform 1 0 14444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_157
timestamp 1676037725
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1676037725
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1676037725
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1676037725
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_206
timestamp 1676037725
transform 1 0 20056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_243
timestamp 1676037725
transform 1 0 23460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1676037725
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_72
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_100
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_111
timestamp 1676037725
transform 1 0 11316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1676037725
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1676037725
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1676037725
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1676037725
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_179
timestamp 1676037725
transform 1 0 17572 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_199
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 1676037725
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1676037725
transform 1 0 20884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_244
timestamp 1676037725
transform 1 0 23552 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1676037725
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_82
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1676037725
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp 1676037725
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp 1676037725
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_115
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_154
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1676037725
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_174
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1676037725
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_204
timestamp 1676037725
transform 1 0 19872 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_217
timestamp 1676037725
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_221
timestamp 1676037725
transform 1 0 21436 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1676037725
transform 1 0 23828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_78
timestamp 1676037725
transform 1 0 8280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_96
timestamp 1676037725
transform 1 0 9936 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1676037725
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1676037725
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1676037725
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1676037725
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_248
timestamp 1676037725
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_259
timestamp 1676037725
transform 1 0 24932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1676037725
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp 1676037725
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1676037725
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_95
timestamp 1676037725
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1676037725
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1676037725
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_132
timestamp 1676037725
transform 1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1676037725
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1676037725
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1676037725
transform 1 0 17296 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1676037725
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1676037725
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_87
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_92
timestamp 1676037725
transform 1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_191
timestamp 1676037725
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_204
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_220
timestamp 1676037725
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_224
timestamp 1676037725
transform 1 0 21712 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_255
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1676037725
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_13
timestamp 1676037725
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_37
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1676037725
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1676037725
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1676037725
transform 1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_150
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1676037725
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_187
timestamp 1676037725
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1676037725
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_208
timestamp 1676037725
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1676037725
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1676037725
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_46
timestamp 1676037725
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1676037725
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1676037725
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_124
timestamp 1676037725
transform 1 0 12512 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_152
timestamp 1676037725
transform 1 0 15088 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_156
timestamp 1676037725
transform 1 0 15456 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_168
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1676037725
transform 1 0 18400 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1676037725
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_199
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_207
timestamp 1676037725
transform 1 0 20148 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_210
timestamp 1676037725
transform 1 0 20424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_222
timestamp 1676037725
transform 1 0 21528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1676037725
transform 1 0 22264 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1676037725
transform 1 0 9568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_139
timestamp 1676037725
transform 1 0 13892 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1676037725
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1676037725
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 1676037725
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_203
timestamp 1676037725
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_215
timestamp 1676037725
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_244
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_13
timestamp 1676037725
transform 1 0 2300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_17
timestamp 1676037725
transform 1 0 2668 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_35
timestamp 1676037725
transform 1 0 4324 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_59
timestamp 1676037725
transform 1 0 6532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1676037725
transform 1 0 7636 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1676037725
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1676037725
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1676037725
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_135
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_160
timestamp 1676037725
transform 1 0 15824 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_166
timestamp 1676037725
transform 1 0 16376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_184
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1676037725
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_228
timestamp 1676037725
transform 1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1676037725
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1676037725
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_132
timestamp 1676037725
transform 1 0 13248 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1676037725
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_148
timestamp 1676037725
transform 1 0 14720 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_174
timestamp 1676037725
transform 1 0 17112 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_183
timestamp 1676037725
transform 1 0 17940 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_192
timestamp 1676037725
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1676037725
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_208
timestamp 1676037725
transform 1 0 20240 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_211
timestamp 1676037725
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_37
timestamp 1676037725
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_49
timestamp 1676037725
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1676037725
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1676037725
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 1676037725
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1676037725
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_129
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_169
timestamp 1676037725
transform 1 0 16652 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1676037725
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_259
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_25
timestamp 1676037725
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_37
timestamp 1676037725
transform 1 0 4508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_61
timestamp 1676037725
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1676037725
transform 1 0 7636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_90
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1676037725
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_116
timestamp 1676037725
transform 1 0 11776 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_127
timestamp 1676037725
transform 1 0 12788 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_133
timestamp 1676037725
transform 1 0 13340 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_157
timestamp 1676037725
transform 1 0 15548 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_177
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_180
timestamp 1676037725
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1676037725
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_210
timestamp 1676037725
transform 1 0 20424 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1676037725
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_263
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1676037725
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1676037725
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_17
timestamp 1676037725
transform 1 0 2668 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_47
timestamp 1676037725
transform 1 0 5428 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_71
timestamp 1676037725
transform 1 0 7636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1676037725
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1676037725
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_107
timestamp 1676037725
transform 1 0 10948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_120
timestamp 1676037725
transform 1 0 12144 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1676037725
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_187
timestamp 1676037725
transform 1 0 18308 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1676037725
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_21
timestamp 1676037725
transform 1 0 3036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_33
timestamp 1676037725
transform 1 0 4140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_59
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1676037725
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1676037725
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_102
timestamp 1676037725
transform 1 0 10488 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1676037725
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1676037725
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_140
timestamp 1676037725
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_152
timestamp 1676037725
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1676037725
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_176
timestamp 1676037725
transform 1 0 17296 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_215
timestamp 1676037725
transform 1 0 20884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_257
timestamp 1676037725
transform 1 0 24748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_13
timestamp 1676037725
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_18
timestamp 1676037725
transform 1 0 2760 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_51
timestamp 1676037725
transform 1 0 5796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_58
timestamp 1676037725
transform 1 0 6440 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1676037725
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1676037725
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_99
timestamp 1676037725
transform 1 0 10212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1676037725
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1676037725
transform 1 0 13432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1676037725
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_175
timestamp 1676037725
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_182
timestamp 1676037725
transform 1 0 17848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1676037725
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1676037725
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_48
timestamp 1676037725
transform 1 0 5520 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1676037725
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_65
timestamp 1676037725
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1676037725
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1676037725
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1676037725
transform 1 0 13248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_143
timestamp 1676037725
transform 1 0 14260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_147
timestamp 1676037725
transform 1 0 14628 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1676037725
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_206
timestamp 1676037725
transform 1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_257
timestamp 1676037725
transform 1 0 24748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_34
timestamp 1676037725
transform 1 0 4232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_46
timestamp 1676037725
transform 1 0 5336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1676037725
transform 1 0 6440 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1676037725
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_87
timestamp 1676037725
transform 1 0 9108 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1676037725
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_106
timestamp 1676037725
transform 1 0 10856 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_110
timestamp 1676037725
transform 1 0 11224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1676037725
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_147
timestamp 1676037725
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_157
timestamp 1676037725
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_181
timestamp 1676037725
transform 1 0 17756 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_187
timestamp 1676037725
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_208
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_220
timestamp 1676037725
transform 1 0 21344 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 1676037725
transform 1 0 22908 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_243
timestamp 1676037725
transform 1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_263
timestamp 1676037725
transform 1 0 25300 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_14
timestamp 1676037725
transform 1 0 2392 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_20
timestamp 1676037725
transform 1 0 2944 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_29
timestamp 1676037725
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_78
timestamp 1676037725
transform 1 0 8280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_82
timestamp 1676037725
transform 1 0 8648 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_86
timestamp 1676037725
transform 1 0 9016 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1676037725
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1676037725
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1676037725
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_121
timestamp 1676037725
transform 1 0 12236 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_146
timestamp 1676037725
transform 1 0 14536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_150
timestamp 1676037725
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_154
timestamp 1676037725
transform 1 0 15272 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1676037725
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_177
timestamp 1676037725
transform 1 0 17388 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_200
timestamp 1676037725
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1676037725
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1676037725
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_33
timestamp 1676037725
transform 1 0 4140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_45
timestamp 1676037725
transform 1 0 5244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_57
timestamp 1676037725
transform 1 0 6348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_78
timestamp 1676037725
transform 1 0 8280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_90
timestamp 1676037725
transform 1 0 9384 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1676037725
transform 1 0 11776 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1676037725
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_146
timestamp 1676037725
transform 1 0 14536 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_154
timestamp 1676037725
transform 1 0 15272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_175
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_181
timestamp 1676037725
transform 1 0 17756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1676037725
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_208
timestamp 1676037725
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1676037725
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_259
timestamp 1676037725
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_263
timestamp 1676037725
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1676037725
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1676037725
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_79
timestamp 1676037725
transform 1 0 8372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_92
timestamp 1676037725
transform 1 0 9568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1676037725
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1676037725
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_144
timestamp 1676037725
transform 1 0 14352 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_157
timestamp 1676037725
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1676037725
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_177
timestamp 1676037725
transform 1 0 17388 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_188
timestamp 1676037725
transform 1 0 18400 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1676037725
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1676037725
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_232
timestamp 1676037725
transform 1 0 22448 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_75
timestamp 1676037725
transform 1 0 8004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1676037725
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_129
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_149
timestamp 1676037725
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_161
timestamp 1676037725
transform 1 0 15916 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_167
timestamp 1676037725
transform 1 0 16468 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_179
timestamp 1676037725
transform 1 0 17572 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_188
timestamp 1676037725
transform 1 0 18400 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1676037725
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_204
timestamp 1676037725
transform 1 0 19872 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1676037725
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_223
timestamp 1676037725
transform 1 0 21620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_247
timestamp 1676037725
transform 1 0 23828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_259
timestamp 1676037725
transform 1 0 24932 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_263
timestamp 1676037725
transform 1 0 25300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_9
timestamp 1676037725
transform 1 0 1932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_13
timestamp 1676037725
transform 1 0 2300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_25
timestamp 1676037725
transform 1 0 3404 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1676037725
transform 1 0 3864 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_42
timestamp 1676037725
transform 1 0 4968 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1676037725
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_77
timestamp 1676037725
transform 1 0 8188 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_98
timestamp 1676037725
transform 1 0 10120 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1676037725
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1676037725
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_128
timestamp 1676037725
transform 1 0 12880 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_146
timestamp 1676037725
transform 1 0 14536 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_154
timestamp 1676037725
transform 1 0 15272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_175
timestamp 1676037725
transform 1 0 17204 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_204
timestamp 1676037725
transform 1 0 19872 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_208
timestamp 1676037725
transform 1 0 20240 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_248
timestamp 1676037725
transform 1 0 23920 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_252
timestamp 1676037725
transform 1 0 24288 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1676037725
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_265
timestamp 1676037725
transform 1 0 25484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_33
timestamp 1676037725
transform 1 0 4140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_55
timestamp 1676037725
transform 1 0 6164 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_79
timestamp 1676037725
transform 1 0 8372 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_123
timestamp 1676037725
transform 1 0 12420 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_152
timestamp 1676037725
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_156
timestamp 1676037725
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_167
timestamp 1676037725
transform 1 0 16468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1676037725
transform 1 0 16836 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1676037725
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_219
timestamp 1676037725
transform 1 0 21252 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_223
timestamp 1676037725
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_235
timestamp 1676037725
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1676037725
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_258
timestamp 1676037725
transform 1 0 24840 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_92
timestamp 1676037725
transform 1 0 9568 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_96
timestamp 1676037725
transform 1 0 9936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1676037725
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_121
timestamp 1676037725
transform 1 0 12236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_133
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1676037725
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_159
timestamp 1676037725
transform 1 0 15732 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_165
timestamp 1676037725
transform 1 0 16284 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_186
timestamp 1676037725
transform 1 0 18216 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_198
timestamp 1676037725
transform 1 0 19320 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_204
timestamp 1676037725
transform 1 0 19872 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_215
timestamp 1676037725
transform 1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_246
timestamp 1676037725
transform 1 0 23736 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_251
timestamp 1676037725
transform 1 0 24196 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_259
timestamp 1676037725
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 1676037725
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_55
timestamp 1676037725
transform 1 0 6164 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp 1676037725
transform 1 0 7636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1676037725
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_89
timestamp 1676037725
transform 1 0 9292 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_100
timestamp 1676037725
transform 1 0 10304 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_134
timestamp 1676037725
transform 1 0 13432 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1676037725
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_181
timestamp 1676037725
transform 1 0 17756 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1676037725
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_210
timestamp 1676037725
transform 1 0 20424 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_214
timestamp 1676037725
transform 1 0 20792 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1676037725
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_231
timestamp 1676037725
transform 1 0 22356 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1676037725
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_87
timestamp 1676037725
transform 1 0 9108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_95
timestamp 1676037725
transform 1 0 9844 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1676037725
transform 1 0 10212 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_118
timestamp 1676037725
transform 1 0 11960 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1676037725
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_188
timestamp 1676037725
transform 1 0 18400 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1676037725
transform 1 0 18952 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_198
timestamp 1676037725
transform 1 0 19320 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1676037725
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1676037725
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_241
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_52
timestamp 1676037725
transform 1 0 5888 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_64
timestamp 1676037725
transform 1 0 6992 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_72
timestamp 1676037725
transform 1 0 7728 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1676037725
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_112
timestamp 1676037725
transform 1 0 11408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1676037725
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_120
timestamp 1676037725
transform 1 0 12144 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_125
timestamp 1676037725
transform 1 0 12604 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_136
timestamp 1676037725
transform 1 0 13616 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_162
timestamp 1676037725
transform 1 0 16008 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_184
timestamp 1676037725
transform 1 0 18032 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1676037725
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_208
timestamp 1676037725
transform 1 0 20240 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_212
timestamp 1676037725
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_224
timestamp 1676037725
transform 1 0 21712 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_236
timestamp 1676037725
transform 1 0 22816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_244
timestamp 1676037725
transform 1 0 23552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1676037725
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_259
timestamp 1676037725
transform 1 0 24932 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1676037725
transform 1 0 7268 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_78
timestamp 1676037725
transform 1 0 8280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_91
timestamp 1676037725
transform 1 0 9476 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_95
timestamp 1676037725
transform 1 0 9844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1676037725
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_148
timestamp 1676037725
transform 1 0 14720 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_152
timestamp 1676037725
transform 1 0 15088 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1676037725
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_172
timestamp 1676037725
transform 1 0 16928 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_183
timestamp 1676037725
transform 1 0 17940 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1676037725
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_209
timestamp 1676037725
transform 1 0 20332 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_215
timestamp 1676037725
transform 1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1676037725
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1676037725
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_75
timestamp 1676037725
transform 1 0 8004 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1676037725
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1676037725
transform 1 0 9200 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_110
timestamp 1676037725
transform 1 0 11224 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_114
timestamp 1676037725
transform 1 0 11592 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_126
timestamp 1676037725
transform 1 0 12696 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_134
timestamp 1676037725
transform 1 0 13432 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_152
timestamp 1676037725
transform 1 0 15088 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_164
timestamp 1676037725
transform 1 0 16192 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_175
timestamp 1676037725
transform 1 0 17204 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1676037725
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_225
timestamp 1676037725
transform 1 0 21804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_235
timestamp 1676037725
transform 1 0 22724 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_35
timestamp 1676037725
transform 1 0 4324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_40
timestamp 1676037725
transform 1 0 4784 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_66
timestamp 1676037725
transform 1 0 7176 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1676037725
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1676037725
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_102
timestamp 1676037725
transform 1 0 10488 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1676037725
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_116
timestamp 1676037725
transform 1 0 11776 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1676037725
transform 1 0 12788 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_134
timestamp 1676037725
transform 1 0 13432 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_180
timestamp 1676037725
transform 1 0 17664 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_199
timestamp 1676037725
transform 1 0 19412 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_209
timestamp 1676037725
transform 1 0 20332 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_227
timestamp 1676037725
transform 1 0 21988 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_232
timestamp 1676037725
transform 1 0 22448 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_243
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_255
timestamp 1676037725
transform 1 0 24564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_259
timestamp 1676037725
transform 1 0 24932 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1676037725
transform 1 0 25392 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1676037725
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_89
timestamp 1676037725
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1676037725
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1676037725
transform 1 0 10948 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_118
timestamp 1676037725
transform 1 0 11960 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_122
timestamp 1676037725
transform 1 0 12328 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_134
timestamp 1676037725
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_152
timestamp 1676037725
transform 1 0 15088 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_158
timestamp 1676037725
transform 1 0 15640 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_161
timestamp 1676037725
transform 1 0 15916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_172
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_178
timestamp 1676037725
transform 1 0 17480 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_184
timestamp 1676037725
transform 1 0 18032 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_201
timestamp 1676037725
transform 1 0 19596 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_212
timestamp 1676037725
transform 1 0 20608 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_225
timestamp 1676037725
transform 1 0 21804 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_232
timestamp 1676037725
transform 1 0 22448 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_238
timestamp 1676037725
transform 1 0 23000 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_259
timestamp 1676037725
transform 1 0 24932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_8
timestamp 1676037725
transform 1 0 1840 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_12
timestamp 1676037725
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_24
timestamp 1676037725
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_36
timestamp 1676037725
transform 1 0 4416 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_44
timestamp 1676037725
transform 1 0 5152 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_49
timestamp 1676037725
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_67
timestamp 1676037725
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_79
timestamp 1676037725
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_91
timestamp 1676037725
transform 1 0 9476 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_97
timestamp 1676037725
transform 1 0 10028 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1676037725
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_121
timestamp 1676037725
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1676037725
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_204
timestamp 1676037725
transform 1 0 19872 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1676037725
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_230
timestamp 1676037725
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_47
timestamp 1676037725
transform 1 0 5428 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_68
timestamp 1676037725
transform 1 0 7360 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_74
timestamp 1676037725
transform 1 0 7912 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1676037725
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1676037725
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_100
timestamp 1676037725
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_125
timestamp 1676037725
transform 1 0 12604 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_143
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_155
timestamp 1676037725
transform 1 0 15364 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_181
timestamp 1676037725
transform 1 0 17756 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1676037725
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_193
timestamp 1676037725
transform 1 0 18860 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_208
timestamp 1676037725
transform 1 0 20240 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_214
timestamp 1676037725
transform 1 0 20792 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1676037725
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_239
timestamp 1676037725
transform 1 0 23092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_243
timestamp 1676037725
transform 1 0 23460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_258
timestamp 1676037725
transform 1 0 24840 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_80
timestamp 1676037725
transform 1 0 8464 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_104
timestamp 1676037725
transform 1 0 10672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1676037725
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_135
timestamp 1676037725
transform 1 0 13524 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_139
timestamp 1676037725
transform 1 0 13892 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_151
timestamp 1676037725
transform 1 0 14996 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_210
timestamp 1676037725
transform 1 0 20424 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1676037725
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_236
timestamp 1676037725
transform 1 0 22816 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_256
timestamp 1676037725
transform 1 0 24656 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_260
timestamp 1676037725
transform 1 0 25024 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_74
timestamp 1676037725
transform 1 0 7912 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1676037725
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_98
timestamp 1676037725
transform 1 0 10120 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_110
timestamp 1676037725
transform 1 0 11224 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_122
timestamp 1676037725
transform 1 0 12328 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_128
timestamp 1676037725
transform 1 0 12880 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_175
timestamp 1676037725
transform 1 0 17204 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_179
timestamp 1676037725
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1676037725
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_219
timestamp 1676037725
transform 1 0 21252 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1676037725
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1676037725
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_255
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_59
timestamp 1676037725
transform 1 0 6532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1676037725
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_75
timestamp 1676037725
transform 1 0 8004 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_96
timestamp 1676037725
transform 1 0 9936 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1676037725
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1676037725
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_148
timestamp 1676037725
transform 1 0 14720 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_160
timestamp 1676037725
transform 1 0 15824 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_177
timestamp 1676037725
transform 1 0 17388 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_212
timestamp 1676037725
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1676037725
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_235
timestamp 1676037725
transform 1 0 22724 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_8
timestamp 1676037725
transform 1 0 1840 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_12
timestamp 1676037725
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1676037725
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1676037725
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_96
timestamp 1676037725
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_108
timestamp 1676037725
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_124
timestamp 1676037725
transform 1 0 12512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_135
timestamp 1676037725
transform 1 0 13524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_152
timestamp 1676037725
transform 1 0 15088 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_158
timestamp 1676037725
transform 1 0 15640 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_161
timestamp 1676037725
transform 1 0 15916 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_172
timestamp 1676037725
transform 1 0 16928 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_179
timestamp 1676037725
transform 1 0 17572 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_191
timestamp 1676037725
transform 1 0 18676 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_208
timestamp 1676037725
transform 1 0 20240 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_223
timestamp 1676037725
transform 1 0 21620 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_235
timestamp 1676037725
transform 1 0 22724 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_250
timestamp 1676037725
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1676037725
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_84
timestamp 1676037725
transform 1 0 8832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_95
timestamp 1676037725
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_115
timestamp 1676037725
transform 1 0 11684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_129
timestamp 1676037725
transform 1 0 12972 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_142
timestamp 1676037725
transform 1 0 14168 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_155
timestamp 1676037725
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_171
timestamp 1676037725
transform 1 0 16836 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_182
timestamp 1676037725
transform 1 0 17848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_194
timestamp 1676037725
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_199
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_214
timestamp 1676037725
transform 1 0 20792 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1676037725
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_256
timestamp 1676037725
transform 1 0 24656 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_260
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_61
timestamp 1676037725
transform 1 0 6716 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1676037725
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_98
timestamp 1676037725
transform 1 0 10120 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_104
timestamp 1676037725
transform 1 0 10672 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_108
timestamp 1676037725
transform 1 0 11040 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_119
timestamp 1676037725
transform 1 0 12052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_126
timestamp 1676037725
transform 1 0 12696 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1676037725
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_148
timestamp 1676037725
transform 1 0 14720 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_159
timestamp 1676037725
transform 1 0 15732 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1676037725
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1676037725
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_192
timestamp 1676037725
transform 1 0 18768 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_210
timestamp 1676037725
transform 1 0 20424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_214
timestamp 1676037725
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_219
timestamp 1676037725
transform 1 0 21252 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_232
timestamp 1676037725
transform 1 0 22448 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_244
timestamp 1676037725
transform 1 0 23552 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_264
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1676037725
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_88
timestamp 1676037725
transform 1 0 9200 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_106
timestamp 1676037725
transform 1 0 10856 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_118
timestamp 1676037725
transform 1 0 11960 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_131
timestamp 1676037725
transform 1 0 13156 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_138
timestamp 1676037725
transform 1 0 13800 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_142
timestamp 1676037725
transform 1 0 14168 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_147
timestamp 1676037725
transform 1 0 14628 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_160
timestamp 1676037725
transform 1 0 15824 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_164
timestamp 1676037725
transform 1 0 16192 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_180
timestamp 1676037725
transform 1 0 17664 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1676037725
transform 1 0 18768 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_203
timestamp 1676037725
transform 1 0 19780 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_207
timestamp 1676037725
transform 1 0 20148 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_236
timestamp 1676037725
transform 1 0 22816 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1676037725
transform 1 0 23368 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_8
timestamp 1676037725
transform 1 0 1840 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_12
timestamp 1676037725
transform 1 0 2208 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1676037725
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_67
timestamp 1676037725
transform 1 0 7268 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_71
timestamp 1676037725
transform 1 0 7636 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1676037725
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_110
timestamp 1676037725
transform 1 0 11224 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_116
timestamp 1676037725
transform 1 0 11776 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_126
timestamp 1676037725
transform 1 0 12696 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_130
timestamp 1676037725
transform 1 0 13064 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_137
timestamp 1676037725
transform 1 0 13708 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_152
timestamp 1676037725
transform 1 0 15088 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_160
timestamp 1676037725
transform 1 0 15824 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_181
timestamp 1676037725
transform 1 0 17756 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 1676037725
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_208
timestamp 1676037725
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_225
timestamp 1676037725
transform 1 0 21804 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_236
timestamp 1676037725
transform 1 0 22816 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1676037725
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_65
timestamp 1676037725
transform 1 0 7084 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_75
timestamp 1676037725
transform 1 0 8004 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_84
timestamp 1676037725
transform 1 0 8832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_96
timestamp 1676037725
transform 1 0 9936 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_100
timestamp 1676037725
transform 1 0 10304 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1676037725
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_115
timestamp 1676037725
transform 1 0 11684 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_139
timestamp 1676037725
transform 1 0 13892 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_146
timestamp 1676037725
transform 1 0 14536 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1676037725
transform 1 0 15732 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_163
timestamp 1676037725
transform 1 0 16100 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_174
timestamp 1676037725
transform 1 0 17112 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1676037725
transform 1 0 17848 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_192
timestamp 1676037725
transform 1 0 18768 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1676037725
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_248
timestamp 1676037725
transform 1 0 23920 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_252
timestamp 1676037725
transform 1 0 24288 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1676037725
transform 1 0 24748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_264
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_61
timestamp 1676037725
transform 1 0 6716 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_67
timestamp 1676037725
transform 1 0 7268 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_79
timestamp 1676037725
transform 1 0 8372 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_90
timestamp 1676037725
transform 1 0 9384 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_103
timestamp 1676037725
transform 1 0 10580 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_127
timestamp 1676037725
transform 1 0 12788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_137
timestamp 1676037725
transform 1 0 13708 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_166
timestamp 1676037725
transform 1 0 16376 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_178
timestamp 1676037725
transform 1 0 17480 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 1676037725
transform 1 0 20240 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_212
timestamp 1676037725
transform 1 0 20608 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_218
timestamp 1676037725
transform 1 0 21160 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_228
timestamp 1676037725
transform 1 0 22080 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_232
timestamp 1676037725
transform 1 0 22448 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_243
timestamp 1676037725
transform 1 0 23460 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1676037725
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_65
timestamp 1676037725
transform 1 0 7084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_76
timestamp 1676037725
transform 1 0 8096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_103
timestamp 1676037725
transform 1 0 10580 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1676037725
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_115
timestamp 1676037725
transform 1 0 11684 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_123
timestamp 1676037725
transform 1 0 12420 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_127
timestamp 1676037725
transform 1 0 12788 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_148
timestamp 1676037725
transform 1 0 14720 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_152
timestamp 1676037725
transform 1 0 15088 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_156
timestamp 1676037725
transform 1 0 15456 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_166
timestamp 1676037725
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_171
timestamp 1676037725
transform 1 0 16836 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_183
timestamp 1676037725
transform 1 0 17940 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_195
timestamp 1676037725
transform 1 0 19044 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_212
timestamp 1676037725
transform 1 0 20608 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 1676037725
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_229
timestamp 1676037725
transform 1 0 22172 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_234
timestamp 1676037725
transform 1 0 22632 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_242
timestamp 1676037725
transform 1 0 23368 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_75
timestamp 1676037725
transform 1 0 8004 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_79
timestamp 1676037725
transform 1 0 8372 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_101
timestamp 1676037725
transform 1 0 10396 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_105
timestamp 1676037725
transform 1 0 10764 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_134
timestamp 1676037725
transform 1 0 13432 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_138
timestamp 1676037725
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1676037725
transform 1 0 14996 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_162
timestamp 1676037725
transform 1 0 16008 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_166
timestamp 1676037725
transform 1 0 16376 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_178
timestamp 1676037725
transform 1 0 17480 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1676037725
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_205
timestamp 1676037725
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_210
timestamp 1676037725
transform 1 0 20424 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_214
timestamp 1676037725
transform 1 0 20792 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_224
timestamp 1676037725
transform 1 0 21712 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_230
timestamp 1676037725
transform 1 0 22264 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_241
timestamp 1676037725
transform 1 0 23276 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_247
timestamp 1676037725
transform 1 0 23828 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_259
timestamp 1676037725
transform 1 0 24932 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_264
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_8
timestamp 1676037725
transform 1 0 1840 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_12
timestamp 1676037725
transform 1 0 2208 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_20
timestamp 1676037725
transform 1 0 2944 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_26
timestamp 1676037725
transform 1 0 3496 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_30
timestamp 1676037725
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_42
timestamp 1676037725
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1676037725
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_77
timestamp 1676037725
transform 1 0 8188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_109
timestamp 1676037725
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_124
timestamp 1676037725
transform 1 0 12512 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_156
timestamp 1676037725
transform 1 0 15456 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_160
timestamp 1676037725
transform 1 0 15824 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_191
timestamp 1676037725
transform 1 0 18676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_197
timestamp 1676037725
transform 1 0 19228 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_208
timestamp 1676037725
transform 1 0 20240 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_212
timestamp 1676037725
transform 1 0 20608 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_222
timestamp 1676037725
transform 1 0 21528 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_230
timestamp 1676037725
transform 1 0 22264 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_257
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_46
timestamp 1676037725
transform 1 0 5336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_50
timestamp 1676037725
transform 1 0 5704 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_72
timestamp 1676037725
transform 1 0 7728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_78
timestamp 1676037725
transform 1 0 8280 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_100
timestamp 1676037725
transform 1 0 10304 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_113
timestamp 1676037725
transform 1 0 11500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_117
timestamp 1676037725
transform 1 0 11868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_129
timestamp 1676037725
transform 1 0 12972 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_161
timestamp 1676037725
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_173
timestamp 1676037725
transform 1 0 17020 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1676037725
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_219
timestamp 1676037725
transform 1 0 21252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_232
timestamp 1676037725
transform 1 0 22448 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_249
timestamp 1676037725
transform 1 0 24012 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_31
timestamp 1676037725
transform 1 0 3956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_37
timestamp 1676037725
transform 1 0 4508 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1676037725
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_63
timestamp 1676037725
transform 1 0 6900 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_67
timestamp 1676037725
transform 1 0 7268 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_102
timestamp 1676037725
transform 1 0 10488 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_106
timestamp 1676037725
transform 1 0 10856 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_138
timestamp 1676037725
transform 1 0 13800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_145
timestamp 1676037725
transform 1 0 14444 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_153
timestamp 1676037725
transform 1 0 15180 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_164
timestamp 1676037725
transform 1 0 16192 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_180
timestamp 1676037725
transform 1 0 17664 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_73_186
timestamp 1676037725
transform 1 0 18216 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_191
timestamp 1676037725
transform 1 0 18676 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_204
timestamp 1676037725
transform 1 0 19872 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_221
timestamp 1676037725
transform 1 0 21436 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_238
timestamp 1676037725
transform 1 0 23000 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_242
timestamp 1676037725
transform 1 0 23368 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_263
timestamp 1676037725
transform 1 0 25300 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_37
timestamp 1676037725
transform 1 0 4508 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_43
timestamp 1676037725
transform 1 0 5060 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_47
timestamp 1676037725
transform 1 0 5428 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_59
timestamp 1676037725
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_71
timestamp 1676037725
transform 1 0 7636 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_79
timestamp 1676037725
transform 1 0 8372 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_93
timestamp 1676037725
transform 1 0 9660 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_101
timestamp 1676037725
transform 1 0 10396 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_125
timestamp 1676037725
transform 1 0 12604 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_129
timestamp 1676037725
transform 1 0 12972 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_137
timestamp 1676037725
transform 1 0 13708 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_145
timestamp 1676037725
transform 1 0 14444 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_169
timestamp 1676037725
transform 1 0 16652 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_173
timestamp 1676037725
transform 1 0 17020 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_183
timestamp 1676037725
transform 1 0 17940 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_220
timestamp 1676037725
transform 1 0 21344 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_224
timestamp 1676037725
transform 1 0 21712 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_234
timestamp 1676037725
transform 1 0 22632 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_74_250
timestamp 1676037725
transform 1 0 24104 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_255
timestamp 1676037725
transform 1 0 24564 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1676037725
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1676037725
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1676037725
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1676037725
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_75
timestamp 1676037725
transform 1 0 8004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_83
timestamp 1676037725
transform 1 0 8740 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_96
timestamp 1676037725
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_100
timestamp 1676037725
transform 1 0 10304 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1676037725
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1676037725
transform 1 0 12236 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_143
timestamp 1676037725
transform 1 0 14260 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_156
timestamp 1676037725
transform 1 0 15456 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_160
timestamp 1676037725
transform 1 0 15824 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_171
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_182
timestamp 1676037725
transform 1 0 17848 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_186
timestamp 1676037725
transform 1 0 18216 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_207
timestamp 1676037725
transform 1 0 20148 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_211
timestamp 1676037725
transform 1 0 20516 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_219
timestamp 1676037725
transform 1 0 21252 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_236
timestamp 1676037725
transform 1 0 22816 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_59
timestamp 1676037725
transform 1 0 6532 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_64
timestamp 1676037725
transform 1 0 6992 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_68
timestamp 1676037725
transform 1 0 7360 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_76
timestamp 1676037725
transform 1 0 8096 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_82
timestamp 1676037725
transform 1 0 8648 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_108
timestamp 1676037725
transform 1 0 11040 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_116
timestamp 1676037725
transform 1 0 11776 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_120
timestamp 1676037725
transform 1 0 12144 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_132
timestamp 1676037725
transform 1 0 13248 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_181
timestamp 1676037725
transform 1 0 17756 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_184
timestamp 1676037725
transform 1 0 18032 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_225
timestamp 1676037725
transform 1 0 21804 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_236
timestamp 1676037725
transform 1 0 22816 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_248
timestamp 1676037725
transform 1 0 23920 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_261
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1676037725
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_63
timestamp 1676037725
transform 1 0 6900 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_71
timestamp 1676037725
transform 1 0 7636 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_78
timestamp 1676037725
transform 1 0 8280 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_77_88
timestamp 1676037725
transform 1 0 9200 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_92
timestamp 1676037725
transform 1 0 9568 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_104
timestamp 1676037725
transform 1 0 10672 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_110
timestamp 1676037725
transform 1 0 11224 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_115
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_126
timestamp 1676037725
transform 1 0 12696 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_130
timestamp 1676037725
transform 1 0 13064 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_157
timestamp 1676037725
transform 1 0 15548 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_165
timestamp 1676037725
transform 1 0 16284 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_191
timestamp 1676037725
transform 1 0 18676 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_195
timestamp 1676037725
transform 1 0 19044 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_199
timestamp 1676037725
transform 1 0 19412 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_220
timestamp 1676037725
transform 1 0 21344 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_229
timestamp 1676037725
transform 1 0 22172 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_250
timestamp 1676037725
transform 1 0 24104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_59
timestamp 1676037725
transform 1 0 6532 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_67
timestamp 1676037725
transform 1 0 7268 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_75
timestamp 1676037725
transform 1 0 8004 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1676037725
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_91
timestamp 1676037725
transform 1 0 9476 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_95
timestamp 1676037725
transform 1 0 9844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_110
timestamp 1676037725
transform 1 0 11224 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_116
timestamp 1676037725
transform 1 0 11776 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_120
timestamp 1676037725
transform 1 0 12144 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_138
timestamp 1676037725
transform 1 0 13800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_149
timestamp 1676037725
transform 1 0 14812 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_172
timestamp 1676037725
transform 1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_176
timestamp 1676037725
transform 1 0 17296 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_188
timestamp 1676037725
transform 1 0 18400 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_78_220
timestamp 1676037725
transform 1 0 21344 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_224
timestamp 1676037725
transform 1 0 21712 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1676037725
transform 1 0 24104 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_255
timestamp 1676037725
transform 1 0 24564 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_263
timestamp 1676037725
transform 1 0 25300 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_5
timestamp 1676037725
transform 1 0 1564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_17
timestamp 1676037725
transform 1 0 2668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_29
timestamp 1676037725
transform 1 0 3772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_41
timestamp 1676037725
transform 1 0 4876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1676037725
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_86
timestamp 1676037725
transform 1 0 9016 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_108
timestamp 1676037725
transform 1 0 11040 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_115
timestamp 1676037725
transform 1 0 11684 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_121
timestamp 1676037725
transform 1 0 12236 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_133
timestamp 1676037725
transform 1 0 13340 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_141
timestamp 1676037725
transform 1 0 14076 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_164
timestamp 1676037725
transform 1 0 16192 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_187
timestamp 1676037725
transform 1 0 18308 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_208
timestamp 1676037725
transform 1 0 20240 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_212
timestamp 1676037725
transform 1 0 20608 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_215
timestamp 1676037725
transform 1 0 20884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_247
timestamp 1676037725
transform 1 0 23828 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_79_251
timestamp 1676037725
transform 1 0 24196 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1676037725
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_78
timestamp 1676037725
transform 1 0 8280 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_90
timestamp 1676037725
transform 1 0 9384 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_96
timestamp 1676037725
transform 1 0 9936 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_100
timestamp 1676037725
transform 1 0 10304 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_113
timestamp 1676037725
transform 1 0 11500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1676037725
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_143
timestamp 1676037725
transform 1 0 14260 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_155
timestamp 1676037725
transform 1 0 15364 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_163
timestamp 1676037725
transform 1 0 16100 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_168
timestamp 1676037725
transform 1 0 16560 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_180
timestamp 1676037725
transform 1 0 17664 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_188
timestamp 1676037725
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_193
timestamp 1676037725
transform 1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_200
timestamp 1676037725
transform 1 0 19504 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_211
timestamp 1676037725
transform 1 0 20516 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_224
timestamp 1676037725
transform 1 0 21712 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_236
timestamp 1676037725
transform 1 0 22816 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1676037725
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_255
timestamp 1676037725
transform 1 0 24564 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_263
timestamp 1676037725
transform 1 0 25300 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_65
timestamp 1676037725
transform 1 0 7084 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_109
timestamp 1676037725
transform 1 0 11132 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1676037725
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1676037725
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_191
timestamp 1676037725
transform 1 0 18676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_215
timestamp 1676037725
transform 1 0 20884 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 1676037725
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_228
timestamp 1676037725
transform 1 0 22080 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_239
timestamp 1676037725
transform 1 0 23092 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_243
timestamp 1676037725
transform 1 0 23460 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_251
timestamp 1676037725
transform 1 0 24196 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_93
timestamp 1676037725
transform 1 0 9660 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_119
timestamp 1676037725
transform 1 0 12052 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_123
timestamp 1676037725
transform 1 0 12420 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1676037725
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_144
timestamp 1676037725
transform 1 0 14352 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_156
timestamp 1676037725
transform 1 0 15456 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_178
timestamp 1676037725
transform 1 0 17480 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_182
timestamp 1676037725
transform 1 0 17848 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1676037725
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_199
timestamp 1676037725
transform 1 0 19412 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_211
timestamp 1676037725
transform 1 0 20516 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_225
timestamp 1676037725
transform 1 0 21804 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_236
timestamp 1676037725
transform 1 0 22816 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1676037725
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_259
timestamp 1676037725
transform 1 0 24932 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_264
timestamp 1676037725
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_90
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_102
timestamp 1676037725
transform 1 0 10488 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1676037725
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_180
timestamp 1676037725
transform 1 0 17664 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_197
timestamp 1676037725
transform 1 0 19228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_209
timestamp 1676037725
transform 1 0 20332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_221
timestamp 1676037725
transform 1 0 21436 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_253
timestamp 1676037725
transform 1 0 24380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1676037725
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1676037725
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_182
timestamp 1676037725
transform 1 0 17848 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1676037725
transform 1 0 18952 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_129
timestamp 1676037725
transform 1 0 12972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_141
timestamp 1676037725
transform 1 0 14076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_153
timestamp 1676037725
transform 1 0 15180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_165
timestamp 1676037725
transform 1 0 16284 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_25
timestamp 1676037725
transform 1 0 3404 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_113
timestamp 1676037725
transform 1 0 11500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_117
timestamp 1676037725
transform 1 0 11868 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_129
timestamp 1676037725
transform 1 0 12972 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_86_137
timestamp 1676037725
transform 1 0 13708 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_259
timestamp 1676037725
transform 1 0 24932 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_25
timestamp 1676037725
transform 1 0 3404 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1676037725
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_61
timestamp 1676037725
transform 1 0 6716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_73
timestamp 1676037725
transform 1 0 7820 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_85
timestamp 1676037725
transform 1 0 8924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_90
timestamp 1676037725
transform 1 0 9384 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_102
timestamp 1676037725
transform 1 0 10488 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_110
timestamp 1676037725
transform 1 0 11224 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 1676037725
transform 1 0 3496 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_45
timestamp 1676037725
transform 1 0 5244 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_57
timestamp 1676037725
transform 1 0 6348 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_61
timestamp 1676037725
transform 1 0 6716 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_91
timestamp 1676037725
transform 1 0 9476 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_103
timestamp 1676037725
transform 1 0 10580 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_115
timestamp 1676037725
transform 1 0 11684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_127
timestamp 1676037725
transform 1 0 12788 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1676037725
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_8
timestamp 1676037725
transform 1 0 1840 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_12
timestamp 1676037725
transform 1 0 2208 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_29
timestamp 1676037725
transform 1 0 3772 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1676037725
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_65
timestamp 1676037725
transform 1 0 7084 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_79
timestamp 1676037725
transform 1 0 8372 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_87
timestamp 1676037725
transform 1 0 9108 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_255
timestamp 1676037725
transform 1 0 24564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_258
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 1676037725
transform 1 0 3496 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_39
timestamp 1676037725
transform 1 0 4692 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_61
timestamp 1676037725
transform 1 0 6716 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_102
timestamp 1676037725
transform 1 0 10488 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_114
timestamp 1676037725
transform 1 0 11592 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_126
timestamp 1676037725
transform 1 0 12696 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1676037725
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_259
timestamp 1676037725
transform 1 0 24932 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_13
timestamp 1676037725
transform 1 0 2300 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_17
timestamp 1676037725
transform 1 0 2668 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_34
timestamp 1676037725
transform 1 0 4232 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_54
timestamp 1676037725
transform 1 0 6072 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_61
timestamp 1676037725
transform 1 0 6716 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_66
timestamp 1676037725
transform 1 0 7176 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_72
timestamp 1676037725
transform 1 0 7728 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_89
timestamp 1676037725
transform 1 0 9292 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_91_109
timestamp 1676037725
transform 1 0 11132 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_118
timestamp 1676037725
transform 1 0 11960 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_91_133
timestamp 1676037725
transform 1 0 13340 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_145
timestamp 1676037725
transform 1 0 14444 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_157
timestamp 1676037725
transform 1 0 15548 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_165
timestamp 1676037725
transform 1 0 16284 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_9
timestamp 1676037725
transform 1 0 1932 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 1676037725
transform 1 0 3496 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_45
timestamp 1676037725
transform 1 0 5244 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_128
timestamp 1676037725
transform 1 0 12880 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_132
timestamp 1676037725
transform 1 0 13248 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1676037725
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_143
timestamp 1676037725
transform 1 0 14260 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_155
timestamp 1676037725
transform 1 0 15364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_167
timestamp 1676037725
transform 1 0 16468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_179
timestamp 1676037725
transform 1 0 17572 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_191
timestamp 1676037725
transform 1 0 18676 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_258
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_14
timestamp 1676037725
transform 1 0 2392 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_34
timestamp 1676037725
transform 1 0 4232 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_73
timestamp 1676037725
transform 1 0 7820 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_90
timestamp 1676037725
transform 1 0 9384 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_133
timestamp 1676037725
transform 1 0 13340 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_141
timestamp 1676037725
transform 1 0 14076 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_148
timestamp 1676037725
transform 1 0 14720 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_152
timestamp 1676037725
transform 1 0 15088 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_160
timestamp 1676037725
transform 1 0 15824 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_164
timestamp 1676037725
transform 1 0 16192 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_93_177
timestamp 1676037725
transform 1 0 17388 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_189
timestamp 1676037725
transform 1 0 18492 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_196
timestamp 1676037725
transform 1 0 19136 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_204
timestamp 1676037725
transform 1 0 19872 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_208
timestamp 1676037725
transform 1 0 20240 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_212
timestamp 1676037725
transform 1 0 20608 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_220
timestamp 1676037725
transform 1 0 21344 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_93_227
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_93_232
timestamp 1676037725
transform 1 0 22448 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_235
timestamp 1676037725
transform 1 0 22724 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_239
timestamp 1676037725
transform 1 0 23092 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_244
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_251
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_255
timestamp 1676037725
transform 1 0 24564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1676037725
transform 1 0 24840 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_39
timestamp 1676037725
transform 1 0 4692 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1676037725
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1676037725
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_147
timestamp 1676037725
transform 1 0 14628 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_151
timestamp 1676037725
transform 1 0 14996 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_94_161
timestamp 1676037725
transform 1 0 15916 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_167
timestamp 1676037725
transform 1 0 16468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_173
timestamp 1676037725
transform 1 0 17020 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_180
timestamp 1676037725
transform 1 0 17664 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_184
timestamp 1676037725
transform 1 0 18032 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_203
timestamp 1676037725
transform 1 0 19780 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_211
timestamp 1676037725
transform 1 0 20516 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_228
timestamp 1676037725
transform 1 0 22080 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_235
timestamp 1676037725
transform 1 0 22724 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_257
timestamp 1676037725
transform 1 0 24748 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_33
timestamp 1676037725
transform 1 0 4140 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_118
timestamp 1676037725
transform 1 0 11960 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_143
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_147
timestamp 1676037725
transform 1 0 14628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_175
timestamp 1676037725
transform 1 0 17204 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_191
timestamp 1676037725
transform 1 0 18676 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_195
timestamp 1676037725
transform 1 0 19044 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_203
timestamp 1676037725
transform 1 0 19780 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_211
timestamp 1676037725
transform 1 0 20516 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_219
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_239
timestamp 1676037725
transform 1 0 23092 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_243
timestamp 1676037725
transform 1 0 23460 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_255
timestamp 1676037725
transform 1 0 24564 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1676037725
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 3956 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1676037725
transform 1 0 3036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1676037725
transform 1 0 1656 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1676037725
transform 1 0 1748 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 25116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 25116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 23184 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 24472 0 -1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 24472 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 24472 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 23184 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 24472 0 -1 47872
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 25116 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 25116 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23920 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 25116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7636 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1676037725
transform 1 0 9016 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 11684 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 16652 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 17572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 18124 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 19412 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 20148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 20148 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 20332 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 20884 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 21068 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 21804 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 22448 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1676037725
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 23092 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 23276 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 23920 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform 1 0 14260 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 14444 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 15548 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1676037725
transform 1 0 25024 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input100
timestamp 1676037725
transform 1 0 25024 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 25024 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform 1 0 23736 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1676037725
transform 1 0 3956 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input110
timestamp 1676037725
transform 1 0 3956 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__conb_1  left_tile_210
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 22632 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 23920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 23920 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 17572 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 19412 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 20516 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 22356 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 14628 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 14996 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 16836 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 1932 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 5336 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 7176 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 7820 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 2024 0 1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 7912 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 10764 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 11868 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 2300 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 2024 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2760 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 2024 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 2760 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 5244 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16192 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15364 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15916 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17572 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 20608 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16192 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14444 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14076 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 12880 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18032 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15364 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17572 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22172 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23552 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23552 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19504 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18308 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18400 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19044 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 16836 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15640 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15088 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14352 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 13616 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12880 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12052 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11684 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10396 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9568 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10580 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12512 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9936 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8280 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6164 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6440 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11500 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15364 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19872 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21712 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18216 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 3956 0 -1 50048
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10212 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11868 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13156 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 12328 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12328 0 -1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10948 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8924 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8464 0 -1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5428 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 5520 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 4232 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6532 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6164 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5244 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7544 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8832 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8096 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6072 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 3956 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6164 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 5888 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14812 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 15916 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11960 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15364 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 13892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__211
timestamp 1676037725
transform 1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 21988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20608 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__216
timestamp 1676037725
transform 1 0 17020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 13432 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__261
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14720 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17572 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 17572 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21528 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__263
timestamp 1676037725
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22080 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16100 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__264
timestamp 1676037725
transform 1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19780 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12788 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20332 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20792 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__213
timestamp 1676037725
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18308 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__215
timestamp 1676037725
transform 1 0 14352 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14996 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20976 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform 1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22908 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21252 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 23828 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23184 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19780 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22264 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20240 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__243
timestamp 1676037725
transform 1 0 22448 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23184 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24380 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20884 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18952 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21804 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 21620 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22448 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20884 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19780 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__218
timestamp 1676037725
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16100 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20608 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22172 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17020 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 16836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18216 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14352 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 14260 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16652 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16192 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 13524 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12880 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16100 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14628 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__224
timestamp 1676037725
transform 1 0 13156 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11960 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__225
timestamp 1676037725
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12604 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15088 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__226
timestamp 1676037725
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__227
timestamp 1676037725
transform 1 0 11960 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14720 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__228
timestamp 1676037725
transform 1 0 9384 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 8740 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__229
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__230
timestamp 1676037725
transform 1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7636 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__231
timestamp 1676037725
transform 1 0 10028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 8832 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10764 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 8188 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__233
timestamp 1676037725
transform 1 0 14720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__235
timestamp 1676037725
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__236
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20424 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__237
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__238
timestamp 1676037725
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23184 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__239
timestamp 1676037725
transform 1 0 20424 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__240
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21068 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22724 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17296 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__242
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14904 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__245
timestamp 1676037725
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10672 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11592 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12696 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15364 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__248
timestamp 1676037725
transform 1 0 14168 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12696 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10672 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__255
timestamp 1676037725
transform 1 0 9844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 8648 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9752 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9292 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 9108 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17296 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 12788 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__246
timestamp 1676037725
transform 1 0 7912 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8004 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7452 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__247
timestamp 1676037725
transform 1 0 6900 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7636 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 9476 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__249
timestamp 1676037725
transform 1 0 9752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9384 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9016 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12328 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12880 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__250
timestamp 1676037725
transform 1 0 5336 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 4968 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform -1 0 12236 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11868 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__251
timestamp 1676037725
transform 1 0 9108 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7176 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__253
timestamp 1676037725
transform 1 0 10948 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19136 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__254
timestamp 1676037725
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1490 56200 1546 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 16946 56200 17002 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 18418 56200 18474 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 19154 56200 19210 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 19890 56200 19946 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 13266 56200 13322 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 20626 56200 20682 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 21362 56200 21418 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 22098 56200 22154 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 23570 56200 23626 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 14002 56200 14058 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 14738 56200 14794 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 15474 56200 15530 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 5906 56200 5962 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 6642 56200 6698 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 8114 56200 8170 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 8850 56200 8906 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 9586 56200 9642 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 10322 56200 10378 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 11058 56200 11114 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 11794 56200 11850 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 2962 56200 3018 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 3698 56200 3754 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 4434 56200 4490 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 prog_reset
port 200 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reset
port 201 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 202 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 203 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 204 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 205 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 206 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 207 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 208 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 209 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 210 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 211 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 212 nsew signal tristate
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 213 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 test_enable
port 214 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal2 6026 24276 6026 24276 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal2 6210 25092 6210 25092 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 4508 23018 4508 23018 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 4232 19482 4232 19482 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 3450 20978 3450 20978 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 7498 19720 7498 19720 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal2 13386 20315 13386 20315 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 11592 18598 11592 18598 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 8326 20060 8326 20060 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal2 9430 16388 9430 16388 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 16008 16626 16008 16626 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 13156 18802 13156 18802 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 10810 14246 10810 14246 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 6900 17102 6900 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 16054 10948 16054 10948 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 12742 15334 12742 15334 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal2 8418 16354 8418 16354 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 14122 19244 14122 19244 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal2 12374 19822 12374 19822 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 8878 21590 8878 21590 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 12926 14586 12926 14586 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7912 21658 7912 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 6762 24174 6762 24174 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13570 16830 13570 16830 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14260 18938 14260 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12742 23018 12742 23018 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11730 19448 11730 19448 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11638 16218 11638 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 11730 20230 11730 20230 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8786 20876 8786 20876 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9246 21658 9246 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9476 20570 9476 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15226 15334 15226 15334 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9798 17306 9798 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 8280 17850 8280 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 14996 15470 14996 15470 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 18734 13662 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13846 18394 13846 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11040 16218 11040 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 14306 16184 14306 16184 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12719 18598 12719 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10350 16218 10350 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11270 17238 11270 17238 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 16762 10350 16762 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 14950 11322 14950 11322 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7084 17578 7084 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 6302 18598 6302 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13616 13294 13616 13294 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12282 18836 12282 18836 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12742 17034 12742 17034 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9338 19482 9338 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 12374 14688 12374 14688 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10580 16150 10580 16150 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7912 17714 7912 17714 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8878 16762 8878 16762 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8142 16218 8142 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12190 16660 12190 16660 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 6256 22746 6256 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 4784 22406 4784 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 13570 18734 13570 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 20264 14306 20264 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12052 21658 12052 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10442 19584 10442 19584 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11270 18122 11270 18122 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10810 21658 10810 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7590 21114 7590 21114 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 8004 22746 8004 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8234 21386 8234 21386 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 4278 24956 4278 24956 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 3036 25806 3036 25806 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal2 3450 26894 3450 26894 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel via1 3795 28186 3795 28186 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 4324 20502 4324 20502 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 2254 20876 2254 20876 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 3036 23290 3036 23290 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 3565 27098 3565 27098 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 5796 20230 5796 20230 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 3634 20400 3634 20400 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 2254 23052 2254 23052 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 4071 25126 4071 25126 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 4094 16728 4094 16728 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 3036 21114 3036 21114 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 4301 23086 4301 23086 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 2338 55420 2338 55420 0 ccff_head
rlabel metal1 1472 2414 1472 2414 0 ccff_head_0
rlabel metal1 20056 6222 20056 6222 0 ccff_tail
rlabel metal1 1794 49266 1794 49266 0 ccff_tail_0
rlabel metal2 25346 24871 25346 24871 0 chanx_right_in[0]
rlabel via2 25346 34187 25346 34187 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal1 25116 36142 25116 36142 0 chanx_right_in[12]
rlabel metal2 25346 36703 25346 36703 0 chanx_right_in[13]
rlabel metal2 25346 37349 25346 37349 0 chanx_right_in[14]
rlabel metal2 25346 38607 25346 38607 0 chanx_right_in[15]
rlabel metal1 24794 38930 24794 38930 0 chanx_right_in[16]
rlabel metal2 25346 40205 25346 40205 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25346 41565 25346 41565 0 chanx_right_in[19]
rlabel metal1 25438 24786 25438 24786 0 chanx_right_in[1]
rlabel metal1 24702 42534 24702 42534 0 chanx_right_in[20]
rlabel metal2 25346 43401 25346 43401 0 chanx_right_in[21]
rlabel metal2 25530 44353 25530 44353 0 chanx_right_in[22]
rlabel metal3 25952 44812 25952 44812 0 chanx_right_in[23]
rlabel metal1 24702 45798 24702 45798 0 chanx_right_in[24]
rlabel metal1 24840 46954 24840 46954 0 chanx_right_in[25]
rlabel metal2 25530 47889 25530 47889 0 chanx_right_in[26]
rlabel via2 25346 48093 25346 48093 0 chanx_right_in[27]
rlabel metal2 25346 49045 25346 49045 0 chanx_right_in[28]
rlabel metal2 25346 49759 25346 49759 0 chanx_right_in[29]
rlabel metal2 24150 28407 24150 28407 0 chanx_right_in[2]
rlabel metal1 24058 28492 24058 28492 0 chanx_right_in[3]
rlabel via2 25530 29291 25530 29291 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel metal2 25346 31127 25346 31127 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal2 25346 32725 25346 32725 0 chanx_right_in[8]
rlabel metal1 25392 32402 25392 32402 0 chanx_right_in[9]
rlabel metal3 25676 9724 25676 9724 0 chanx_right_out[10]
rlabel metal2 24610 9469 24610 9469 0 chanx_right_out[11]
rlabel metal2 24702 10421 24702 10421 0 chanx_right_out[12]
rlabel metal2 24794 11373 24794 11373 0 chanx_right_out[13]
rlabel metal3 25768 12988 25768 12988 0 chanx_right_out[14]
rlabel metal2 24794 13277 24794 13277 0 chanx_right_out[15]
rlabel metal2 25162 14297 25162 14297 0 chanx_right_out[16]
rlabel metal3 26228 15436 26228 15436 0 chanx_right_out[17]
rlabel metal2 24702 15589 24702 15589 0 chanx_right_out[18]
rlabel metal2 24794 16541 24794 16541 0 chanx_right_out[19]
rlabel metal3 24020 2380 24020 2380 0 chanx_right_out[1]
rlabel metal1 23368 18190 23368 18190 0 chanx_right_out[20]
rlabel metal2 24702 17901 24702 17901 0 chanx_right_out[21]
rlabel metal2 24794 18853 24794 18853 0 chanx_right_out[22]
rlabel metal1 24426 19890 24426 19890 0 chanx_right_out[23]
rlabel metal1 23368 20502 23368 20502 0 chanx_right_out[24]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[25]
rlabel metal3 24848 22780 24848 22780 0 chanx_right_out[26]
rlabel metal2 23874 23341 23874 23341 0 chanx_right_out[27]
rlabel metal1 24380 24242 24380 24242 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal3 24480 3196 24480 3196 0 chanx_right_out[2]
rlabel metal1 19274 5270 19274 5270 0 chanx_right_out[3]
rlabel metal3 24894 4828 24894 4828 0 chanx_right_out[4]
rlabel metal2 25162 4913 25162 4913 0 chanx_right_out[5]
rlabel metal3 25676 6460 25676 6460 0 chanx_right_out[6]
rlabel metal3 25584 7276 25584 7276 0 chanx_right_out[7]
rlabel metal3 25492 8092 25492 8092 0 chanx_right_out[8]
rlabel metal2 24702 8109 24702 8109 0 chanx_right_out[9]
rlabel metal2 1702 2098 1702 2098 0 chany_bottom_in[0]
rlabel metal1 5198 3026 5198 3026 0 chany_bottom_in[10]
rlabel metal1 5934 2346 5934 2346 0 chany_bottom_in[11]
rlabel metal2 6118 3706 6118 3706 0 chany_bottom_in[12]
rlabel metal2 6486 1761 6486 1761 0 chany_bottom_in[13]
rlabel metal2 6854 3196 6854 3196 0 chany_bottom_in[14]
rlabel metal2 7222 1588 7222 1588 0 chany_bottom_in[15]
rlabel metal1 7636 2414 7636 2414 0 chany_bottom_in[16]
rlabel metal2 7912 1972 7912 1972 0 chany_bottom_in[17]
rlabel metal1 7912 3026 7912 3026 0 chany_bottom_in[18]
rlabel metal1 8510 3026 8510 3026 0 chany_bottom_in[19]
rlabel metal1 1978 4522 1978 4522 0 chany_bottom_in[1]
rlabel metal2 9062 3502 9062 3502 0 chany_bottom_in[20]
rlabel metal2 9430 1761 9430 1761 0 chany_bottom_in[21]
rlabel metal1 9844 3502 9844 3502 0 chany_bottom_in[22]
rlabel metal1 9890 2414 9890 2414 0 chany_bottom_in[23]
rlabel metal2 10534 1761 10534 1761 0 chany_bottom_in[24]
rlabel metal1 10764 3502 10764 3502 0 chany_bottom_in[25]
rlabel metal2 11730 3196 11730 3196 0 chany_bottom_in[26]
rlabel metal1 11684 4046 11684 4046 0 chany_bottom_in[27]
rlabel metal1 11914 2448 11914 2448 0 chany_bottom_in[28]
rlabel metal1 10350 2380 10350 2380 0 chany_bottom_in[29]
rlabel metal2 2438 2438 2438 2438 0 chany_bottom_in[2]
rlabel metal2 2806 1761 2806 1761 0 chany_bottom_in[3]
rlabel metal2 3358 748 3358 748 0 chany_bottom_in[4]
rlabel metal1 1794 3536 1794 3536 0 chany_bottom_in[5]
rlabel metal1 3542 2414 3542 2414 0 chany_bottom_in[6]
rlabel metal1 4140 2414 4140 2414 0 chany_bottom_in[7]
rlabel metal1 4692 2414 4692 2414 0 chany_bottom_in[8]
rlabel metal1 4922 3366 4922 3366 0 chany_bottom_in[9]
rlabel metal2 12742 2166 12742 2166 0 chany_bottom_out[0]
rlabel metal2 16422 2404 16422 2404 0 chany_bottom_out[10]
rlabel metal2 16790 1792 16790 1792 0 chany_bottom_out[11]
rlabel metal2 17158 1826 17158 1826 0 chany_bottom_out[12]
rlabel metal2 17526 2404 17526 2404 0 chany_bottom_out[13]
rlabel metal2 17894 2166 17894 2166 0 chany_bottom_out[14]
rlabel metal2 18262 959 18262 959 0 chany_bottom_out[15]
rlabel metal2 18630 1792 18630 1792 0 chany_bottom_out[16]
rlabel metal2 18998 2098 18998 2098 0 chany_bottom_out[17]
rlabel metal2 19366 823 19366 823 0 chany_bottom_out[18]
rlabel metal2 19734 1826 19734 1826 0 chany_bottom_out[19]
rlabel metal2 13110 823 13110 823 0 chany_bottom_out[1]
rlabel metal2 20102 2404 20102 2404 0 chany_bottom_out[20]
rlabel metal2 20470 3254 20470 3254 0 chany_bottom_out[21]
rlabel metal2 20838 1826 20838 1826 0 chany_bottom_out[22]
rlabel metal2 21206 1775 21206 1775 0 chany_bottom_out[23]
rlabel metal2 21574 3254 21574 3254 0 chany_bottom_out[24]
rlabel metal2 21942 3492 21942 3492 0 chany_bottom_out[25]
rlabel metal1 22448 7310 22448 7310 0 chany_bottom_out[26]
rlabel metal2 22678 1792 22678 1792 0 chany_bottom_out[27]
rlabel metal2 23046 1639 23046 1639 0 chany_bottom_out[28]
rlabel metal2 23414 1860 23414 1860 0 chany_bottom_out[29]
rlabel metal2 13478 2404 13478 2404 0 chany_bottom_out[2]
rlabel metal2 13846 1554 13846 1554 0 chany_bottom_out[3]
rlabel metal2 14214 1860 14214 1860 0 chany_bottom_out[4]
rlabel metal2 14582 1622 14582 1622 0 chany_bottom_out[5]
rlabel metal2 14950 2166 14950 2166 0 chany_bottom_out[6]
rlabel metal2 15318 1622 15318 1622 0 chany_bottom_out[7]
rlabel metal2 15686 1860 15686 1860 0 chany_bottom_out[8]
rlabel metal2 16054 2166 16054 2166 0 chany_bottom_out[9]
rlabel metal1 11914 54196 11914 54196 0 chany_top_in_0[0]
rlabel metal1 16652 53550 16652 53550 0 chany_top_in_0[10]
rlabel metal1 17296 54162 17296 54162 0 chany_top_in_0[11]
rlabel metal1 17480 53550 17480 53550 0 chany_top_in_0[12]
rlabel metal1 18078 54230 18078 54230 0 chany_top_in_0[13]
rlabel metal2 18262 56236 18262 56236 0 chany_top_in_0[14]
rlabel metal1 19458 54128 19458 54128 0 chany_top_in_0[15]
rlabel metal1 18952 53074 18952 53074 0 chany_top_in_0[16]
rlabel metal1 19320 53550 19320 53550 0 chany_top_in_0[17]
rlabel metal1 19872 54162 19872 54162 0 chany_top_in_0[18]
rlabel metal1 20102 53550 20102 53550 0 chany_top_in_0[19]
rlabel metal2 13294 55711 13294 55711 0 chany_top_in_0[1]
rlabel metal1 20424 53074 20424 53074 0 chany_top_in_0[20]
rlabel metal2 20654 55711 20654 55711 0 chany_top_in_0[21]
rlabel metal1 21068 53550 21068 53550 0 chany_top_in_0[22]
rlabel metal1 21712 54162 21712 54162 0 chany_top_in_0[23]
rlabel metal1 21896 53550 21896 53550 0 chany_top_in_0[24]
rlabel metal1 22218 53210 22218 53210 0 chany_top_in_0[25]
rlabel metal1 22632 54162 22632 54162 0 chany_top_in_0[26]
rlabel metal1 23092 53550 23092 53550 0 chany_top_in_0[27]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[28]
rlabel metal1 23874 53074 23874 53074 0 chany_top_in_0[29]
rlabel metal1 13754 53142 13754 53142 0 chany_top_in_0[2]
rlabel metal1 14168 53550 14168 53550 0 chany_top_in_0[3]
rlabel metal1 14536 53074 14536 53074 0 chany_top_in_0[4]
rlabel metal1 14674 54298 14674 54298 0 chany_top_in_0[5]
rlabel metal1 15410 54162 15410 54162 0 chany_top_in_0[6]
rlabel metal1 15594 53550 15594 53550 0 chany_top_in_0[7]
rlabel metal1 16008 53074 16008 53074 0 chany_top_in_0[8]
rlabel metal1 16721 54162 16721 54162 0 chany_top_in_0[9]
rlabel metal1 2714 52938 2714 52938 0 chany_top_out_0[0]
rlabel metal1 5566 53652 5566 53652 0 chany_top_out_0[10]
rlabel metal1 4600 54094 4600 54094 0 chany_top_out_0[11]
rlabel metal1 6072 53142 6072 53142 0 chany_top_out_0[12]
rlabel metal1 6624 52462 6624 52462 0 chany_top_out_0[13]
rlabel metal1 7314 51442 7314 51442 0 chany_top_out_0[14]
rlabel metal1 6992 53618 6992 53618 0 chany_top_out_0[15]
rlabel metal2 7774 54376 7774 54376 0 chany_top_out_0[16]
rlabel metal2 7958 56236 7958 56236 0 chany_top_out_0[17]
rlabel metal2 8510 54070 8510 54070 0 chany_top_out_0[18]
rlabel metal1 8648 53618 8648 53618 0 chany_top_out_0[19]
rlabel metal1 2852 52666 2852 52666 0 chany_top_out_0[1]
rlabel metal1 9200 53142 9200 53142 0 chany_top_out_0[20]
rlabel metal2 9706 53550 9706 53550 0 chany_top_out_0[21]
rlabel metal1 9982 54264 9982 54264 0 chany_top_out_0[22]
rlabel metal2 10350 54614 10350 54614 0 chany_top_out_0[23]
rlabel metal1 10994 52530 10994 52530 0 chany_top_out_0[24]
rlabel metal2 11086 54920 11086 54920 0 chany_top_out_0[25]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[26]
rlabel metal1 12098 53006 12098 53006 0 chany_top_out_0[27]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[28]
rlabel metal1 12696 54094 12696 54094 0 chany_top_out_0[29]
rlabel metal2 2714 52972 2714 52972 0 chany_top_out_0[2]
rlabel metal2 2990 55711 2990 55711 0 chany_top_out_0[3]
rlabel metal2 3358 54070 3358 54070 0 chany_top_out_0[4]
rlabel metal1 3496 52530 3496 52530 0 chany_top_out_0[5]
rlabel metal2 4232 53244 4232 53244 0 chany_top_out_0[6]
rlabel metal1 4232 53142 4232 53142 0 chany_top_out_0[7]
rlabel metal2 4830 55711 4830 55711 0 chany_top_out_0[8]
rlabel metal1 5704 53210 5704 53210 0 chany_top_out_0[9]
rlabel metal1 20976 18734 20976 18734 0 clknet_0_prog_clk
rlabel metal1 8004 13362 8004 13362 0 clknet_4_0_0_prog_clk
rlabel metal1 6026 39474 6026 39474 0 clknet_4_10_0_prog_clk
rlabel metal1 12880 40018 12880 40018 0 clknet_4_11_0_prog_clk
rlabel metal1 19596 35122 19596 35122 0 clknet_4_12_0_prog_clk
rlabel metal1 22172 37230 22172 37230 0 clknet_4_13_0_prog_clk
rlabel metal2 19274 41854 19274 41854 0 clknet_4_14_0_prog_clk
rlabel metal1 22908 41038 22908 41038 0 clknet_4_15_0_prog_clk
rlabel metal2 11362 17340 11362 17340 0 clknet_4_1_0_prog_clk
rlabel metal1 9016 19890 9016 19890 0 clknet_4_2_0_prog_clk
rlabel metal1 10258 20978 10258 20978 0 clknet_4_3_0_prog_clk
rlabel metal1 18630 18190 18630 18190 0 clknet_4_4_0_prog_clk
rlabel metal1 18308 11866 18308 11866 0 clknet_4_5_0_prog_clk
rlabel metal2 15410 26180 15410 26180 0 clknet_4_6_0_prog_clk
rlabel metal1 22908 23698 22908 23698 0 clknet_4_7_0_prog_clk
rlabel metal1 6854 37162 6854 37162 0 clknet_4_8_0_prog_clk
rlabel metal1 12972 31246 12972 31246 0 clknet_4_9_0_prog_clk
rlabel metal3 1004 13804 1004 13804 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 16252 1004 16252 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18700 1004 18700 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 21148 1004 21148 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 1564 33490 1564 33490 0 gfpga_pad_io_soc_in[0]
rlabel metal1 1932 36142 1932 36142 0 gfpga_pad_io_soc_in[1]
rlabel metal1 1564 38318 1564 38318 0 gfpga_pad_io_soc_in[2]
rlabel metal1 1564 41106 1564 41106 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 23596 1004 23596 0 gfpga_pad_io_soc_out[0]
rlabel metal2 2806 26163 2806 26163 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 28492 1004 28492 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 30940 1004 30940 0 gfpga_pad_io_soc_out[3]
rlabel metal1 1518 43282 1518 43282 0 isol_n
rlabel metal1 2806 51034 2806 51034 0 net1
rlabel metal1 23299 39066 23299 39066 0 net10
rlabel metal3 23805 51068 23805 51068 0 net100
rlabel metal1 25116 38862 25116 38862 0 net101
rlabel metal2 22494 25738 22494 25738 0 net102
rlabel metal1 22494 40426 22494 40426 0 net103
rlabel metal2 23598 38403 23598 38403 0 net104
rlabel metal1 15870 14926 15870 14926 0 net105
rlabel metal1 22908 25874 22908 25874 0 net106
rlabel metal1 9614 40358 9614 40358 0 net107
rlabel metal1 14536 37366 14536 37366 0 net108
rlabel metal1 15686 40596 15686 40596 0 net109
rlabel metal1 20332 41242 20332 41242 0 net11
rlabel metal1 7682 52496 7682 52496 0 net110
rlabel metal1 18124 6290 18124 6290 0 net111
rlabel metal2 10994 37927 10994 37927 0 net112
rlabel metal1 22678 9996 22678 9996 0 net113
rlabel metal2 23966 9758 23966 9758 0 net114
rlabel metal1 23966 9588 23966 9588 0 net115
rlabel metal1 23920 10642 23920 10642 0 net116
rlabel metal2 22678 15164 22678 15164 0 net117
rlabel metal1 23644 12818 23644 12818 0 net118
rlabel metal2 22770 16048 22770 16048 0 net119
rlabel metal1 21298 41242 21298 41242 0 net12
rlabel metal1 23552 15470 23552 15470 0 net120
rlabel metal1 23828 14994 23828 14994 0 net121
rlabel metal2 24150 19040 24150 19040 0 net122
rlabel metal1 22862 5882 22862 5882 0 net123
rlabel metal2 22126 21148 22126 21148 0 net124
rlabel metal1 23644 25738 23644 25738 0 net125
rlabel metal2 23966 21692 23966 21692 0 net126
rlabel metal1 24978 27370 24978 27370 0 net127
rlabel metal1 24426 25126 24426 25126 0 net128
rlabel metal1 25300 25942 25300 25942 0 net129
rlabel metal1 22310 39576 22310 39576 0 net13
rlabel metal1 24564 26350 24564 26350 0 net130
rlabel metal2 23000 26860 23000 26860 0 net131
rlabel metal1 23046 24174 23046 24174 0 net132
rlabel metal1 23920 25874 23920 25874 0 net133
rlabel metal1 22310 8398 22310 8398 0 net134
rlabel metal1 20838 4794 20838 4794 0 net135
rlabel metal1 23184 7854 23184 7854 0 net136
rlabel metal2 24702 5372 24702 5372 0 net137
rlabel metal2 22770 7004 22770 7004 0 net138
rlabel metal1 24426 9894 24426 9894 0 net139
rlabel via2 25162 24667 25162 24667 0 net14
rlabel metal2 22218 5100 22218 5100 0 net140
rlabel metal1 23644 7378 23644 7378 0 net141
rlabel metal1 13018 15674 13018 15674 0 net142
rlabel metal1 16790 4114 16790 4114 0 net143
rlabel metal2 19458 6222 19458 6222 0 net144
rlabel metal1 18676 2618 18676 2618 0 net145
rlabel metal2 18814 4063 18814 4063 0 net146
rlabel metal1 19412 3502 19412 3502 0 net147
rlabel metal1 19826 2550 19826 2550 0 net148
rlabel metal1 19044 4590 19044 4590 0 net149
rlabel metal2 18354 40528 18354 40528 0 net15
rlabel metal1 21252 3502 21252 3502 0 net150
rlabel metal2 19550 6051 19550 6051 0 net151
rlabel metal1 21114 8330 21114 8330 0 net152
rlabel metal2 12650 3740 12650 3740 0 net153
rlabel metal2 22126 5507 22126 5507 0 net154
rlabel metal1 20470 5678 20470 5678 0 net155
rlabel metal1 21942 5202 21942 5202 0 net156
rlabel metal1 18400 9350 18400 9350 0 net157
rlabel metal1 21528 5678 21528 5678 0 net158
rlabel metal1 21712 6290 21712 6290 0 net159
rlabel metal3 24127 44268 24127 44268 0 net16
rlabel metal1 22080 7378 22080 7378 0 net160
rlabel metal1 20700 6290 20700 6290 0 net161
rlabel metal1 20562 7718 20562 7718 0 net162
rlabel metal1 19044 6630 19044 6630 0 net163
rlabel metal1 13616 4250 13616 4250 0 net164
rlabel metal1 12696 2414 12696 2414 0 net165
rlabel metal1 14122 12682 14122 12682 0 net166
rlabel metal2 14674 7548 14674 7548 0 net167
rlabel metal1 15364 3502 15364 3502 0 net168
rlabel metal2 16974 6188 16974 6188 0 net169
rlabel metal3 22724 36244 22724 36244 0 net17
rlabel metal1 16974 11526 16974 11526 0 net170
rlabel metal1 16606 3502 16606 3502 0 net171
rlabel metal2 1978 45526 1978 45526 0 net172
rlabel metal1 3082 53550 3082 53550 0 net173
rlabel metal1 2300 54162 2300 54162 0 net174
rlabel metal1 6348 44982 6348 44982 0 net175
rlabel metal1 5750 52462 5750 52462 0 net176
rlabel metal2 7130 51217 7130 51217 0 net177
rlabel metal1 6210 50490 6210 50490 0 net178
rlabel metal1 8372 45050 8372 45050 0 net179
rlabel metal1 24702 46478 24702 46478 0 net18
rlabel metal1 5106 54162 5106 54162 0 net180
rlabel metal1 8050 51918 8050 51918 0 net181
rlabel metal1 8234 53550 8234 53550 0 net182
rlabel metal1 2254 50218 2254 50218 0 net183
rlabel metal1 7636 53074 7636 53074 0 net184
rlabel metal1 10396 44506 10396 44506 0 net185
rlabel metal1 7406 54128 7406 54128 0 net186
rlabel metal1 9568 53074 9568 53074 0 net187
rlabel metal1 10212 52462 10212 52462 0 net188
rlabel metal1 11362 53550 11362 53550 0 net189
rlabel metal1 23598 45934 23598 45934 0 net19
rlabel metal1 10120 51578 10120 51578 0 net190
rlabel metal1 11822 52122 11822 52122 0 net191
rlabel metal2 12650 53108 12650 53108 0 net192
rlabel metal2 12374 53142 12374 53142 0 net193
rlabel metal1 2898 50830 2898 50830 0 net194
rlabel metal1 3082 51374 3082 51374 0 net195
rlabel metal1 2990 51884 2990 51884 0 net196
rlabel metal1 3726 52462 3726 52462 0 net197
rlabel metal1 4876 50898 4876 50898 0 net198
rlabel metal1 3588 53074 3588 53074 0 net199
rlabel metal2 2898 5814 2898 5814 0 net2
rlabel metal1 25392 47158 25392 47158 0 net20
rlabel metal2 7222 51646 7222 51646 0 net200
rlabel metal1 6118 51374 6118 51374 0 net201
rlabel metal2 1794 14892 1794 14892 0 net202
rlabel metal1 1794 19482 1794 19482 0 net203
rlabel metal2 1794 19754 1794 19754 0 net204
rlabel metal1 1840 21522 1840 21522 0 net205
rlabel metal1 1932 22746 1932 22746 0 net206
rlabel metal1 1932 26350 1932 26350 0 net207
rlabel metal1 1978 26010 1978 26010 0 net208
rlabel metal1 2024 28186 2024 28186 0 net209
rlabel metal2 22402 38420 22402 38420 0 net21
rlabel metal1 24472 2482 24472 2482 0 net210
rlabel metal2 17618 21182 17618 21182 0 net211
rlabel metal1 12926 28186 12926 28186 0 net212
rlabel metal2 21482 33728 21482 33728 0 net213
rlabel metal1 24978 23120 24978 23120 0 net214
rlabel metal1 14904 37842 14904 37842 0 net215
rlabel metal1 17158 21998 17158 21998 0 net216
rlabel metal2 20930 29376 20930 29376 0 net217
rlabel metal1 16928 36074 16928 36074 0 net218
rlabel metal1 17986 36890 17986 36890 0 net219
rlabel metal1 20516 36890 20516 36890 0 net22
rlabel metal1 17066 38862 17066 38862 0 net220
rlabel metal1 14674 39066 14674 39066 0 net221
rlabel metal1 13432 37230 13432 37230 0 net222
rlabel metal1 23460 39338 23460 39338 0 net223
rlabel metal1 12788 32402 12788 32402 0 net224
rlabel metal1 11270 30226 11270 30226 0 net225
rlabel metal1 13018 24242 13018 24242 0 net226
rlabel metal2 11822 25534 11822 25534 0 net227
rlabel metal2 9430 25602 9430 25602 0 net228
rlabel metal2 9154 26690 9154 26690 0 net229
rlabel metal1 18722 39610 18722 39610 0 net23
rlabel metal1 7958 24922 7958 24922 0 net230
rlabel metal1 10074 24820 10074 24820 0 net231
rlabel metal1 6394 9554 6394 9554 0 net232
rlabel metal2 14766 11458 14766 11458 0 net233
rlabel metal1 20608 32878 20608 32878 0 net234
rlabel metal2 17250 13056 17250 13056 0 net235
rlabel metal1 18768 15130 18768 15130 0 net236
rlabel metal2 20470 16830 20470 16830 0 net237
rlabel metal1 22356 15130 22356 15130 0 net238
rlabel metal1 20056 16082 20056 16082 0 net239
rlabel metal1 21114 41038 21114 41038 0 net24
rlabel metal1 21758 12206 21758 12206 0 net240
rlabel metal1 19596 10778 19596 10778 0 net241
rlabel metal1 19826 13260 19826 13260 0 net242
rlabel metal1 23046 34714 23046 34714 0 net243
rlabel metal2 22034 41344 22034 41344 0 net244
rlabel metal1 9936 37842 9936 37842 0 net245
rlabel metal1 7912 30770 7912 30770 0 net246
rlabel metal1 7406 32538 7406 32538 0 net247
rlabel metal1 13800 42194 13800 42194 0 net248
rlabel metal2 9798 33150 9798 33150 0 net249
rlabel metal2 23966 29546 23966 29546 0 net25
rlabel metal2 5382 32980 5382 32980 0 net250
rlabel metal1 8280 38318 8280 38318 0 net251
rlabel metal1 11270 37978 11270 37978 0 net252
rlabel metal1 10902 39066 10902 39066 0 net253
rlabel metal1 14582 35802 14582 35802 0 net254
rlabel metal1 9476 31450 9476 31450 0 net255
rlabel metal1 11316 23086 11316 23086 0 net256
rlabel metal1 12880 20434 12880 20434 0 net257
rlabel metal1 9568 16558 9568 16558 0 net258
rlabel metal1 9844 23766 9844 23766 0 net259
rlabel metal1 18124 26894 18124 26894 0 net26
rlabel metal2 13938 22100 13938 22100 0 net260
rlabel metal1 14076 24106 14076 24106 0 net261
rlabel metal1 20332 26962 20332 26962 0 net262
rlabel metal2 21666 25534 21666 25534 0 net263
rlabel metal2 17250 29716 17250 29716 0 net264
rlabel metal2 24610 2890 24610 2890 0 net265
rlabel metal1 22993 44778 22993 44778 0 net266
rlabel metal1 24334 3502 24334 3502 0 net267
rlabel metal1 25300 2618 25300 2618 0 net268
rlabel metal1 23828 8058 23828 8058 0 net269
rlabel metal1 25162 30804 25162 30804 0 net27
rlabel metal1 1978 52122 1978 52122 0 net270
rlabel metal1 4462 51238 4462 51238 0 net271
rlabel metal2 2254 3638 2254 3638 0 net272
rlabel metal1 4048 6426 4048 6426 0 net273
rlabel metal1 1610 52020 1610 52020 0 net274
rlabel metal2 1794 51884 1794 51884 0 net275
rlabel metal1 1932 2618 1932 2618 0 net276
rlabel metal1 2116 4250 2116 4250 0 net277
rlabel metal1 25162 29512 25162 29512 0 net28
rlabel metal2 23966 33456 23966 33456 0 net29
rlabel metal1 19826 24718 19826 24718 0 net3
rlabel metal1 20102 39066 20102 39066 0 net30
rlabel metal1 16238 37638 16238 37638 0 net31
rlabel metal1 17342 32402 17342 32402 0 net32
rlabel metal1 3772 3706 3772 3706 0 net33
rlabel metal1 7912 18938 7912 18938 0 net34
rlabel metal1 13202 36074 13202 36074 0 net35
rlabel metal1 16146 4046 16146 4046 0 net36
rlabel metal2 12466 38029 12466 38029 0 net37
rlabel metal1 7268 16966 7268 16966 0 net38
rlabel metal1 13064 17646 13064 17646 0 net39
rlabel metal1 13616 33626 13616 33626 0 net4
rlabel metal1 9890 2550 9890 2550 0 net40
rlabel via2 16698 36771 16698 36771 0 net41
rlabel via2 15778 36227 15778 36227 0 net42
rlabel metal2 18630 36669 18630 36669 0 net43
rlabel metal1 5934 18054 5934 18054 0 net44
rlabel metal1 14812 19686 14812 19686 0 net45
rlabel metal1 14950 20910 14950 20910 0 net46
rlabel metal2 13938 10409 13938 10409 0 net47
rlabel metal1 9844 2618 9844 2618 0 net48
rlabel metal1 15410 12206 15410 12206 0 net49
rlabel metal1 23598 30634 23598 30634 0 net5
rlabel metal1 15088 16626 15088 16626 0 net50
rlabel metal1 14076 19482 14076 19482 0 net51
rlabel metal2 15962 11050 15962 11050 0 net52
rlabel metal1 13570 2618 13570 2618 0 net53
rlabel metal1 11178 2482 11178 2482 0 net54
rlabel metal1 6118 20774 6118 20774 0 net55
rlabel metal2 2714 8058 2714 8058 0 net56
rlabel metal1 12650 13872 12650 13872 0 net57
rlabel metal2 1978 6035 1978 6035 0 net58
rlabel metal1 7176 25874 7176 25874 0 net59
rlabel metal3 21482 32300 21482 32300 0 net6
rlabel metal1 10442 33082 10442 33082 0 net60
rlabel metal1 5520 2414 5520 2414 0 net61
rlabel metal1 13386 36006 13386 36006 0 net62
rlabel metal1 12006 53958 12006 53958 0 net63
rlabel metal1 15318 12886 15318 12886 0 net64
rlabel metal1 16698 54026 16698 54026 0 net65
rlabel metal1 17940 47770 17940 47770 0 net66
rlabel metal1 18492 53958 18492 53958 0 net67
rlabel metal1 18492 53482 18492 53482 0 net68
rlabel metal1 19504 53958 19504 53958 0 net69
rlabel metal2 20102 36822 20102 36822 0 net7
rlabel metal1 18768 52870 18768 52870 0 net70
rlabel metal1 17158 18394 17158 18394 0 net71
rlabel metal1 20654 53958 20654 53958 0 net72
rlabel metal1 20562 53482 20562 53482 0 net73
rlabel metal1 13616 52462 13616 52462 0 net74
rlabel metal1 20286 52870 20286 52870 0 net75
rlabel metal1 21390 53958 21390 53958 0 net76
rlabel metal1 21436 53686 21436 53686 0 net77
rlabel metal2 22126 49827 22126 49827 0 net78
rlabel metal1 21620 53414 21620 53414 0 net79
rlabel metal1 25162 37128 25162 37128 0 net8
rlabel metal2 22494 50252 22494 50252 0 net80
rlabel metal1 20884 11798 20884 11798 0 net81
rlabel metal1 22448 43418 22448 43418 0 net82
rlabel metal1 22356 43826 22356 43826 0 net83
rlabel metal1 23092 46682 23092 46682 0 net84
rlabel via3 14053 52564 14053 52564 0 net85
rlabel metal3 14559 52564 14559 52564 0 net86
rlabel metal1 14628 52870 14628 52870 0 net87
rlabel metal1 13984 12410 13984 12410 0 net88
rlabel metal1 15502 53958 15502 53958 0 net89
rlabel metal1 23782 36686 23782 36686 0 net9
rlabel via3 16445 52564 16445 52564 0 net90
rlabel metal1 16606 47770 16606 47770 0 net91
rlabel via2 17526 11883 17526 11883 0 net92
rlabel metal1 2576 33286 2576 33286 0 net93
rlabel metal1 2898 36006 2898 36006 0 net94
rlabel metal2 1610 33932 1610 33932 0 net95
rlabel metal1 1656 40902 1656 40902 0 net96
rlabel metal2 8786 17340 8786 17340 0 net97
rlabel metal1 25116 3162 25116 3162 0 net98
rlabel metal1 23276 37910 23276 37910 0 net99
rlabel metal2 21390 17959 21390 17959 0 prog_clk
rlabel metal2 24150 1792 24150 1792 0 prog_reset
rlabel metal2 25070 50711 25070 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 25530 51561 25530 51561 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24794 52309 24794 52309 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 24978 53975 24978 53975 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 24932 53550 24932 53550 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25446 55420 25446 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel via2 4094 4029 4094 4029 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 20148 27302 20148 27302 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 18446 21862 18446 21862 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1211 11356 1211 11356 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18630 14042 18630 14042 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel via1 16054 22073 16054 22073 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 17250 18802 17250 18802 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 14398 21930 14398 21930 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal1 20562 21862 20562 21862 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 17388 25126 17388 25126 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal1 19550 34034 19550 34034 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal1 17480 26554 17480 26554 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal1 22310 26554 22310 26554 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 20608 34442 20608 34442 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal2 21206 29172 21206 29172 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal1 25162 24276 25162 24276 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal2 22678 32946 22678 32946 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal1 23000 25330 23000 25330 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 15548 30158 15548 30158 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 19366 36720 19366 36720 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 17664 32334 17664 32334 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal2 21666 20570 21666 20570 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 19872 27982 19872 27982 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 20102 20978 20102 20978 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal2 15548 32810 15548 32810 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 20378 35666 20378 35666 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 14674 33286 14674 33286 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 19504 33626 19504 33626 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal1 19872 34986 19872 34986 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal2 21666 33694 21666 33694 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 23966 21454 23966 21454 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 23690 22746 23690 22746 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 24196 23494 24196 23494 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 15916 37774 15916 37774 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 24334 23596 24334 23596 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 19218 22202 19218 22202 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal2 17710 36992 17710 36992 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 23690 29682 23690 29682 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal2 21620 32946 21620 32946 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 23644 30294 23644 30294 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 23736 44710 23736 44710 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal2 21206 43010 21206 43010 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 23230 45594 23230 45594 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 16606 36210 16606 36210 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal2 20102 44404 20102 44404 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal2 19826 44642 19826 44642 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal2 17342 38658 17342 38658 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal2 18630 45492 18630 45492 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 19366 46036 19366 46036 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 17664 37774 17664 37774 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 17112 40630 17112 40630 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal1 18538 46682 18538 46682 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 15364 39474 15364 39474 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 15594 40970 15594 40970 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal2 16330 45866 16330 45866 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal1 13984 41038 13984 41038 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 25254 43078 25254 43078 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 22770 41174 22770 41174 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 23460 41650 23460 41650 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 14168 34510 14168 34510 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel metal2 14674 39338 14674 39338 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal2 14030 37740 14030 37740 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal1 12811 29682 12811 29682 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 13524 35530 13524 35530 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 13570 34068 13570 34068 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 14352 26758 14352 26758 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal2 12834 27200 12834 27200 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal2 12926 27098 12926 27098 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal2 14490 27744 14490 27744 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 10672 27914 10672 27914 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal2 14858 27540 14858 27540 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 9108 28594 9108 28594 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 12742 29070 12742 29070 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 9016 26826 9016 26826 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 7912 27574 7912 27574 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal2 8602 24718 8602 24718 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 15502 29138 15502 29138 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal2 8786 12954 8786 12954 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 8142 23494 8142 23494 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 7728 18190 7728 18190 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 13616 11662 13616 11662 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal1 12926 13770 12926 13770 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 23414 34816 23414 34816 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 24288 42330 24288 42330 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 23230 38726 23230 38726 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal1 16146 13498 16146 13498 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal2 14858 14076 14858 14076 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal2 18630 16660 18630 16660 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 17158 16932 17158 16932 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal2 20194 17816 20194 17816 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal1 19274 18326 19274 18326 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 23230 17850 23230 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal1 21482 17850 21482 17850 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal2 21942 18054 21942 18054 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 22448 25806 22448 25806 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal1 21804 12274 21804 12274 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 21206 15436 21206 15436 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal2 20010 12070 20010 12070 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal1 19182 13362 19182 13362 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 18216 12410 18216 12410 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 24932 37774 24932 37774 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 22770 37774 22770 37774 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal2 23874 38148 23874 38148 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal1 23874 40154 23874 40154 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal2 22586 44642 22586 44642 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 12190 46444 12190 46444 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal1 15456 37298 15456 37298 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal1 12466 44268 12466 44268 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 7544 38386 7544 38386 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal2 6026 36244 6026 36244 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal1 7590 33966 7590 33966 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 9476 34034 9476 34034 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal1 7728 32334 7728 32334 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal1 14904 31790 14904 31790 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 8234 32946 8234 32946 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 13110 44914 13110 44914 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal2 19274 39219 19274 39219 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 14720 44506 14720 44506 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal2 9614 36125 9614 36125 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 18676 31790 18676 31790 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal1 9929 34374 9929 34374 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal2 5842 38522 5842 38522 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 13478 34612 13478 34612 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal2 7866 35904 7866 35904 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal1 10258 42092 10258 42092 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 7360 40562 7360 40562 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal1 8510 38318 8510 38318 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 10350 40902 10350 40902 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 19550 36210 19550 36210 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal1 14858 38420 14858 38420 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 12558 42568 12558 42568 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal2 16146 39780 16146 39780 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal1 18078 41038 18078 41038 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 15640 38386 15640 38386 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 18538 37978 18538 37978 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal2 8602 37944 8602 37944 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 19872 6766 19872 6766 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal1 15732 26010 15732 26010 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18400 32198 18400 32198 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13432 21590 13432 21590 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15226 24208 15226 24208 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13708 21658 13708 21658 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15180 17646 15180 17646 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 17342 9792 17342 9792 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 17434 28594 17434 28594 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19274 33830 19274 33830 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16882 25024 16882 25024 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14306 24650 14306 24650 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16928 24242 16928 24242 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16790 24820 16790 24820 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 17170 16882 17170 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 18860 9554 18860 9554 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal1 20102 29716 20102 29716 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 29614 20378 29614 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 27098 18814 27098 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20378 27744 20378 27744 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19918 26010 19918 26010 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18860 19822 18860 19822 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21206 8534 21206 8534 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 21988 29478 21988 29478 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21988 29614 21988 29614 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21114 26452 21114 26452 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24748 24174 24748 24174 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 24978 24752 24978 24752 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23506 24038 23506 24038 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16698 9622 16698 9622 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 16744 32538 16744 32538 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17250 34510 17250 34510 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17434 29274 17434 29274 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16928 32198 16928 32198 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 16054 28764 16054 28764 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15732 28390 15732 28390 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 20148 7854 20148 7854 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal1 19504 25330 19504 25330 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 25262 19642 25262 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19412 20570 19412 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19412 20434 19412 20434 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 17612 19826 17612 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14030 10030 14030 10030 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal1 17250 34646 17250 34646 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17894 34714 17894 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 34714 14904 34714 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13478 28730 13478 28730 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13340 21998 13340 21998 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17802 9894 17802 9894 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal2 21298 37468 21298 37468 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 31790 20378 31790 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20470 34102 20470 34102 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal3 19067 20604 19067 20604 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20930 7854 20930 7854 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal2 21666 27710 21666 27710 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22724 26282 22724 26282 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24242 23018 24242 23018 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22724 26486 22724 26486 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24058 22950 24058 22950 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 20838 18394 20838 18394 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9798 16422 9798 16422 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 13110 37128 13110 37128 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11776 37230 11776 37230 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10672 37230 10672 37230 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19136 8534 19136 8534 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 19458 26418 19458 26418 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20470 31926 20470 31926 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18308 24582 18308 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16882 21964 16882 21964 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19734 24582 19734 24582 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18722 21998 18722 21998 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19044 19414 19044 19414 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 22632 26962 22632 26962 0 sb_0__1_.mux_right_track_0.out
rlabel metal2 21390 32028 21390 32028 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21160 32742 21160 32742 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 30804 23414 30804 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23322 29240 23322 29240 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24794 28560 24794 28560 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22494 25738 22494 25738 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 20746 42160 20746 42160 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20240 40154 20240 40154 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 38386 20700 38386 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17572 36278 17572 36278 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22264 32402 22264 32402 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24702 27472 24702 27472 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 19826 45798 19826 45798 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19688 39474 19688 39474 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17066 36856 17066 36856 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19918 39270 19918 39270 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23138 25194 23138 25194 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 18584 41650 18584 41650 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18584 40154 18584 40154 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17618 37638 17618 37638 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22402 33609 22402 33609 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21528 28900 21528 28900 0 sb_0__1_.mux_right_track_16.out
rlabel metal2 17526 45424 17526 45424 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 40562 17112 40562 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14766 39270 14766 39270 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19780 32402 19780 32402 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21896 24174 21896 24174 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 16652 41650 16652 41650 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16422 37298 16422 37298 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14858 37162 14858 37162 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17434 37162 17434 37162 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24656 29206 24656 29206 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 23000 41650 23000 41650 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22218 40562 22218 40562 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21160 37706 21160 37706 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 25070 40596 25070 40596 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24978 39474 24978 39474 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24472 39270 24472 39270 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 21298 21760 21298 21760 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 13800 36890 13800 36890 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14628 32946 14628 32946 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 32640 14674 32640 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15686 33014 15686 33014 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21390 19822 21390 19822 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 13064 34034 13064 34034 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12926 33830 12926 33830 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10442 29818 10442 29818 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17802 24140 17802 24140 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21482 20808 21482 20808 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 15180 24786 15180 24786 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 24922 13938 24922 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17618 24650 17618 24650 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21206 18326 21206 18326 0 sb_0__1_.mux_right_track_26.out
rlabel metal1 15916 27098 15916 27098 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11500 25466 11500 25466 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18078 21522 18078 21522 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 19312 22494 19312 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 13478 26350 13478 26350 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12558 26078 12558 26078 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13938 21454 13938 21454 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19182 17136 19182 17136 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 10902 27506 10902 27506 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10672 26010 10672 26010 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16238 21454 16238 21454 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21160 16150 21160 16150 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 10672 25262 10672 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8050 24650 8050 24650 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14674 20434 14674 20434 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21850 15640 21850 15640 0 sb_0__1_.mux_right_track_34.out
rlabel metal2 12650 24412 12650 24412 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11178 24378 11178 24378 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13754 19550 13754 19550 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19826 10642 19826 10642 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 8142 24582 8142 24582 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8694 15504 8694 15504 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 12818 7590 12818 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14858 11696 14858 11696 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22218 10064 22218 10064 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 15364 11866 15364 11866 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15778 11084 15778 11084 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25070 27030 25070 27030 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 22218 38386 22218 38386 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22816 38250 22816 38250 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22770 36244 22770 36244 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 33320 22494 33320 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23092 30702 23092 30702 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23414 10676 23414 10676 0 sb_0__1_.mux_right_track_40.out
rlabel metal2 17342 14042 17342 14042 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 12614 20194 12614 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23736 9962 23736 9962 0 sb_0__1_.mux_right_track_44.out
rlabel metal2 18906 16456 18906 16456 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19918 12206 19918 12206 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24886 8976 24886 8976 0 sb_0__1_.mux_right_track_46.out
rlabel metal2 20562 17986 20562 17986 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20102 16456 20102 16456 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24518 6766 24518 6766 0 sb_0__1_.mux_right_track_48.out
rlabel metal2 20746 17680 20746 17680 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23414 12240 23414 12240 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23690 8942 23690 8942 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 21620 25670 21620 25670 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19596 16218 19596 16218 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 16660 21482 16660 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23414 4590 23414 4590 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 21068 12274 21068 12274 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22908 9554 22908 9554 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24012 4522 24012 4522 0 sb_0__1_.mux_right_track_54.out
rlabel metal1 19596 10642 19596 10642 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21206 8942 21206 8942 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23598 5678 23598 5678 0 sb_0__1_.mux_right_track_56.out
rlabel metal1 19642 13158 19642 13158 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21390 10030 21390 10030 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24610 26282 24610 26282 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 25024 38318 25024 38318 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24702 38080 24702 38080 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23690 34034 23690 34034 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23782 37196 23782 37196 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 23690 35943 23690 35943 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 23874 36278 23874 36278 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 24702 31416 24702 31416 0 sb_0__1_.mux_right_track_8.out
rlabel metal2 22034 44812 22034 44812 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 40698 21022 40698 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19964 37978 19964 37978 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22540 40562 22540 40562 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22954 40494 22954 40494 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 22586 40358 22586 40358 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12282 51986 12282 51986 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 10166 43146 10166 43146 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17158 42568 17158 42568 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12282 38131 12282 38131 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10304 37978 10304 37978 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11546 44506 11546 44506 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11408 45866 11408 45866 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10718 47668 10718 47668 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 7958 44506 7958 44506 0 sb_0__1_.mux_top_track_10.out
rlabel metal1 9430 38386 9430 38386 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17204 37366 17204 37366 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10810 33830 10810 33830 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8602 33898 8602 33898 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8234 36890 8234 36890 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9154 35462 9154 35462 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7866 44370 7866 44370 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7774 46614 7774 46614 0 sb_0__1_.mux_top_track_12.out
rlabel metal1 10856 33626 10856 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11638 32742 11638 32742 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7866 32810 7866 32810 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10396 33626 10396 33626 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 7498 34544 7498 34544 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7820 43282 7820 43282 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12788 48858 12788 48858 0 sb_0__1_.mux_top_track_2.out
rlabel metal1 16376 42330 16376 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18446 38522 18446 38522 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13064 36346 13064 36346 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15364 42330 15364 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13202 42330 13202 42330 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12926 45050 12926 45050 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8924 43962 8924 43962 0 sb_0__1_.mux_top_track_20.out
rlabel metal1 14030 35054 14030 35054 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15870 31450 15870 31450 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9706 32742 9706 32742 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 11086 36006 11086 36006 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9384 33082 9384 33082 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8832 43758 8832 43758 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5842 47396 5842 47396 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 10718 36142 10718 36142 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11270 34816 11270 34816 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9062 36346 9062 36346 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 5014 35190 5014 35190 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 5658 44370 5658 44370 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7360 46682 7360 46682 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 12282 38386 12282 38386 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11040 42262 11040 42262 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7728 38522 7728 38522 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9660 42330 9660 42330 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11408 51986 11408 51986 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 15088 38318 15088 38318 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19504 36346 19504 36346 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11040 33082 11040 33082 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14260 38522 14260 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10764 38522 10764 38522 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10902 41786 10902 41786 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 8004 52054 8004 52054 0 sb_0__1_.mux_top_track_44.out
rlabel metal2 15594 41208 15594 41208 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10810 38794 10810 38794 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11822 44982 11822 44982 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8878 46070 8878 46070 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 20240 38998 20240 38998 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17618 39066 17618 39066 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 36346 14904 36346 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14168 39542 14168 39542 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9844 51374 9844 51374 0 sb_0__1_.mux_top_track_6.out
rlabel metal2 10258 40052 10258 40052 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18032 38454 18032 38454 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 33456 14306 33456 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9200 34986 9200 34986 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8786 39610 8786 39610 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8372 35258 8372 35258 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7360 40154 7360 40154 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 1380 45594 1380 45594 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1518 48042 1518 48042 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 1334 50439 1334 50439 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 4002 52564 4002 52564 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
