magic
tech sky130A
magscale 1 2
timestamp 1656942999
<< obsli1 >>
rect 1104 2159 16008 17425
<< obsm1 >>
rect 290 1368 16914 17536
<< metal2 >>
rect 294 19200 350 20000
rect 662 19200 718 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11702 19200 11758 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14646 19200 14702 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16854 19200 16910 20000
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2870 0 2926 800
rect 3146 0 3202 800
rect 3422 0 3478 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
<< obsm2 >>
rect 406 19144 606 19258
rect 774 19144 974 19258
rect 1142 19144 1342 19258
rect 1510 19144 1710 19258
rect 1878 19144 2078 19258
rect 2246 19144 2446 19258
rect 2614 19144 2814 19258
rect 2982 19144 3182 19258
rect 3350 19144 3550 19258
rect 3718 19144 3918 19258
rect 4086 19144 4286 19258
rect 4454 19144 4654 19258
rect 4822 19144 5022 19258
rect 5190 19144 5390 19258
rect 5558 19144 5758 19258
rect 5926 19144 6126 19258
rect 6294 19144 6494 19258
rect 6662 19144 6862 19258
rect 7030 19144 7230 19258
rect 7398 19144 7598 19258
rect 7766 19144 7966 19258
rect 8134 19144 8334 19258
rect 8502 19144 8702 19258
rect 8870 19144 9070 19258
rect 9238 19144 9438 19258
rect 9606 19144 9806 19258
rect 9974 19144 10174 19258
rect 10342 19144 10542 19258
rect 10710 19144 10910 19258
rect 11078 19144 11278 19258
rect 11446 19144 11646 19258
rect 11814 19144 12014 19258
rect 12182 19144 12382 19258
rect 12550 19144 12750 19258
rect 12918 19144 13118 19258
rect 13286 19144 13486 19258
rect 13654 19144 13854 19258
rect 14022 19144 14222 19258
rect 14390 19144 14590 19258
rect 14758 19144 14958 19258
rect 15126 19144 15326 19258
rect 15494 19144 15694 19258
rect 15862 19144 16062 19258
rect 16230 19144 16430 19258
rect 16598 19144 16798 19258
rect 296 856 16908 19144
rect 296 800 1710 856
rect 1878 800 1986 856
rect 2154 800 2262 856
rect 2430 800 2538 856
rect 2706 800 2814 856
rect 2982 800 3090 856
rect 3258 800 3366 856
rect 3534 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4194 856
rect 4362 800 4470 856
rect 4638 800 4746 856
rect 4914 800 5022 856
rect 5190 800 5298 856
rect 5466 800 5574 856
rect 5742 800 5850 856
rect 6018 800 6126 856
rect 6294 800 6402 856
rect 6570 800 6678 856
rect 6846 800 6954 856
rect 7122 800 7230 856
rect 7398 800 7506 856
rect 7674 800 7782 856
rect 7950 800 8058 856
rect 8226 800 8334 856
rect 8502 800 8610 856
rect 8778 800 8886 856
rect 9054 800 9162 856
rect 9330 800 9438 856
rect 9606 800 9714 856
rect 9882 800 9990 856
rect 10158 800 10266 856
rect 10434 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11094 856
rect 11262 800 11370 856
rect 11538 800 11646 856
rect 11814 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12474 856
rect 12642 800 12750 856
rect 12918 800 13026 856
rect 13194 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13854 856
rect 14022 800 14130 856
rect 14298 800 14406 856
rect 14574 800 14682 856
rect 14850 800 14958 856
rect 15126 800 15234 856
rect 15402 800 16908 856
<< metal3 >>
rect 0 18912 800 19032
rect 0 17960 800 18080
rect 0 17008 800 17128
rect 16400 16600 17200 16720
rect 0 16056 800 16176
rect 0 15104 800 15224
rect 0 14152 800 14272
rect 0 13200 800 13320
rect 0 12248 800 12368
rect 0 11296 800 11416
rect 0 10344 800 10464
rect 16400 9936 17200 10056
rect 0 9392 800 9512
rect 0 8440 800 8560
rect 0 7488 800 7608
rect 0 6536 800 6656
rect 0 5584 800 5704
rect 0 4632 800 4752
rect 0 3680 800 3800
rect 16400 3272 17200 3392
rect 0 2728 800 2848
rect 0 1776 800 1896
rect 0 824 800 944
<< obsm3 >>
rect 880 18832 16400 19005
rect 800 18160 16400 18832
rect 880 17880 16400 18160
rect 800 17208 16400 17880
rect 880 16928 16400 17208
rect 800 16800 16400 16928
rect 800 16520 16320 16800
rect 800 16256 16400 16520
rect 880 15976 16400 16256
rect 800 15304 16400 15976
rect 880 15024 16400 15304
rect 800 14352 16400 15024
rect 880 14072 16400 14352
rect 800 13400 16400 14072
rect 880 13120 16400 13400
rect 800 12448 16400 13120
rect 880 12168 16400 12448
rect 800 11496 16400 12168
rect 880 11216 16400 11496
rect 800 10544 16400 11216
rect 880 10264 16400 10544
rect 800 10136 16400 10264
rect 800 9856 16320 10136
rect 800 9592 16400 9856
rect 880 9312 16400 9592
rect 800 8640 16400 9312
rect 880 8360 16400 8640
rect 800 7688 16400 8360
rect 880 7408 16400 7688
rect 800 6736 16400 7408
rect 880 6456 16400 6736
rect 800 5784 16400 6456
rect 880 5504 16400 5784
rect 800 4832 16400 5504
rect 880 4552 16400 4832
rect 800 3880 16400 4552
rect 880 3600 16400 3880
rect 800 3472 16400 3600
rect 800 3192 16320 3472
rect 800 2928 16400 3192
rect 880 2648 16400 2928
rect 800 1976 16400 2648
rect 880 1696 16400 1976
rect 800 1024 16400 1696
rect 880 851 16400 1024
<< metal4 >>
rect 2818 2128 3138 17456
rect 4692 2128 5012 17456
rect 6566 2128 6886 17456
rect 8440 2128 8760 17456
rect 10314 2128 10634 17456
rect 12188 2128 12508 17456
rect 14062 2128 14382 17456
<< obsm4 >>
rect 3371 2048 4612 17101
rect 5092 2048 6486 17101
rect 6966 2048 8360 17101
rect 8840 2048 10234 17101
rect 10714 2048 12108 17101
rect 12588 2048 13982 17101
rect 14462 2048 15029 17101
rect 3371 1803 15029 2048
<< labels >>
rlabel metal3 s 16400 16600 17200 16720 6 Test_en_E_in
port 1 nsew signal input
rlabel metal3 s 16400 9936 17200 10056 6 Test_en_E_out
port 2 nsew signal output
rlabel metal2 s 2134 19200 2190 20000 6 Test_en_N_out
port 3 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 Test_en_S_in
port 4 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 Test_en_W_in
port 5 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 Test_en_W_out
port 6 nsew signal output
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 7 nsew ground bidirectional
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 8 nsew power bidirectional
rlabel metal3 s 0 824 800 944 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 16400 3272 17200 3392 6 ccff_tail
port 10 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[0]
port 11 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[10]
port 12 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[11]
port 13 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[12]
port 14 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[13]
port 15 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[14]
port 16 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[15]
port 17 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_in[16]
port 18 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 chany_bottom_in[17]
port 19 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[18]
port 20 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_in[19]
port 21 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[1]
port 22 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[2]
port 23 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[3]
port 24 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_in[4]
port 25 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[5]
port 26 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[6]
port 27 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[7]
port 28 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[8]
port 29 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[9]
port 30 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[0]
port 31 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[10]
port 32 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[11]
port 33 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_out[12]
port 34 nsew signal output
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_out[13]
port 35 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_out[14]
port 36 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_out[15]
port 37 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[16]
port 38 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_out[17]
port 39 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_out[18]
port 40 nsew signal output
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[19]
port 41 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 chany_bottom_out[1]
port 42 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[2]
port 43 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 chany_bottom_out[3]
port 44 nsew signal output
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_out[4]
port 45 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[5]
port 46 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_out[6]
port 47 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_out[7]
port 48 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[8]
port 49 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_out[9]
port 50 nsew signal output
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[0]
port 51 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[10]
port 52 nsew signal input
rlabel metal2 s 13910 19200 13966 20000 6 chany_top_in[11]
port 53 nsew signal input
rlabel metal2 s 14278 19200 14334 20000 6 chany_top_in[12]
port 54 nsew signal input
rlabel metal2 s 14646 19200 14702 20000 6 chany_top_in[13]
port 55 nsew signal input
rlabel metal2 s 15014 19200 15070 20000 6 chany_top_in[14]
port 56 nsew signal input
rlabel metal2 s 15382 19200 15438 20000 6 chany_top_in[15]
port 57 nsew signal input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[16]
port 58 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[17]
port 59 nsew signal input
rlabel metal2 s 16486 19200 16542 20000 6 chany_top_in[18]
port 60 nsew signal input
rlabel metal2 s 16854 19200 16910 20000 6 chany_top_in[19]
port 61 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[1]
port 62 nsew signal input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[2]
port 63 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[3]
port 64 nsew signal input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[4]
port 65 nsew signal input
rlabel metal2 s 11702 19200 11758 20000 6 chany_top_in[5]
port 66 nsew signal input
rlabel metal2 s 12070 19200 12126 20000 6 chany_top_in[6]
port 67 nsew signal input
rlabel metal2 s 12438 19200 12494 20000 6 chany_top_in[7]
port 68 nsew signal input
rlabel metal2 s 12806 19200 12862 20000 6 chany_top_in[8]
port 69 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[9]
port 70 nsew signal input
rlabel metal2 s 2502 19200 2558 20000 6 chany_top_out[0]
port 71 nsew signal output
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[10]
port 72 nsew signal output
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[11]
port 73 nsew signal output
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[12]
port 74 nsew signal output
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[13]
port 75 nsew signal output
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[14]
port 76 nsew signal output
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[15]
port 77 nsew signal output
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[16]
port 78 nsew signal output
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_out[17]
port 79 nsew signal output
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_out[18]
port 80 nsew signal output
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_out[19]
port 81 nsew signal output
rlabel metal2 s 2870 19200 2926 20000 6 chany_top_out[1]
port 82 nsew signal output
rlabel metal2 s 3238 19200 3294 20000 6 chany_top_out[2]
port 83 nsew signal output
rlabel metal2 s 3606 19200 3662 20000 6 chany_top_out[3]
port 84 nsew signal output
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[4]
port 85 nsew signal output
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[5]
port 86 nsew signal output
rlabel metal2 s 4710 19200 4766 20000 6 chany_top_out[6]
port 87 nsew signal output
rlabel metal2 s 5078 19200 5134 20000 6 chany_top_out[7]
port 88 nsew signal output
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[8]
port 89 nsew signal output
rlabel metal2 s 5814 19200 5870 20000 6 chany_top_out[9]
port 90 nsew signal output
rlabel metal2 s 294 19200 350 20000 6 clk_2_N_out
port 91 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 clk_2_S_in
port 92 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 clk_2_S_out
port 93 nsew signal output
rlabel metal2 s 662 19200 718 20000 6 clk_3_N_out
port 94 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 clk_3_S_in
port 95 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 clk_3_S_out
port 96 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 left_grid_pin_16_
port 97 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 left_grid_pin_17_
port 98 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 left_grid_pin_18_
port 99 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 left_grid_pin_19_
port 100 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 left_grid_pin_20_
port 101 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 left_grid_pin_21_
port 102 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 left_grid_pin_22_
port 103 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 left_grid_pin_23_
port 104 nsew signal output
rlabel metal3 s 0 9392 800 9512 6 left_grid_pin_24_
port 105 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 left_grid_pin_25_
port 106 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 left_grid_pin_26_
port 107 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 left_grid_pin_27_
port 108 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 left_grid_pin_28_
port 109 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 left_grid_pin_29_
port 110 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 left_grid_pin_30_
port 111 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 left_grid_pin_31_
port 112 nsew signal output
rlabel metal2 s 1030 19200 1086 20000 6 prog_clk_0_N_out
port 113 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 prog_clk_0_S_out
port 114 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 prog_clk_0_W_in
port 115 nsew signal input
rlabel metal2 s 1398 19200 1454 20000 6 prog_clk_2_N_out
port 116 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 prog_clk_2_S_in
port 117 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 prog_clk_2_S_out
port 118 nsew signal output
rlabel metal2 s 1766 19200 1822 20000 6 prog_clk_3_N_out
port 119 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 prog_clk_3_S_in
port 120 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 prog_clk_3_S_out
port 121 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 17200 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1169466
string GDS_FILE /home/marwan/clear_signoff_final/openlane/cby_1__1_/runs/cby_1__1_/results/signoff/cby_1__1_.magic.gds
string GDS_START 65030
<< end >>

