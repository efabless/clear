magic
tech sky130A
magscale 1 2
timestamp 1625785166
<< locali >>
rect 8861 16507 8895 16677
rect 7205 14263 7239 14365
rect 10241 12835 10275 12937
rect 3341 10999 3375 11305
rect 9965 10999 9999 11237
rect 12541 10455 12575 10557
rect 8953 5763 8987 5865
rect 9873 5083 9907 5321
rect 5365 3451 5399 3621
<< viali >>
rect 2237 20553 2271 20587
rect 2605 20553 2639 20587
rect 4169 20553 4203 20587
rect 5089 20553 5123 20587
rect 8217 20553 8251 20587
rect 12909 20553 12943 20587
rect 19625 20553 19659 20587
rect 2881 20485 2915 20519
rect 3249 20485 3283 20519
rect 6285 20485 6319 20519
rect 8861 20485 8895 20519
rect 11621 20485 11655 20519
rect 12633 20485 12667 20519
rect 13093 20485 13127 20519
rect 13553 20485 13587 20519
rect 14013 20485 14047 20519
rect 14565 20485 14599 20519
rect 14933 20485 14967 20519
rect 15393 20485 15427 20519
rect 15853 20485 15887 20519
rect 16313 20485 16347 20519
rect 16773 20485 16807 20519
rect 17693 20485 17727 20519
rect 18153 20485 18187 20519
rect 18613 20485 18647 20519
rect 19073 20485 19107 20519
rect 19901 20485 19935 20519
rect 20269 20485 20303 20519
rect 20637 20485 20671 20519
rect 21005 20485 21039 20519
rect 5641 20417 5675 20451
rect 6193 20417 6227 20451
rect 7481 20417 7515 20451
rect 9781 20417 9815 20451
rect 17601 20417 17635 20451
rect 1501 20349 1535 20383
rect 4077 20349 4111 20383
rect 4537 20349 4571 20383
rect 4813 20349 4847 20383
rect 5549 20349 5583 20383
rect 6009 20349 6043 20383
rect 6653 20349 6687 20383
rect 8309 20349 8343 20383
rect 8677 20349 8711 20383
rect 9045 20349 9079 20383
rect 10241 20349 10275 20383
rect 10885 20349 10919 20383
rect 11437 20349 11471 20383
rect 12449 20349 12483 20383
rect 12817 20349 12851 20383
rect 14197 20349 14231 20383
rect 15117 20349 15151 20383
rect 21189 20349 21223 20383
rect 21557 20349 21591 20383
rect 1685 20281 1719 20315
rect 1961 20281 1995 20315
rect 2329 20281 2363 20315
rect 2697 20281 2731 20315
rect 3065 20281 3099 20315
rect 3433 20281 3467 20315
rect 3709 20281 3743 20315
rect 4997 20281 5031 20315
rect 7757 20281 7791 20315
rect 7941 20281 7975 20315
rect 9689 20281 9723 20315
rect 10609 20281 10643 20315
rect 11069 20281 11103 20315
rect 12081 20281 12115 20315
rect 13277 20281 13311 20315
rect 13737 20281 13771 20315
rect 14749 20281 14783 20315
rect 15577 20281 15611 20315
rect 16037 20281 16071 20315
rect 16497 20281 16531 20315
rect 16957 20281 16991 20315
rect 17417 20281 17451 20315
rect 17877 20281 17911 20315
rect 18337 20281 18371 20315
rect 18797 20281 18831 20315
rect 19257 20281 19291 20315
rect 19533 20281 19567 20315
rect 20085 20281 20119 20315
rect 20453 20281 20487 20315
rect 20821 20281 20855 20315
rect 1869 20213 1903 20247
rect 3893 20213 3927 20247
rect 4353 20213 4387 20247
rect 5457 20213 5491 20247
rect 6745 20213 6779 20247
rect 6929 20213 6963 20247
rect 7297 20213 7331 20247
rect 7389 20213 7423 20247
rect 8585 20213 8619 20247
rect 9229 20213 9263 20247
rect 9597 20213 9631 20247
rect 10149 20213 10183 20247
rect 10517 20213 10551 20247
rect 11345 20213 11379 20247
rect 11989 20213 12023 20247
rect 12357 20213 12391 20247
rect 21373 20213 21407 20247
rect 1869 20009 1903 20043
rect 2145 20009 2179 20043
rect 2605 20009 2639 20043
rect 3157 20009 3191 20043
rect 4353 20009 4387 20043
rect 6929 20009 6963 20043
rect 8861 20009 8895 20043
rect 13461 20009 13495 20043
rect 13645 20009 13679 20043
rect 16957 20009 16991 20043
rect 21557 20009 21591 20043
rect 1961 19941 1995 19975
rect 8585 19941 8619 19975
rect 10876 19941 10910 19975
rect 13829 19941 13863 19975
rect 17233 19941 17267 19975
rect 1593 19873 1627 19907
rect 2329 19873 2363 19907
rect 2421 19873 2455 19907
rect 2881 19873 2915 19907
rect 2973 19873 3007 19907
rect 3249 19873 3283 19907
rect 4261 19873 4295 19907
rect 4997 19873 5031 19907
rect 6213 19873 6247 19907
rect 6653 19873 6687 19907
rect 8042 19873 8076 19907
rect 10250 19873 10284 19907
rect 12081 19873 12115 19907
rect 12449 19873 12483 19907
rect 12909 19873 12943 19907
rect 13369 19873 13403 19907
rect 16773 19873 16807 19907
rect 17417 19873 17451 19907
rect 3525 19805 3559 19839
rect 4537 19805 4571 19839
rect 6469 19805 6503 19839
rect 8309 19805 8343 19839
rect 10517 19805 10551 19839
rect 10609 19805 10643 19839
rect 12725 19805 12759 19839
rect 1409 19737 1443 19771
rect 2697 19737 2731 19771
rect 3893 19737 3927 19771
rect 6837 19737 6871 19771
rect 8401 19737 8435 19771
rect 13185 19737 13219 19771
rect 3433 19669 3467 19703
rect 4813 19669 4847 19703
rect 5089 19669 5123 19703
rect 9137 19669 9171 19703
rect 11989 19669 12023 19703
rect 12265 19669 12299 19703
rect 12633 19669 12667 19703
rect 13093 19669 13127 19703
rect 14381 19669 14415 19703
rect 16589 19669 16623 19703
rect 1777 19465 1811 19499
rect 2053 19465 2087 19499
rect 3065 19465 3099 19499
rect 7113 19465 7147 19499
rect 9137 19465 9171 19499
rect 10609 19465 10643 19499
rect 13369 19465 13403 19499
rect 13645 19465 13679 19499
rect 13921 19465 13955 19499
rect 15301 19465 15335 19499
rect 15853 19465 15887 19499
rect 16497 19465 16531 19499
rect 18245 19465 18279 19499
rect 18521 19465 18555 19499
rect 19809 19465 19843 19499
rect 15025 19397 15059 19431
rect 19257 19397 19291 19431
rect 2513 19329 2547 19363
rect 7021 19329 7055 19363
rect 8493 19329 8527 19363
rect 9045 19329 9079 19363
rect 11437 19329 11471 19363
rect 1961 19261 1995 19295
rect 2237 19261 2271 19295
rect 2697 19261 2731 19295
rect 4270 19261 4304 19295
rect 4537 19261 4571 19295
rect 4629 19261 4663 19295
rect 6101 19261 6135 19295
rect 6745 19261 6779 19295
rect 8769 19261 8803 19295
rect 10517 19261 10551 19295
rect 11713 19261 11747 19295
rect 11980 19261 12014 19295
rect 13185 19261 13219 19295
rect 13461 19261 13495 19295
rect 13737 19261 13771 19295
rect 14013 19261 14047 19295
rect 14473 19261 14507 19295
rect 14841 19261 14875 19295
rect 15117 19261 15151 19295
rect 15393 19261 15427 19295
rect 15669 19261 15703 19295
rect 15945 19261 15979 19295
rect 16313 19261 16347 19295
rect 16589 19261 16623 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 18613 19261 18647 19295
rect 19073 19261 19107 19295
rect 19349 19261 19383 19295
rect 19625 19261 19659 19295
rect 1409 19193 1443 19227
rect 1593 19193 1627 19227
rect 4874 19193 4908 19227
rect 8248 19193 8282 19227
rect 10272 19193 10306 19227
rect 14381 19193 14415 19227
rect 17141 19193 17175 19227
rect 18981 19193 19015 19227
rect 2605 19125 2639 19159
rect 3157 19125 3191 19159
rect 6009 19125 6043 19159
rect 6561 19125 6595 19159
rect 8585 19125 8619 19159
rect 10793 19125 10827 19159
rect 11161 19125 11195 19159
rect 11253 19125 11287 19159
rect 13093 19125 13127 19159
rect 14197 19125 14231 19159
rect 14657 19125 14691 19159
rect 16129 19125 16163 19159
rect 16773 19125 16807 19159
rect 18797 19125 18831 19159
rect 1777 18921 1811 18955
rect 2053 18921 2087 18955
rect 2605 18921 2639 18955
rect 2881 18921 2915 18955
rect 6561 18921 6595 18955
rect 7021 18921 7055 18955
rect 7389 18921 7423 18955
rect 8217 18921 8251 18955
rect 8401 18921 8435 18955
rect 9321 18921 9355 18955
rect 10609 18921 10643 18955
rect 11069 18921 11103 18955
rect 11529 18921 11563 18955
rect 11713 18921 11747 18955
rect 12173 18921 12207 18955
rect 12541 18921 12575 18955
rect 13645 18921 13679 18955
rect 14197 18921 14231 18955
rect 15025 18921 15059 18955
rect 16865 18921 16899 18955
rect 18889 18921 18923 18955
rect 4261 18853 4295 18887
rect 6202 18853 6236 18887
rect 6929 18853 6963 18887
rect 8585 18853 8619 18887
rect 9781 18853 9815 18887
rect 12817 18853 12851 18887
rect 15577 18853 15611 18887
rect 1409 18785 1443 18819
rect 1593 18785 1627 18819
rect 1961 18785 1995 18819
rect 2237 18785 2271 18819
rect 2329 18785 2363 18819
rect 2789 18785 2823 18819
rect 3065 18785 3099 18819
rect 3157 18785 3191 18819
rect 3433 18785 3467 18819
rect 4721 18785 4755 18819
rect 7757 18785 7791 18819
rect 7849 18785 7883 18819
rect 9229 18785 9263 18819
rect 9689 18785 9723 18819
rect 10333 18785 10367 18819
rect 11161 18785 11195 18819
rect 12081 18785 12115 18819
rect 14013 18785 14047 18819
rect 14473 18785 14507 18819
rect 14565 18785 14599 18819
rect 14841 18785 14875 18819
rect 16681 18785 16715 18819
rect 18705 18785 18739 18819
rect 4353 18717 4387 18751
rect 4537 18717 4571 18751
rect 6469 18717 6503 18751
rect 7113 18717 7147 18751
rect 8033 18717 8067 18751
rect 9965 18717 9999 18751
rect 10517 18717 10551 18751
rect 10977 18717 11011 18751
rect 12357 18717 12391 18751
rect 2513 18649 2547 18683
rect 3341 18649 3375 18683
rect 3893 18649 3927 18683
rect 4905 18649 4939 18683
rect 10149 18649 10183 18683
rect 14749 18649 14783 18683
rect 3617 18581 3651 18615
rect 5089 18581 5123 18615
rect 16129 18581 16163 18615
rect 16405 18581 16439 18615
rect 17969 18581 18003 18615
rect 18429 18581 18463 18615
rect 1777 18377 1811 18411
rect 3985 18377 4019 18411
rect 4353 18377 4387 18411
rect 5273 18377 5307 18411
rect 5733 18377 5767 18411
rect 6469 18377 6503 18411
rect 7021 18377 7055 18411
rect 2513 18309 2547 18343
rect 5365 18309 5399 18343
rect 1409 18241 1443 18275
rect 4261 18241 4295 18275
rect 4813 18241 4847 18275
rect 4905 18241 4939 18275
rect 9413 18241 9447 18275
rect 11161 18241 11195 18275
rect 12265 18241 12299 18275
rect 1961 18173 1995 18207
rect 2053 18173 2087 18207
rect 2329 18173 2363 18207
rect 2605 18173 2639 18207
rect 2872 18173 2906 18207
rect 6009 18173 6043 18207
rect 1593 18105 1627 18139
rect 8769 18105 8803 18139
rect 9321 18105 9355 18139
rect 2237 18037 2271 18071
rect 4721 18037 4755 18071
rect 5549 18037 5583 18071
rect 6653 18037 6687 18071
rect 7297 18037 7331 18071
rect 8861 18037 8895 18071
rect 9229 18037 9263 18071
rect 11713 18037 11747 18071
rect 12081 18037 12115 18071
rect 12173 18037 12207 18071
rect 1501 17833 1535 17867
rect 1777 17833 1811 17867
rect 2329 17833 2363 17867
rect 2605 17833 2639 17867
rect 3157 17833 3191 17867
rect 3525 17833 3559 17867
rect 4445 17833 4479 17867
rect 4813 17833 4847 17867
rect 4997 17833 5031 17867
rect 8217 17833 8251 17867
rect 8585 17833 8619 17867
rect 9229 17833 9263 17867
rect 13185 17833 13219 17867
rect 13737 17833 13771 17867
rect 7205 17765 7239 17799
rect 1593 17697 1627 17731
rect 1961 17697 1995 17731
rect 2053 17697 2087 17731
rect 2513 17697 2547 17731
rect 2789 17697 2823 17731
rect 3065 17697 3099 17731
rect 3433 17697 3467 17731
rect 4353 17697 4387 17731
rect 7113 17697 7147 17731
rect 10037 17697 10071 17731
rect 12072 17697 12106 17731
rect 13553 17697 13587 17731
rect 4629 17629 4663 17663
rect 7297 17629 7331 17663
rect 7573 17629 7607 17663
rect 8677 17629 8711 17663
rect 8861 17629 8895 17663
rect 9781 17629 9815 17663
rect 11805 17629 11839 17663
rect 2237 17561 2271 17595
rect 2881 17561 2915 17595
rect 3985 17561 4019 17595
rect 6745 17561 6779 17595
rect 5273 17493 5307 17527
rect 11161 17493 11195 17527
rect 1869 17289 1903 17323
rect 2145 17289 2179 17323
rect 3341 17289 3375 17323
rect 4813 17289 4847 17323
rect 7849 17289 7883 17323
rect 9413 17289 9447 17323
rect 10977 17289 11011 17323
rect 13093 17289 13127 17323
rect 13369 17289 13403 17323
rect 9321 17221 9355 17255
rect 2421 17153 2455 17187
rect 2789 17153 2823 17187
rect 2881 17153 2915 17187
rect 11713 17153 11747 17187
rect 21557 17153 21591 17187
rect 2329 17085 2363 17119
rect 3433 17085 3467 17119
rect 3700 17085 3734 17119
rect 4905 17085 4939 17119
rect 5161 17085 5195 17119
rect 6469 17085 6503 17119
rect 7941 17085 7975 17119
rect 8197 17085 8231 17119
rect 10526 17085 10560 17119
rect 10793 17085 10827 17119
rect 11253 17085 11287 17119
rect 11980 17085 12014 17119
rect 13185 17085 13219 17119
rect 1593 17017 1627 17051
rect 1961 17017 1995 17051
rect 6736 17017 6770 17051
rect 21097 17017 21131 17051
rect 21373 17017 21407 17051
rect 1501 16949 1535 16983
rect 2973 16949 3007 16983
rect 6285 16949 6319 16983
rect 11069 16949 11103 16983
rect 11345 16949 11379 16983
rect 1961 16745 1995 16779
rect 2237 16745 2271 16779
rect 2329 16745 2363 16779
rect 3525 16745 3559 16779
rect 7389 16745 7423 16779
rect 7665 16745 7699 16779
rect 9781 16745 9815 16779
rect 10149 16745 10183 16779
rect 11069 16745 11103 16779
rect 11437 16745 11471 16779
rect 12265 16745 12299 16779
rect 12449 16745 12483 16779
rect 2513 16677 2547 16711
rect 3433 16677 3467 16711
rect 4445 16677 4479 16711
rect 8033 16677 8067 16711
rect 8861 16677 8895 16711
rect 11897 16677 11931 16711
rect 1593 16609 1627 16643
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 4353 16609 4387 16643
rect 5437 16609 5471 16643
rect 6929 16609 6963 16643
rect 7021 16609 7055 16643
rect 8125 16609 8159 16643
rect 4629 16541 4663 16575
rect 5181 16541 5215 16575
rect 6837 16541 6871 16575
rect 8217 16541 8251 16575
rect 9689 16609 9723 16643
rect 10241 16609 10275 16643
rect 12633 16609 12667 16643
rect 10425 16541 10459 16575
rect 10885 16541 10919 16575
rect 10977 16541 11011 16575
rect 11713 16541 11747 16575
rect 11805 16541 11839 16575
rect 6561 16473 6595 16507
rect 8585 16473 8619 16507
rect 8861 16473 8895 16507
rect 1501 16405 1535 16439
rect 3985 16405 4019 16439
rect 8769 16405 8803 16439
rect 1777 16201 1811 16235
rect 2145 16201 2179 16235
rect 5273 16201 5307 16235
rect 6745 16201 6779 16235
rect 7941 16201 7975 16235
rect 9045 16201 9079 16235
rect 11161 16201 11195 16235
rect 13461 16201 13495 16235
rect 8493 16065 8527 16099
rect 10425 16065 10459 16099
rect 11897 16065 11931 16099
rect 12909 16065 12943 16099
rect 1961 15997 1995 16031
rect 2329 15997 2363 16031
rect 3893 15997 3927 16031
rect 4160 15997 4194 16031
rect 6929 15997 6963 16031
rect 8401 15997 8435 16031
rect 11989 15997 12023 16031
rect 13093 15997 13127 16031
rect 1409 15929 1443 15963
rect 1593 15929 1627 15963
rect 8309 15929 8343 15963
rect 8861 15929 8895 15963
rect 12081 15929 12115 15963
rect 6469 15861 6503 15895
rect 10517 15861 10551 15895
rect 10609 15861 10643 15895
rect 10977 15861 11011 15895
rect 12449 15861 12483 15895
rect 13001 15861 13035 15895
rect 1777 15657 1811 15691
rect 2329 15657 2363 15691
rect 4721 15657 4755 15691
rect 8125 15657 8159 15691
rect 9321 15657 9355 15691
rect 9781 15657 9815 15691
rect 9873 15657 9907 15691
rect 10793 15657 10827 15691
rect 14105 15657 14139 15691
rect 4261 15589 4295 15623
rect 5181 15589 5215 15623
rect 6990 15589 7024 15623
rect 10701 15589 10735 15623
rect 11498 15589 11532 15623
rect 14626 15589 14660 15623
rect 1593 15521 1627 15555
rect 1961 15521 1995 15555
rect 2237 15521 2271 15555
rect 2513 15521 2547 15555
rect 4353 15521 4387 15555
rect 4813 15521 4847 15555
rect 6745 15521 6779 15555
rect 11253 15521 11287 15555
rect 12725 15521 12759 15555
rect 12992 15521 13026 15555
rect 4077 15453 4111 15487
rect 9689 15453 9723 15487
rect 10609 15453 10643 15487
rect 14381 15453 14415 15487
rect 1409 15385 1443 15419
rect 2053 15317 2087 15351
rect 8217 15317 8251 15351
rect 10241 15317 10275 15351
rect 11161 15317 11195 15351
rect 12633 15317 12667 15351
rect 15761 15317 15795 15351
rect 2053 15113 2087 15147
rect 2329 15113 2363 15147
rect 5549 15113 5583 15147
rect 6469 15113 6503 15147
rect 9781 15113 9815 15147
rect 11253 15113 11287 15147
rect 12449 15113 12483 15147
rect 13369 15113 13403 15147
rect 4261 15045 4295 15079
rect 1409 14977 1443 15011
rect 6193 14977 6227 15011
rect 8493 14977 8527 15011
rect 9229 14977 9263 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12633 14977 12667 15011
rect 13921 14977 13955 15011
rect 14473 14977 14507 15011
rect 2237 14909 2271 14943
rect 2513 14909 2547 14943
rect 2697 14909 2731 14943
rect 7849 14909 7883 14943
rect 8401 14909 8435 14943
rect 9321 14909 9355 14943
rect 9413 14909 9447 14943
rect 9873 14909 9907 14943
rect 12081 14909 12115 14943
rect 14565 14909 14599 14943
rect 15117 14909 15151 14943
rect 1593 14841 1627 14875
rect 2964 14841 2998 14875
rect 5917 14841 5951 14875
rect 7582 14841 7616 14875
rect 10140 14841 10174 14875
rect 12817 14841 12851 14875
rect 13829 14841 13863 14875
rect 4077 14773 4111 14807
rect 6009 14773 6043 14807
rect 7941 14773 7975 14807
rect 8309 14773 8343 14807
rect 12909 14773 12943 14807
rect 13277 14773 13311 14807
rect 13737 14773 13771 14807
rect 14657 14773 14691 14807
rect 15025 14773 15059 14807
rect 1777 14569 1811 14603
rect 2053 14569 2087 14603
rect 3249 14569 3283 14603
rect 7297 14569 7331 14603
rect 7757 14569 7791 14603
rect 8217 14569 8251 14603
rect 8677 14569 8711 14603
rect 9689 14569 9723 14603
rect 10425 14569 10459 14603
rect 10885 14569 10919 14603
rect 11437 14569 11471 14603
rect 13093 14569 13127 14603
rect 13461 14569 13495 14603
rect 4138 14501 4172 14535
rect 7113 14501 7147 14535
rect 12633 14501 12667 14535
rect 13921 14501 13955 14535
rect 14740 14501 14774 14535
rect 1409 14433 1443 14467
rect 1593 14433 1627 14467
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 3341 14433 3375 14467
rect 3893 14433 3927 14467
rect 5632 14433 5666 14467
rect 7665 14433 7699 14467
rect 8585 14433 8619 14467
rect 9321 14433 9355 14467
rect 10793 14433 10827 14467
rect 11253 14433 11287 14467
rect 13553 14433 13587 14467
rect 3065 14365 3099 14399
rect 5365 14365 5399 14399
rect 7205 14365 7239 14399
rect 7849 14365 7883 14399
rect 8769 14365 8803 14399
rect 11069 14365 11103 14399
rect 12357 14365 12391 14399
rect 12541 14365 12575 14399
rect 13645 14365 13679 14399
rect 14473 14365 14507 14399
rect 5273 14297 5307 14331
rect 9505 14297 9539 14331
rect 13001 14297 13035 14331
rect 2789 14229 2823 14263
rect 3709 14229 3743 14263
rect 6745 14229 6779 14263
rect 7205 14229 7239 14263
rect 9137 14229 9171 14263
rect 12173 14229 12207 14263
rect 15853 14229 15887 14263
rect 1501 14025 1535 14059
rect 2605 14025 2639 14059
rect 3157 14025 3191 14059
rect 11805 14025 11839 14059
rect 12633 14025 12667 14059
rect 12725 14025 12759 14059
rect 2053 13957 2087 13991
rect 2329 13957 2363 13991
rect 3065 13957 3099 13991
rect 4721 13957 4755 13991
rect 7849 13957 7883 13991
rect 3617 13889 3651 13923
rect 3801 13889 3835 13923
rect 5273 13889 5307 13923
rect 7021 13889 7055 13923
rect 9229 13889 9263 13923
rect 9781 13889 9815 13923
rect 9965 13889 9999 13923
rect 12081 13889 12115 13923
rect 13185 13889 13219 13923
rect 13369 13889 13403 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 1593 13821 1627 13855
rect 1961 13821 1995 13855
rect 2237 13821 2271 13855
rect 2513 13821 2547 13855
rect 2789 13821 2823 13855
rect 2881 13821 2915 13855
rect 3525 13821 3559 13855
rect 3985 13821 4019 13855
rect 5181 13821 5215 13855
rect 7113 13821 7147 13855
rect 7757 13821 7791 13855
rect 11529 13821 11563 13855
rect 13553 13821 13587 13855
rect 8984 13753 9018 13787
rect 9689 13753 9723 13787
rect 15025 13753 15059 13787
rect 1777 13685 1811 13719
rect 5089 13685 5123 13719
rect 7205 13685 7239 13719
rect 7573 13685 7607 13719
rect 9321 13685 9355 13719
rect 12173 13685 12207 13719
rect 12265 13685 12299 13719
rect 13093 13685 13127 13719
rect 13737 13685 13771 13719
rect 14657 13685 14691 13719
rect 1501 13481 1535 13515
rect 2421 13481 2455 13515
rect 2881 13481 2915 13515
rect 4537 13481 4571 13515
rect 6009 13481 6043 13515
rect 6837 13481 6871 13515
rect 7849 13481 7883 13515
rect 8217 13481 8251 13515
rect 8677 13481 8711 13515
rect 9597 13481 9631 13515
rect 12909 13481 12943 13515
rect 13277 13481 13311 13515
rect 13737 13481 13771 13515
rect 14841 13481 14875 13515
rect 15577 13481 15611 13515
rect 1593 13413 1627 13447
rect 7757 13413 7791 13447
rect 9505 13413 9539 13447
rect 15669 13413 15703 13447
rect 2329 13345 2363 13379
rect 3249 13345 3283 13379
rect 5650 13345 5684 13379
rect 5917 13345 5951 13379
rect 6377 13345 6411 13379
rect 7021 13345 7055 13379
rect 8585 13345 8619 13379
rect 9965 13345 9999 13379
rect 11437 13345 11471 13379
rect 11704 13345 11738 13379
rect 13369 13345 13403 13379
rect 14933 13345 14967 13379
rect 2513 13277 2547 13311
rect 3341 13277 3375 13311
rect 3433 13277 3467 13311
rect 6469 13277 6503 13311
rect 6561 13277 6595 13311
rect 7941 13277 7975 13311
rect 8769 13277 8803 13311
rect 9689 13277 9723 13311
rect 13553 13277 13587 13311
rect 14657 13277 14691 13311
rect 7205 13209 7239 13243
rect 10149 13209 10183 13243
rect 10241 13209 10275 13243
rect 12817 13209 12851 13243
rect 1777 13141 1811 13175
rect 1961 13141 1995 13175
rect 7389 13141 7423 13175
rect 9137 13141 9171 13175
rect 15301 13141 15335 13175
rect 1409 12937 1443 12971
rect 3525 12937 3559 12971
rect 4445 12937 4479 12971
rect 7849 12937 7883 12971
rect 10241 12937 10275 12971
rect 15853 12937 15887 12971
rect 16957 12869 16991 12903
rect 2789 12801 2823 12835
rect 4077 12801 4111 12835
rect 6469 12801 6503 12835
rect 9505 12801 9539 12835
rect 9689 12801 9723 12835
rect 10241 12801 10275 12835
rect 10517 12801 10551 12835
rect 12265 12801 12299 12835
rect 16405 12801 16439 12835
rect 2881 12733 2915 12767
rect 3157 12733 3191 12767
rect 3985 12733 4019 12767
rect 7941 12733 7975 12767
rect 8197 12733 8231 12767
rect 9781 12733 9815 12767
rect 12532 12733 12566 12767
rect 14381 12733 14415 12767
rect 18337 12733 18371 12767
rect 2544 12665 2578 12699
rect 6736 12665 6770 12699
rect 14648 12665 14682 12699
rect 18092 12665 18126 12699
rect 3065 12597 3099 12631
rect 3893 12597 3927 12631
rect 9321 12597 9355 12631
rect 10149 12597 10183 12631
rect 10609 12597 10643 12631
rect 10701 12597 10735 12631
rect 11069 12597 11103 12631
rect 13645 12597 13679 12631
rect 15761 12597 15795 12631
rect 16221 12597 16255 12631
rect 16313 12597 16347 12631
rect 1593 12393 1627 12427
rect 1869 12393 1903 12427
rect 2053 12393 2087 12427
rect 5549 12393 5583 12427
rect 7205 12393 7239 12427
rect 7665 12393 7699 12427
rect 8125 12393 8159 12427
rect 12265 12393 12299 12427
rect 12725 12393 12759 12427
rect 13093 12393 13127 12427
rect 14381 12393 14415 12427
rect 16313 12393 16347 12427
rect 4414 12325 4448 12359
rect 7573 12325 7607 12359
rect 9566 12325 9600 12359
rect 13553 12325 13587 12359
rect 1409 12257 1443 12291
rect 1685 12257 1719 12291
rect 3166 12257 3200 12291
rect 5641 12257 5675 12291
rect 5908 12257 5942 12291
rect 9321 12257 9355 12291
rect 10793 12257 10827 12291
rect 11049 12257 11083 12291
rect 12633 12257 12667 12291
rect 13461 12257 13495 12291
rect 15494 12257 15528 12291
rect 15761 12257 15795 12291
rect 16221 12257 16255 12291
rect 3433 12189 3467 12223
rect 4169 12189 4203 12223
rect 7757 12189 7791 12223
rect 12817 12189 12851 12223
rect 13645 12189 13679 12223
rect 16405 12189 16439 12223
rect 12173 12121 12207 12155
rect 3617 12053 3651 12087
rect 7021 12053 7055 12087
rect 10701 12053 10735 12087
rect 15853 12053 15887 12087
rect 2329 11849 2363 11883
rect 3617 11849 3651 11883
rect 5733 11849 5767 11883
rect 11253 11849 11287 11883
rect 12541 11849 12575 11883
rect 14933 11849 14967 11883
rect 1777 11713 1811 11747
rect 3065 11713 3099 11747
rect 4169 11713 4203 11747
rect 5181 11713 5215 11747
rect 7205 11713 7239 11747
rect 9137 11713 9171 11747
rect 9321 11713 9355 11747
rect 10701 11713 10735 11747
rect 11805 11713 11839 11747
rect 11989 11713 12023 11747
rect 13093 11713 13127 11747
rect 14381 11713 14415 11747
rect 16497 11713 16531 11747
rect 2881 11645 2915 11679
rect 9413 11645 9447 11679
rect 10793 11645 10827 11679
rect 16241 11645 16275 11679
rect 1869 11577 1903 11611
rect 2789 11577 2823 11611
rect 7472 11577 7506 11611
rect 10333 11577 10367 11611
rect 12081 11577 12115 11611
rect 13001 11577 13035 11611
rect 1409 11509 1443 11543
rect 1961 11509 1995 11543
rect 2421 11509 2455 11543
rect 3249 11509 3283 11543
rect 3985 11509 4019 11543
rect 4077 11509 4111 11543
rect 4537 11509 4571 11543
rect 5273 11509 5307 11543
rect 5365 11509 5399 11543
rect 6929 11509 6963 11543
rect 8585 11509 8619 11543
rect 9781 11509 9815 11543
rect 10885 11509 10919 11543
rect 12449 11509 12483 11543
rect 12909 11509 12943 11543
rect 14473 11509 14507 11543
rect 14565 11509 14599 11543
rect 15117 11509 15151 11543
rect 1869 11305 1903 11339
rect 2329 11305 2363 11339
rect 2697 11305 2731 11339
rect 3341 11305 3375 11339
rect 3985 11305 4019 11339
rect 5457 11305 5491 11339
rect 8493 11305 8527 11339
rect 9137 11305 9171 11339
rect 9597 11305 9631 11339
rect 14105 11305 14139 11339
rect 14473 11305 14507 11339
rect 1409 11169 1443 11203
rect 1685 11169 1719 11203
rect 2145 11101 2179 11135
rect 2789 11101 2823 11135
rect 2881 11101 2915 11135
rect 3157 11101 3191 11135
rect 1593 11033 1627 11067
rect 9965 11237 9999 11271
rect 11805 11237 11839 11271
rect 14933 11237 14967 11271
rect 5089 11169 5123 11203
rect 6828 11169 6862 11203
rect 8585 11169 8619 11203
rect 9505 11169 9539 11203
rect 3617 11101 3651 11135
rect 4905 11101 4939 11135
rect 4997 11101 5031 11135
rect 6561 11101 6595 11135
rect 8401 11101 8435 11135
rect 9689 11101 9723 11135
rect 3525 11033 3559 11067
rect 7941 11033 7975 11067
rect 8953 11033 8987 11067
rect 1961 10965 1995 10999
rect 3341 10965 3375 10999
rect 12173 11169 12207 11203
rect 12265 11169 12299 11203
rect 13093 11169 13127 11203
rect 14841 11169 14875 11203
rect 15301 11169 15335 11203
rect 10057 11101 10091 11135
rect 12081 11101 12115 11135
rect 13185 11101 13219 11135
rect 13277 11101 13311 11135
rect 15025 11101 15059 11135
rect 9965 10965 9999 10999
rect 12633 10965 12667 10999
rect 12725 10965 12759 10999
rect 1593 10761 1627 10795
rect 5089 10761 5123 10795
rect 8125 10761 8159 10795
rect 10517 10761 10551 10795
rect 14933 10761 14967 10795
rect 4077 10693 4111 10727
rect 4721 10625 4755 10659
rect 4905 10625 4939 10659
rect 5641 10625 5675 10659
rect 5917 10625 5951 10659
rect 6745 10625 6779 10659
rect 7573 10625 7607 10659
rect 11161 10625 11195 10659
rect 12449 10625 12483 10659
rect 14381 10625 14415 10659
rect 1409 10557 1443 10591
rect 1777 10557 1811 10591
rect 5549 10557 5583 10591
rect 6929 10557 6963 10591
rect 8401 10557 8435 10591
rect 8657 10557 8691 10591
rect 12541 10557 12575 10591
rect 12725 10557 12759 10591
rect 2044 10489 2078 10523
rect 6837 10489 6871 10523
rect 7757 10489 7791 10523
rect 10885 10489 10919 10523
rect 12970 10489 13004 10523
rect 3157 10421 3191 10455
rect 4261 10421 4295 10455
rect 4629 10421 4663 10455
rect 5457 10421 5491 10455
rect 7297 10421 7331 10455
rect 7665 10421 7699 10455
rect 9781 10421 9815 10455
rect 10333 10421 10367 10455
rect 10977 10421 11011 10455
rect 11805 10421 11839 10455
rect 12541 10421 12575 10455
rect 14105 10421 14139 10455
rect 14473 10421 14507 10455
rect 14565 10421 14599 10455
rect 1593 10217 1627 10251
rect 1869 10217 1903 10251
rect 2145 10217 2179 10251
rect 2329 10217 2363 10251
rect 3893 10217 3927 10251
rect 5365 10217 5399 10251
rect 7113 10217 7147 10251
rect 9413 10217 9447 10251
rect 9965 10217 9999 10251
rect 10425 10217 10459 10251
rect 14473 10217 14507 10251
rect 5006 10149 5040 10183
rect 10333 10149 10367 10183
rect 13185 10149 13219 10183
rect 15586 10149 15620 10183
rect 1409 10081 1443 10115
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 3453 10081 3487 10115
rect 5273 10081 5307 10115
rect 6745 10081 6779 10115
rect 7665 10081 7699 10115
rect 9505 10081 9539 10115
rect 11437 10081 11471 10115
rect 11693 10081 11727 10115
rect 13369 10081 13403 10115
rect 13829 10081 13863 10115
rect 13921 10081 13955 10115
rect 3709 10013 3743 10047
rect 6561 10013 6595 10047
rect 6653 10013 6687 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 9229 10013 9263 10047
rect 10517 10013 10551 10047
rect 14105 10013 14139 10047
rect 15853 10013 15887 10047
rect 7297 9877 7331 9911
rect 9873 9877 9907 9911
rect 12817 9877 12851 9911
rect 13461 9877 13495 9911
rect 1869 9605 1903 9639
rect 3985 9605 4019 9639
rect 4905 9605 4939 9639
rect 6837 9605 6871 9639
rect 11529 9605 11563 9639
rect 14565 9605 14599 9639
rect 2237 9537 2271 9571
rect 4537 9537 4571 9571
rect 5549 9537 5583 9571
rect 9321 9537 9355 9571
rect 10885 9537 10919 9571
rect 11069 9537 11103 9571
rect 11805 9537 11839 9571
rect 13093 9537 13127 9571
rect 13277 9537 13311 9571
rect 14013 9537 14047 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 1961 9469 1995 9503
rect 2421 9469 2455 9503
rect 2697 9469 2731 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 6193 9469 6227 9503
rect 8217 9469 8251 9503
rect 9237 9469 9271 9503
rect 13369 9469 13403 9503
rect 14197 9469 14231 9503
rect 2789 9401 2823 9435
rect 7950 9401 7984 9435
rect 9566 9401 9600 9435
rect 11989 9401 12023 9435
rect 12081 9401 12115 9435
rect 12541 9401 12575 9435
rect 1593 9333 1627 9367
rect 2145 9333 2179 9367
rect 2973 9333 3007 9367
rect 5273 9333 5307 9367
rect 5365 9333 5399 9367
rect 6009 9333 6043 9367
rect 9045 9333 9079 9367
rect 10701 9333 10735 9367
rect 11161 9333 11195 9367
rect 12449 9333 12483 9367
rect 13737 9333 13771 9367
rect 14105 9333 14139 9367
rect 1869 9129 1903 9163
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 4261 9129 4295 9163
rect 5733 9129 5767 9163
rect 7665 9129 7699 9163
rect 8125 9129 8159 9163
rect 11253 9129 11287 9163
rect 11713 9129 11747 9163
rect 12081 9129 12115 9163
rect 12173 9129 12207 9163
rect 12541 9129 12575 9163
rect 14657 9129 14691 9163
rect 6070 9061 6104 9095
rect 8769 9061 8803 9095
rect 10250 9061 10284 9095
rect 1409 8993 1443 9027
rect 1685 8993 1719 9027
rect 2237 8993 2271 9027
rect 3157 8993 3191 9027
rect 4620 8993 4654 9027
rect 8033 8993 8067 9027
rect 11345 8993 11379 9027
rect 13001 8993 13035 9027
rect 13645 8993 13679 9027
rect 2421 8925 2455 8959
rect 3249 8925 3283 8959
rect 3341 8925 3375 8959
rect 4353 8925 4387 8959
rect 5825 8925 5859 8959
rect 8217 8925 8251 8959
rect 8493 8925 8527 8959
rect 10517 8925 10551 8959
rect 11069 8925 11103 8959
rect 11989 8925 12023 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 14381 8925 14415 8959
rect 1593 8857 1627 8891
rect 7205 8857 7239 8891
rect 3709 8789 3743 8823
rect 9137 8789 9171 8823
rect 13185 8789 13219 8823
rect 14013 8789 14047 8823
rect 14933 8789 14967 8823
rect 1593 8585 1627 8619
rect 3525 8585 3559 8619
rect 5549 8585 5583 8619
rect 7849 8585 7883 8619
rect 8309 8585 8343 8619
rect 9137 8585 9171 8619
rect 9229 8585 9263 8619
rect 13645 8585 13679 8619
rect 6469 8517 6503 8551
rect 10701 8517 10735 8551
rect 11897 8517 11931 8551
rect 4077 8449 4111 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 6009 8449 6043 8483
rect 6101 8449 6135 8483
rect 7021 8449 7055 8483
rect 8585 8449 8619 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 11161 8449 11195 8483
rect 11253 8449 11287 8483
rect 12909 8449 12943 8483
rect 14197 8449 14231 8483
rect 15117 8449 15151 8483
rect 1409 8381 1443 8415
rect 2993 8381 3027 8415
rect 3249 8381 3283 8415
rect 8033 8381 8067 8415
rect 11713 8381 11747 8415
rect 13185 8381 13219 8415
rect 14013 8381 14047 8415
rect 14933 8381 14967 8415
rect 1685 8313 1719 8347
rect 3893 8313 3927 8347
rect 4629 8313 4663 8347
rect 5089 8313 5123 8347
rect 6837 8313 6871 8347
rect 7389 8313 7423 8347
rect 8769 8313 8803 8347
rect 10057 8313 10091 8347
rect 12725 8313 12759 8347
rect 13093 8313 13127 8347
rect 14105 8313 14139 8347
rect 15025 8313 15059 8347
rect 1869 8245 1903 8279
rect 3341 8245 3375 8279
rect 3985 8245 4019 8279
rect 5457 8245 5491 8279
rect 5917 8245 5951 8279
rect 6929 8245 6963 8279
rect 8677 8245 8711 8279
rect 9597 8245 9631 8279
rect 11069 8245 11103 8279
rect 13553 8245 13587 8279
rect 14565 8245 14599 8279
rect 1409 8041 1443 8075
rect 13921 8041 13955 8075
rect 2544 7973 2578 8007
rect 5580 7973 5614 8007
rect 7021 7973 7055 8007
rect 9689 7973 9723 8007
rect 10692 7973 10726 8007
rect 14626 7973 14660 8007
rect 2789 7905 2823 7939
rect 3249 7905 3283 7939
rect 3341 7905 3375 7939
rect 5825 7905 5859 7939
rect 6929 7905 6963 7939
rect 7757 7905 7791 7939
rect 9597 7905 9631 7939
rect 12541 7905 12575 7939
rect 12808 7905 12842 7939
rect 14381 7905 14415 7939
rect 16109 7905 16143 7939
rect 3433 7837 3467 7871
rect 4169 7837 4203 7871
rect 7205 7837 7239 7871
rect 7849 7837 7883 7871
rect 8033 7837 8067 7871
rect 9873 7837 9907 7871
rect 10425 7837 10459 7871
rect 15853 7837 15887 7871
rect 4445 7769 4479 7803
rect 6469 7769 6503 7803
rect 9229 7769 9263 7803
rect 2881 7701 2915 7735
rect 3893 7701 3927 7735
rect 4261 7701 4295 7735
rect 6561 7701 6595 7735
rect 7389 7701 7423 7735
rect 11805 7701 11839 7735
rect 15761 7701 15795 7735
rect 17233 7701 17267 7735
rect 1593 7497 1627 7531
rect 3525 7497 3559 7531
rect 4353 7497 4387 7531
rect 4629 7497 4663 7531
rect 6285 7497 6319 7531
rect 8953 7497 8987 7531
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 4077 7361 4111 7395
rect 5733 7361 5767 7395
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 9689 7361 9723 7395
rect 12173 7361 12207 7395
rect 14197 7361 14231 7395
rect 14381 7361 14415 7395
rect 15117 7361 15151 7395
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 1961 7293 1995 7327
rect 3893 7293 3927 7327
rect 3985 7293 4019 7327
rect 5917 7293 5951 7327
rect 6837 7293 6871 7327
rect 7573 7293 7607 7327
rect 9781 7293 9815 7327
rect 15301 7293 15335 7327
rect 2697 7225 2731 7259
rect 3157 7225 3191 7259
rect 4721 7225 4755 7259
rect 5825 7225 5859 7259
rect 7840 7225 7874 7259
rect 12357 7225 12391 7259
rect 14473 7225 14507 7259
rect 1869 7157 1903 7191
rect 2145 7157 2179 7191
rect 2329 7157 2363 7191
rect 4905 7157 4939 7191
rect 5181 7157 5215 7191
rect 5457 7157 5491 7191
rect 6469 7157 6503 7191
rect 6929 7157 6963 7191
rect 9873 7157 9907 7191
rect 10241 7157 10275 7191
rect 12265 7157 12299 7191
rect 12725 7157 12759 7191
rect 14841 7157 14875 7191
rect 15209 7157 15243 7191
rect 15669 7157 15703 7191
rect 2421 6953 2455 6987
rect 3341 6953 3375 6987
rect 5273 6953 5307 6987
rect 8309 6953 8343 6987
rect 10149 6953 10183 6987
rect 10885 6953 10919 6987
rect 14749 6953 14783 6987
rect 4261 6885 4295 6919
rect 6592 6885 6626 6919
rect 11998 6885 12032 6919
rect 1409 6817 1443 6851
rect 1685 6817 1719 6851
rect 2513 6817 2547 6851
rect 4353 6817 4387 6851
rect 4905 6817 4939 6851
rect 7196 6817 7230 6851
rect 9689 6817 9723 6851
rect 12357 6817 12391 6851
rect 14657 6817 14691 6851
rect 2605 6749 2639 6783
rect 3157 6749 3191 6783
rect 3249 6749 3283 6783
rect 4537 6749 4571 6783
rect 6837 6749 6871 6783
rect 6929 6749 6963 6783
rect 9413 6749 9447 6783
rect 9597 6749 9631 6783
rect 12265 6749 12299 6783
rect 14565 6749 14599 6783
rect 1593 6681 1627 6715
rect 1869 6681 1903 6715
rect 3893 6681 3927 6715
rect 5457 6681 5491 6715
rect 2053 6613 2087 6647
rect 3709 6613 3743 6647
rect 4721 6613 4755 6647
rect 5089 6613 5123 6647
rect 10057 6613 10091 6647
rect 12541 6613 12575 6647
rect 15117 6613 15151 6647
rect 1593 6409 1627 6443
rect 3249 6409 3283 6443
rect 7849 6409 7883 6443
rect 18337 6409 18371 6443
rect 5457 6341 5491 6375
rect 10517 6341 10551 6375
rect 12541 6341 12575 6375
rect 3985 6273 4019 6307
rect 4813 6273 4847 6307
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 6101 6273 6135 6307
rect 6561 6273 6595 6307
rect 7205 6273 7239 6307
rect 8401 6273 8435 6307
rect 10977 6273 11011 6307
rect 11069 6273 11103 6307
rect 11989 6273 12023 6307
rect 1409 6205 1443 6239
rect 1869 6205 1903 6239
rect 5733 6205 5767 6239
rect 6745 6205 6779 6239
rect 10425 6205 10459 6239
rect 10885 6205 10919 6239
rect 15209 6205 15243 6239
rect 16957 6205 16991 6239
rect 2114 6137 2148 6171
rect 4721 6137 4755 6171
rect 7297 6137 7331 6171
rect 8309 6137 8343 6171
rect 10180 6137 10214 6171
rect 12173 6137 12207 6171
rect 14942 6137 14976 6171
rect 17224 6137 17258 6171
rect 1685 6069 1719 6103
rect 3433 6069 3467 6103
rect 3801 6069 3835 6103
rect 3893 6069 3927 6103
rect 4353 6069 4387 6103
rect 5825 6069 5859 6103
rect 6929 6069 6963 6103
rect 7389 6069 7423 6103
rect 7757 6069 7791 6103
rect 8217 6069 8251 6103
rect 9045 6069 9079 6103
rect 12081 6069 12115 6103
rect 13829 6069 13863 6103
rect 15301 6069 15335 6103
rect 16773 6069 16807 6103
rect 1777 5865 1811 5899
rect 3893 5865 3927 5899
rect 4261 5865 4295 5899
rect 6101 5865 6135 5899
rect 6469 5865 6503 5899
rect 7941 5865 7975 5899
rect 8401 5865 8435 5899
rect 8953 5865 8987 5899
rect 9137 5865 9171 5899
rect 9321 5865 9355 5899
rect 10793 5865 10827 5899
rect 11161 5865 11195 5899
rect 11253 5865 11287 5899
rect 11897 5865 11931 5899
rect 14197 5865 14231 5899
rect 15117 5865 15151 5899
rect 15577 5865 15611 5899
rect 17877 5865 17911 5899
rect 21373 5865 21407 5899
rect 3617 5797 3651 5831
rect 4353 5797 4387 5831
rect 6285 5797 6319 5831
rect 7604 5797 7638 5831
rect 8309 5797 8343 5831
rect 8861 5797 8895 5831
rect 10456 5797 10490 5831
rect 11713 5797 11747 5831
rect 14749 5797 14783 5831
rect 15485 5797 15519 5831
rect 17969 5797 18003 5831
rect 1409 5729 1443 5763
rect 2901 5729 2935 5763
rect 3433 5729 3467 5763
rect 4988 5729 5022 5763
rect 8953 5729 8987 5763
rect 12633 5729 12667 5763
rect 12900 5729 12934 5763
rect 14657 5729 14691 5763
rect 16304 5729 16338 5763
rect 21281 5729 21315 5763
rect 21557 5729 21591 5763
rect 3157 5661 3191 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 7849 5661 7883 5695
rect 8493 5661 8527 5695
rect 10701 5661 10735 5695
rect 11345 5661 11379 5695
rect 14565 5661 14599 5695
rect 15301 5661 15335 5695
rect 16037 5661 16071 5695
rect 18061 5661 18095 5695
rect 1593 5593 1627 5627
rect 14013 5593 14047 5627
rect 17417 5593 17451 5627
rect 3341 5525 3375 5559
rect 15945 5525 15979 5559
rect 17509 5525 17543 5559
rect 4629 5321 4663 5355
rect 6469 5321 6503 5355
rect 7389 5321 7423 5355
rect 9873 5321 9907 5355
rect 1685 5253 1719 5287
rect 4077 5253 4111 5287
rect 7481 5253 7515 5287
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 5181 5185 5215 5219
rect 5549 5185 5583 5219
rect 6837 5185 6871 5219
rect 1501 5117 1535 5151
rect 1869 5117 1903 5151
rect 2136 5117 2170 5151
rect 3709 5117 3743 5151
rect 6101 5117 6135 5151
rect 8861 5117 8895 5151
rect 16773 5253 16807 5287
rect 10517 5185 10551 5219
rect 11345 5185 11379 5219
rect 12265 5185 12299 5219
rect 13093 5185 13127 5219
rect 14749 5185 14783 5219
rect 15393 5185 15427 5219
rect 17509 5185 17543 5219
rect 10333 5117 10367 5151
rect 12173 5117 12207 5151
rect 13360 5117 13394 5151
rect 17325 5117 17359 5151
rect 17785 5117 17819 5151
rect 19165 5117 19199 5151
rect 4353 5049 4387 5083
rect 4997 5049 5031 5083
rect 5089 5049 5123 5083
rect 5917 5049 5951 5083
rect 6929 5049 6963 5083
rect 8616 5049 8650 5083
rect 9045 5049 9079 5083
rect 9873 5049 9907 5083
rect 12081 5049 12115 5083
rect 14933 5049 14967 5083
rect 15638 5049 15672 5083
rect 3249 4981 3283 5015
rect 4169 4981 4203 5015
rect 5733 4981 5767 5015
rect 6193 4981 6227 5015
rect 7021 4981 7055 5015
rect 9965 4981 9999 5015
rect 10425 4981 10459 5015
rect 10793 4981 10827 5015
rect 11161 4981 11195 5015
rect 11253 4981 11287 5015
rect 11713 4981 11747 5015
rect 14473 4981 14507 5015
rect 14841 4981 14875 5015
rect 15301 4981 15335 5015
rect 16957 4981 16991 5015
rect 17417 4981 17451 5015
rect 17969 4981 18003 5015
rect 19349 4981 19383 5015
rect 2053 4777 2087 4811
rect 3065 4777 3099 4811
rect 3341 4777 3375 4811
rect 4537 4777 4571 4811
rect 6285 4777 6319 4811
rect 7021 4777 7055 4811
rect 7297 4777 7331 4811
rect 8217 4777 8251 4811
rect 8585 4777 8619 4811
rect 9965 4777 9999 4811
rect 10057 4777 10091 4811
rect 11253 4777 11287 4811
rect 12081 4777 12115 4811
rect 13277 4777 13311 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15117 4777 15151 4811
rect 15669 4777 15703 4811
rect 16773 4777 16807 4811
rect 17141 4777 17175 4811
rect 17233 4777 17267 4811
rect 1501 4709 1535 4743
rect 4353 4709 4387 4743
rect 7757 4709 7791 4743
rect 9137 4709 9171 4743
rect 12541 4709 12575 4743
rect 15577 4709 15611 4743
rect 16313 4709 16347 4743
rect 1777 4641 1811 4675
rect 2421 4641 2455 4675
rect 2873 4641 2907 4675
rect 3157 4641 3191 4675
rect 4077 4641 4111 4675
rect 5661 4641 5695 4675
rect 6193 4641 6227 4675
rect 6653 4641 6687 4675
rect 6929 4641 6963 4675
rect 7205 4641 7239 4675
rect 7665 4641 7699 4675
rect 8309 4641 8343 4675
rect 8677 4641 8711 4675
rect 9321 4641 9355 4675
rect 10609 4641 10643 4675
rect 11621 4641 11655 4675
rect 12449 4641 12483 4675
rect 13185 4641 13219 4675
rect 14749 4641 14783 4675
rect 16405 4641 16439 4675
rect 19993 4641 20027 4675
rect 1685 4573 1719 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 3617 4573 3651 4607
rect 5917 4573 5951 4607
rect 7849 4573 7883 4607
rect 9781 4573 9815 4607
rect 11713 4573 11747 4607
rect 11805 4573 11839 4607
rect 12725 4573 12759 4607
rect 13093 4573 13127 4607
rect 14473 4573 14507 4607
rect 14657 4573 14691 4607
rect 15761 4573 15795 4607
rect 16221 4573 16255 4607
rect 17049 4573 17083 4607
rect 1961 4505 1995 4539
rect 3893 4505 3927 4539
rect 9505 4505 9539 4539
rect 3433 4437 3467 4471
rect 4169 4437 4203 4471
rect 6009 4437 6043 4471
rect 6469 4437 6503 4471
rect 8953 4437 8987 4471
rect 10425 4437 10459 4471
rect 15209 4437 15243 4471
rect 17601 4437 17635 4471
rect 20177 4437 20211 4471
rect 3985 4233 4019 4267
rect 4445 4233 4479 4267
rect 6469 4233 6503 4267
rect 13645 4233 13679 4267
rect 3157 4165 3191 4199
rect 3709 4165 3743 4199
rect 1777 4097 1811 4131
rect 7021 4097 7055 4131
rect 7573 4097 7607 4131
rect 8493 4097 8527 4131
rect 9505 4097 9539 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 11437 4097 11471 4131
rect 11989 4097 12023 4131
rect 13277 4097 13311 4131
rect 15025 4097 15059 4131
rect 1501 4029 1535 4063
rect 3249 4029 3283 4063
rect 3525 4029 3559 4063
rect 3801 4029 3835 4063
rect 4077 4029 4111 4063
rect 5825 4029 5859 4063
rect 7297 4029 7331 4063
rect 7757 4029 7791 4063
rect 8677 4029 8711 4063
rect 12173 4029 12207 4063
rect 12817 4029 12851 4063
rect 13093 4029 13127 4063
rect 17141 4029 17175 4063
rect 2044 3961 2078 3995
rect 5558 3961 5592 3995
rect 6193 3961 6227 3995
rect 6929 3961 6963 3995
rect 8585 3961 8619 3995
rect 9689 3961 9723 3995
rect 10517 3961 10551 3995
rect 10977 3961 11011 3995
rect 14758 3961 14792 3995
rect 1593 3893 1627 3927
rect 3433 3893 3467 3927
rect 4261 3893 4295 3927
rect 5917 3893 5951 3927
rect 6837 3893 6871 3927
rect 7849 3893 7883 3927
rect 8217 3893 8251 3927
rect 9045 3893 9079 3927
rect 9137 3893 9171 3927
rect 9597 3893 9631 3927
rect 10057 3893 10091 3927
rect 10149 3893 10183 3927
rect 11253 3893 11287 3927
rect 12081 3893 12115 3927
rect 12541 3893 12575 3927
rect 12633 3893 12667 3927
rect 12909 3893 12943 3927
rect 15117 3893 15151 3927
rect 17325 3893 17359 3927
rect 1593 3689 1627 3723
rect 6193 3689 6227 3723
rect 6561 3689 6595 3723
rect 7021 3689 7055 3723
rect 7941 3689 7975 3723
rect 8769 3689 8803 3723
rect 9505 3689 9539 3723
rect 9873 3689 9907 3723
rect 12081 3689 12115 3723
rect 13369 3689 13403 3723
rect 14105 3689 14139 3723
rect 14381 3689 14415 3723
rect 15669 3689 15703 3723
rect 18337 3689 18371 3723
rect 2820 3621 2854 3655
rect 4160 3621 4194 3655
rect 5365 3621 5399 3655
rect 9413 3621 9447 3655
rect 14841 3621 14875 3655
rect 16037 3621 16071 3655
rect 1409 3553 1443 3587
rect 3249 3553 3283 3587
rect 3893 3553 3927 3587
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 5825 3553 5859 3587
rect 6653 3553 6687 3587
rect 7297 3553 7331 3587
rect 8677 3553 8711 3587
rect 10149 3553 10183 3587
rect 10405 3553 10439 3587
rect 11989 3553 12023 3587
rect 12449 3553 12483 3587
rect 12817 3553 12851 3587
rect 13093 3553 13127 3587
rect 13553 3553 13587 3587
rect 14749 3553 14783 3587
rect 15393 3553 15427 3587
rect 18061 3553 18095 3587
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6377 3485 6411 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 9321 3485 9355 3519
rect 12173 3485 12207 3519
rect 13829 3485 13863 3519
rect 14933 3485 14967 3519
rect 5273 3417 5307 3451
rect 5365 3417 5399 3451
rect 7113 3417 7147 3451
rect 11621 3417 11655 3451
rect 12633 3417 12667 3451
rect 15209 3417 15243 3451
rect 15577 3417 15611 3451
rect 18245 3417 18279 3451
rect 1685 3349 1719 3383
rect 3341 3349 3375 3383
rect 7573 3349 7607 3383
rect 8493 3349 8527 3383
rect 9965 3349 9999 3383
rect 11529 3349 11563 3383
rect 13001 3349 13035 3383
rect 13277 3349 13311 3383
rect 13645 3349 13679 3383
rect 15853 3349 15887 3383
rect 3525 3145 3559 3179
rect 5273 3145 5307 3179
rect 6193 3145 6227 3179
rect 7481 3145 7515 3179
rect 10333 3145 10367 3179
rect 10609 3145 10643 3179
rect 11897 3145 11931 3179
rect 13645 3145 13679 3179
rect 15761 3145 15795 3179
rect 21005 3145 21039 3179
rect 1685 3077 1719 3111
rect 4445 3077 4479 3111
rect 6469 3077 6503 3111
rect 14841 3077 14875 3111
rect 16037 3077 16071 3111
rect 16405 3077 16439 3111
rect 17325 3077 17359 3111
rect 18797 3077 18831 3111
rect 19625 3077 19659 3111
rect 20177 3077 20211 3111
rect 2605 3009 2639 3043
rect 2881 3009 2915 3043
rect 3801 3009 3835 3043
rect 4997 3009 5031 3043
rect 5641 3009 5675 3043
rect 5733 3009 5767 3043
rect 7113 3009 7147 3043
rect 8861 3009 8895 3043
rect 8953 3009 8987 3043
rect 11345 3009 11379 3043
rect 12265 3009 12299 3043
rect 1501 2941 1535 2975
rect 2329 2941 2363 2975
rect 3157 2941 3191 2975
rect 4813 2941 4847 2975
rect 5825 2941 5859 2975
rect 9220 2941 9254 2975
rect 10517 2941 10551 2975
rect 11161 2941 11195 2975
rect 12081 2941 12115 2975
rect 12521 2941 12555 2975
rect 13737 2941 13771 2975
rect 14013 2941 14047 2975
rect 14289 2941 14323 2975
rect 14657 2941 14691 2975
rect 14933 2941 14967 2975
rect 15301 2941 15335 2975
rect 15577 2941 15611 2975
rect 15853 2941 15887 2975
rect 16221 2941 16255 2975
rect 16497 2941 16531 2975
rect 16957 2941 16991 2975
rect 17141 2941 17175 2975
rect 17693 2941 17727 2975
rect 17877 2941 17911 2975
rect 18337 2941 18371 2975
rect 18613 2941 18647 2975
rect 19073 2941 19107 2975
rect 19441 2941 19475 2975
rect 19901 2941 19935 2975
rect 20361 2941 20395 2975
rect 20913 2941 20947 2975
rect 21189 2941 21223 2975
rect 4905 2873 4939 2907
rect 7297 2873 7331 2907
rect 8594 2873 8628 2907
rect 11805 2873 11839 2907
rect 17509 2873 17543 2907
rect 18429 2873 18463 2907
rect 21373 2873 21407 2907
rect 21557 2873 21591 2907
rect 1777 2805 1811 2839
rect 1961 2805 1995 2839
rect 2421 2805 2455 2839
rect 3065 2805 3099 2839
rect 3893 2805 3927 2839
rect 3985 2805 4019 2839
rect 4353 2805 4387 2839
rect 6837 2805 6871 2839
rect 6929 2805 6963 2839
rect 10793 2805 10827 2839
rect 11253 2805 11287 2839
rect 13921 2805 13955 2839
rect 14197 2805 14231 2839
rect 14473 2805 14507 2839
rect 15117 2805 15151 2839
rect 15485 2805 15519 2839
rect 16681 2805 16715 2839
rect 18061 2805 18095 2839
rect 18153 2805 18187 2839
rect 18889 2805 18923 2839
rect 19257 2805 19291 2839
rect 19717 2805 19751 2839
rect 20545 2805 20579 2839
rect 1777 2601 1811 2635
rect 2237 2601 2271 2635
rect 2605 2601 2639 2635
rect 3985 2601 4019 2635
rect 4629 2601 4663 2635
rect 4997 2601 5031 2635
rect 5273 2601 5307 2635
rect 5917 2601 5951 2635
rect 6285 2601 6319 2635
rect 7481 2601 7515 2635
rect 7573 2601 7607 2635
rect 8033 2601 8067 2635
rect 8493 2601 8527 2635
rect 9229 2601 9263 2635
rect 9781 2601 9815 2635
rect 10333 2601 10367 2635
rect 10793 2601 10827 2635
rect 11253 2601 11287 2635
rect 12265 2601 12299 2635
rect 12633 2601 12667 2635
rect 13185 2601 13219 2635
rect 14381 2601 14415 2635
rect 17049 2601 17083 2635
rect 1685 2533 1719 2567
rect 2697 2533 2731 2567
rect 3433 2533 3467 2567
rect 4721 2533 4755 2567
rect 5825 2533 5859 2567
rect 6837 2533 6871 2567
rect 8401 2533 8435 2567
rect 10701 2533 10735 2567
rect 13645 2533 13679 2567
rect 14013 2533 14047 2567
rect 14749 2533 14783 2567
rect 15485 2533 15519 2567
rect 16313 2533 16347 2567
rect 16773 2533 16807 2567
rect 17417 2533 17451 2567
rect 17693 2533 17727 2567
rect 18613 2533 18647 2567
rect 19165 2533 19199 2567
rect 19625 2533 19659 2567
rect 20545 2533 20579 2567
rect 21465 2533 21499 2567
rect 3249 2465 3283 2499
rect 3617 2465 3651 2499
rect 4077 2465 4111 2499
rect 4261 2465 4295 2499
rect 5089 2465 5123 2499
rect 5457 2465 5491 2499
rect 6653 2465 6687 2499
rect 6929 2465 6963 2499
rect 9045 2465 9079 2499
rect 9413 2465 9447 2499
rect 9873 2465 9907 2499
rect 11345 2465 11379 2499
rect 11713 2465 11747 2499
rect 12909 2465 12943 2499
rect 13277 2465 13311 2499
rect 14197 2465 14231 2499
rect 15117 2465 15151 2499
rect 15853 2465 15887 2499
rect 18153 2465 18187 2499
rect 20085 2465 20119 2499
rect 21005 2465 21039 2499
rect 1593 2397 1627 2431
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 5641 2397 5675 2431
rect 7389 2397 7423 2431
rect 8677 2397 8711 2431
rect 9689 2397 9723 2431
rect 10885 2397 10919 2431
rect 12081 2397 12115 2431
rect 12173 2397 12207 2431
rect 17877 2397 17911 2431
rect 2145 2329 2179 2363
rect 7941 2329 7975 2363
rect 10241 2329 10275 2363
rect 13461 2329 13495 2363
rect 13829 2329 13863 2363
rect 14565 2329 14599 2363
rect 14933 2329 14967 2363
rect 15301 2329 15335 2363
rect 15669 2329 15703 2363
rect 16129 2329 16163 2363
rect 16589 2329 16623 2363
rect 17233 2329 17267 2363
rect 17969 2329 18003 2363
rect 18981 2329 19015 2363
rect 19441 2329 19475 2363
rect 19901 2329 19935 2363
rect 20361 2329 20395 2363
rect 20821 2329 20855 2363
rect 21281 2329 21315 2363
rect 4445 2261 4479 2295
rect 7113 2261 7147 2295
rect 8861 2261 8895 2295
rect 11529 2261 11563 2295
rect 12817 2261 12851 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2774 20584 2780 20596
rect 2639 20556 2780 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 3878 20544 3884 20596
rect 3936 20584 3942 20596
rect 4062 20584 4068 20596
rect 3936 20556 4068 20584
rect 3936 20544 3942 20556
rect 4062 20544 4068 20556
rect 4120 20584 4126 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 4120 20556 4169 20584
rect 4120 20544 4126 20556
rect 4157 20553 4169 20556
rect 4203 20553 4215 20587
rect 5077 20587 5135 20593
rect 5077 20584 5089 20587
rect 4157 20547 4215 20553
rect 4264 20556 5089 20584
rect 2866 20516 2872 20528
rect 2827 20488 2872 20516
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 3234 20516 3240 20528
rect 3195 20488 3240 20516
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 3510 20476 3516 20528
rect 3568 20516 3574 20528
rect 4264 20516 4292 20556
rect 5077 20553 5089 20556
rect 5123 20553 5135 20587
rect 5077 20547 5135 20553
rect 5166 20544 5172 20596
rect 5224 20584 5230 20596
rect 5224 20556 6408 20584
rect 5224 20544 5230 20556
rect 3568 20488 4292 20516
rect 3568 20476 3574 20488
rect 4338 20476 4344 20528
rect 4396 20516 4402 20528
rect 6273 20519 6331 20525
rect 6273 20516 6285 20519
rect 4396 20488 6285 20516
rect 4396 20476 4402 20488
rect 6273 20485 6285 20488
rect 6319 20485 6331 20519
rect 6273 20479 6331 20485
rect 1118 20408 1124 20460
rect 1176 20448 1182 20460
rect 3694 20448 3700 20460
rect 1176 20420 3700 20448
rect 1176 20408 1182 20420
rect 3694 20408 3700 20420
rect 3752 20408 3758 20460
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20448 5687 20451
rect 5810 20448 5816 20460
rect 5675 20420 5816 20448
rect 5675 20417 5687 20420
rect 5629 20411 5687 20417
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6181 20451 6239 20457
rect 6181 20448 6193 20451
rect 6144 20420 6193 20448
rect 6144 20408 6150 20420
rect 6181 20417 6193 20420
rect 6227 20417 6239 20451
rect 6380 20448 6408 20556
rect 7190 20544 7196 20596
rect 7248 20584 7254 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7248 20556 8217 20584
rect 7248 20544 7254 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 10134 20584 10140 20596
rect 8205 20547 8263 20553
rect 8956 20556 10140 20584
rect 6454 20476 6460 20528
rect 6512 20516 6518 20528
rect 8849 20519 8907 20525
rect 8849 20516 8861 20519
rect 6512 20488 8861 20516
rect 6512 20476 6518 20488
rect 8849 20485 8861 20488
rect 8895 20485 8907 20519
rect 8849 20479 8907 20485
rect 7466 20448 7472 20460
rect 6380 20420 7328 20448
rect 7427 20420 7472 20448
rect 6181 20411 6239 20417
rect 198 20340 204 20392
rect 256 20380 262 20392
rect 1489 20383 1547 20389
rect 1489 20380 1501 20383
rect 256 20352 1501 20380
rect 256 20340 262 20352
rect 1489 20349 1501 20352
rect 1535 20380 1547 20383
rect 1578 20380 1584 20392
rect 1535 20352 1584 20380
rect 1535 20349 1547 20352
rect 1489 20343 1547 20349
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 4062 20340 4068 20392
rect 4120 20380 4126 20392
rect 4120 20352 4165 20380
rect 4120 20340 4126 20352
rect 4338 20340 4344 20392
rect 4396 20380 4402 20392
rect 4525 20383 4583 20389
rect 4525 20380 4537 20383
rect 4396 20352 4537 20380
rect 4396 20340 4402 20352
rect 4525 20349 4537 20352
rect 4571 20349 4583 20383
rect 4798 20380 4804 20392
rect 4759 20352 4804 20380
rect 4525 20343 4583 20349
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 5534 20380 5540 20392
rect 5495 20352 5540 20380
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 5997 20383 6055 20389
rect 5997 20380 6009 20383
rect 5776 20352 6009 20380
rect 5776 20340 5782 20352
rect 5997 20349 6009 20352
rect 6043 20349 6055 20383
rect 5997 20343 6055 20349
rect 6270 20340 6276 20392
rect 6328 20380 6334 20392
rect 6641 20383 6699 20389
rect 6641 20380 6653 20383
rect 6328 20352 6653 20380
rect 6328 20340 6334 20352
rect 6641 20349 6653 20352
rect 6687 20349 6699 20383
rect 6641 20343 6699 20349
rect 6914 20340 6920 20392
rect 6972 20340 6978 20392
rect 7300 20380 7328 20420
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 8956 20448 8984 20556
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 10594 20544 10600 20596
rect 10652 20584 10658 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 10652 20556 12909 20584
rect 10652 20544 10658 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 19613 20587 19671 20593
rect 19613 20553 19625 20587
rect 19659 20584 19671 20587
rect 21358 20584 21364 20596
rect 19659 20556 21364 20584
rect 19659 20553 19671 20556
rect 19613 20547 19671 20553
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 11609 20519 11667 20525
rect 11609 20516 11621 20519
rect 7576 20420 8984 20448
rect 9048 20488 11621 20516
rect 7576 20380 7604 20420
rect 7300 20352 7604 20380
rect 7650 20340 7656 20392
rect 7708 20380 7714 20392
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 7708 20352 8309 20380
rect 7708 20340 7714 20352
rect 8297 20349 8309 20352
rect 8343 20380 8355 20383
rect 8386 20380 8392 20392
rect 8343 20352 8392 20380
rect 8343 20349 8355 20352
rect 8297 20343 8355 20349
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8478 20340 8484 20392
rect 8536 20380 8542 20392
rect 8665 20383 8723 20389
rect 8665 20380 8677 20383
rect 8536 20352 8677 20380
rect 8536 20340 8542 20352
rect 8665 20349 8677 20352
rect 8711 20349 8723 20383
rect 8665 20343 8723 20349
rect 8938 20340 8944 20392
rect 8996 20380 9002 20392
rect 9048 20389 9076 20488
rect 11609 20485 11621 20488
rect 11655 20485 11667 20519
rect 11609 20479 11667 20485
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 12621 20519 12679 20525
rect 12621 20516 12633 20519
rect 11848 20488 12633 20516
rect 11848 20476 11854 20488
rect 12621 20485 12633 20488
rect 12667 20485 12679 20519
rect 13078 20516 13084 20528
rect 13039 20488 13084 20516
rect 12621 20479 12679 20485
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 13538 20516 13544 20528
rect 13499 20488 13544 20516
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 13998 20516 14004 20528
rect 13959 20488 14004 20516
rect 13998 20476 14004 20488
rect 14056 20476 14062 20528
rect 14458 20476 14464 20528
rect 14516 20516 14522 20528
rect 14553 20519 14611 20525
rect 14553 20516 14565 20519
rect 14516 20488 14565 20516
rect 14516 20476 14522 20488
rect 14553 20485 14565 20488
rect 14599 20485 14611 20519
rect 14918 20516 14924 20528
rect 14879 20488 14924 20516
rect 14553 20479 14611 20485
rect 14918 20476 14924 20488
rect 14976 20476 14982 20528
rect 15378 20516 15384 20528
rect 15339 20488 15384 20516
rect 15378 20476 15384 20488
rect 15436 20476 15442 20528
rect 15838 20516 15844 20528
rect 15799 20488 15844 20516
rect 15838 20476 15844 20488
rect 15896 20476 15902 20528
rect 16298 20516 16304 20528
rect 16259 20488 16304 20516
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 16758 20516 16764 20528
rect 16719 20488 16764 20516
rect 16758 20476 16764 20488
rect 16816 20476 16822 20528
rect 17678 20516 17684 20528
rect 17639 20488 17684 20516
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 18138 20516 18144 20528
rect 18099 20488 18144 20516
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 18598 20516 18604 20528
rect 18559 20488 18604 20516
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 19058 20516 19064 20528
rect 19019 20488 19064 20516
rect 19058 20476 19064 20488
rect 19116 20476 19122 20528
rect 19518 20476 19524 20528
rect 19576 20516 19582 20528
rect 19889 20519 19947 20525
rect 19889 20516 19901 20519
rect 19576 20488 19901 20516
rect 19576 20476 19582 20488
rect 19889 20485 19901 20488
rect 19935 20485 19947 20519
rect 19889 20479 19947 20485
rect 19978 20476 19984 20528
rect 20036 20516 20042 20528
rect 20257 20519 20315 20525
rect 20257 20516 20269 20519
rect 20036 20488 20269 20516
rect 20036 20476 20042 20488
rect 20257 20485 20269 20488
rect 20303 20485 20315 20519
rect 20257 20479 20315 20485
rect 20438 20476 20444 20528
rect 20496 20516 20502 20528
rect 20625 20519 20683 20525
rect 20625 20516 20637 20519
rect 20496 20488 20637 20516
rect 20496 20476 20502 20488
rect 20625 20485 20637 20488
rect 20671 20485 20683 20519
rect 20625 20479 20683 20485
rect 20898 20476 20904 20528
rect 20956 20516 20962 20528
rect 20993 20519 21051 20525
rect 20993 20516 21005 20519
rect 20956 20488 21005 20516
rect 20956 20476 20962 20488
rect 20993 20485 21005 20488
rect 21039 20485 21051 20519
rect 20993 20479 21051 20485
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9769 20451 9827 20457
rect 9769 20448 9781 20451
rect 9180 20420 9781 20448
rect 9180 20408 9186 20420
rect 9769 20417 9781 20420
rect 9815 20417 9827 20451
rect 9769 20411 9827 20417
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 17589 20451 17647 20457
rect 11112 20420 12848 20448
rect 11112 20408 11118 20420
rect 12360 20392 12388 20420
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8996 20352 9045 20380
rect 8996 20340 9002 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 9398 20340 9404 20392
rect 9456 20380 9462 20392
rect 10226 20380 10232 20392
rect 9456 20352 10232 20380
rect 9456 20340 9462 20352
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10376 20352 10885 20380
rect 10376 20340 10382 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 11296 20352 11437 20380
rect 11296 20340 11302 20352
rect 11425 20349 11437 20352
rect 11471 20380 11483 20383
rect 11471 20352 12204 20380
rect 11471 20349 11483 20352
rect 11425 20343 11483 20349
rect 1670 20312 1676 20324
rect 1631 20284 1676 20312
rect 1670 20272 1676 20284
rect 1728 20272 1734 20324
rect 1946 20312 1952 20324
rect 1907 20284 1952 20312
rect 1946 20272 1952 20284
rect 2004 20272 2010 20324
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 2682 20312 2688 20324
rect 2643 20284 2688 20312
rect 2682 20272 2688 20284
rect 2740 20272 2746 20324
rect 2958 20272 2964 20324
rect 3016 20312 3022 20324
rect 3053 20315 3111 20321
rect 3053 20312 3065 20315
rect 3016 20284 3065 20312
rect 3016 20272 3022 20284
rect 3053 20281 3065 20284
rect 3099 20281 3111 20315
rect 3053 20275 3111 20281
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 3421 20315 3479 20321
rect 3421 20312 3433 20315
rect 3384 20284 3433 20312
rect 3384 20272 3390 20284
rect 3421 20281 3433 20284
rect 3467 20281 3479 20315
rect 3421 20275 3479 20281
rect 3697 20315 3755 20321
rect 3697 20281 3709 20315
rect 3743 20312 3755 20315
rect 4816 20312 4844 20340
rect 3743 20284 4844 20312
rect 4985 20315 5043 20321
rect 3743 20281 3755 20284
rect 3697 20275 3755 20281
rect 4985 20281 4997 20315
rect 5031 20312 5043 20315
rect 5350 20312 5356 20324
rect 5031 20284 5356 20312
rect 5031 20281 5043 20284
rect 4985 20275 5043 20281
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 6932 20312 6960 20340
rect 7742 20312 7748 20324
rect 6932 20284 7604 20312
rect 7703 20284 7748 20312
rect 1854 20244 1860 20256
rect 1815 20216 1860 20244
rect 1854 20204 1860 20216
rect 1912 20204 1918 20256
rect 2774 20204 2780 20256
rect 2832 20244 2838 20256
rect 3510 20244 3516 20256
rect 2832 20216 3516 20244
rect 2832 20204 2838 20216
rect 3510 20204 3516 20216
rect 3568 20204 3574 20256
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4341 20247 4399 20253
rect 4341 20244 4353 20247
rect 4212 20216 4353 20244
rect 4212 20204 4218 20216
rect 4341 20213 4353 20216
rect 4387 20213 4399 20247
rect 4341 20207 4399 20213
rect 5445 20247 5503 20253
rect 5445 20213 5457 20247
rect 5491 20244 5503 20247
rect 5902 20244 5908 20256
rect 5491 20216 5908 20244
rect 5491 20213 5503 20216
rect 5445 20207 5503 20213
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6733 20247 6791 20253
rect 6733 20244 6745 20247
rect 6328 20216 6745 20244
rect 6328 20204 6334 20216
rect 6733 20213 6745 20216
rect 6779 20213 6791 20247
rect 6914 20244 6920 20256
rect 6875 20216 6920 20244
rect 6733 20207 6791 20213
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 7282 20244 7288 20256
rect 7243 20216 7288 20244
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7576 20244 7604 20284
rect 7742 20272 7748 20284
rect 7800 20272 7806 20324
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20281 7987 20315
rect 7929 20275 7987 20281
rect 7650 20244 7656 20256
rect 7432 20216 7477 20244
rect 7563 20216 7656 20244
rect 7432 20204 7438 20216
rect 7650 20204 7656 20216
rect 7708 20244 7714 20256
rect 7944 20244 7972 20275
rect 9306 20272 9312 20324
rect 9364 20312 9370 20324
rect 9677 20315 9735 20321
rect 9677 20312 9689 20315
rect 9364 20284 9689 20312
rect 9364 20272 9370 20284
rect 9677 20281 9689 20284
rect 9723 20281 9735 20315
rect 9677 20275 9735 20281
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 10594 20312 10600 20324
rect 9916 20284 10600 20312
rect 9916 20272 9922 20284
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 11054 20312 11060 20324
rect 11015 20284 11060 20312
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 11698 20272 11704 20324
rect 11756 20312 11762 20324
rect 12066 20312 12072 20324
rect 11756 20284 12072 20312
rect 11756 20272 11762 20284
rect 12066 20272 12072 20284
rect 12124 20272 12130 20324
rect 12176 20312 12204 20352
rect 12342 20340 12348 20392
rect 12400 20340 12406 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 12820 20389 12848 20420
rect 17589 20417 17601 20451
rect 17635 20448 17647 20451
rect 21818 20448 21824 20460
rect 17635 20420 21824 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 12805 20383 12863 20389
rect 12492 20352 12537 20380
rect 12492 20340 12498 20352
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 14185 20383 14243 20389
rect 14185 20380 14197 20383
rect 13688 20352 14197 20380
rect 13688 20340 13694 20352
rect 14185 20349 14197 20352
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 15105 20383 15163 20389
rect 15105 20349 15117 20383
rect 15151 20380 15163 20383
rect 15378 20380 15384 20392
rect 15151 20352 15384 20380
rect 15151 20349 15163 20352
rect 15105 20343 15163 20349
rect 15378 20340 15384 20352
rect 15436 20340 15442 20392
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 18012 20352 21189 20380
rect 18012 20340 18018 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21542 20380 21548 20392
rect 21455 20352 21548 20380
rect 21177 20343 21235 20349
rect 21542 20340 21548 20352
rect 21600 20380 21606 20392
rect 22738 20380 22744 20392
rect 21600 20352 22744 20380
rect 21600 20340 21606 20352
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 12894 20312 12900 20324
rect 12176 20284 12900 20312
rect 12894 20272 12900 20284
rect 12952 20272 12958 20324
rect 13262 20312 13268 20324
rect 13223 20284 13268 20312
rect 13262 20272 13268 20284
rect 13320 20272 13326 20324
rect 13722 20312 13728 20324
rect 13683 20284 13728 20312
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 14366 20272 14372 20324
rect 14424 20312 14430 20324
rect 14737 20315 14795 20321
rect 14737 20312 14749 20315
rect 14424 20284 14749 20312
rect 14424 20272 14430 20284
rect 14737 20281 14749 20284
rect 14783 20281 14795 20315
rect 14737 20275 14795 20281
rect 15194 20272 15200 20324
rect 15252 20312 15258 20324
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 15252 20284 15577 20312
rect 15252 20272 15258 20284
rect 15565 20281 15577 20284
rect 15611 20281 15623 20315
rect 15565 20275 15623 20281
rect 15654 20272 15660 20324
rect 15712 20312 15718 20324
rect 16025 20315 16083 20321
rect 16025 20312 16037 20315
rect 15712 20284 16037 20312
rect 15712 20272 15718 20284
rect 16025 20281 16037 20284
rect 16071 20281 16083 20315
rect 16025 20275 16083 20281
rect 16206 20272 16212 20324
rect 16264 20312 16270 20324
rect 16485 20315 16543 20321
rect 16485 20312 16497 20315
rect 16264 20284 16497 20312
rect 16264 20272 16270 20284
rect 16485 20281 16497 20284
rect 16531 20281 16543 20315
rect 16485 20275 16543 20281
rect 16666 20272 16672 20324
rect 16724 20312 16730 20324
rect 16945 20315 17003 20321
rect 16945 20312 16957 20315
rect 16724 20284 16957 20312
rect 16724 20272 16730 20284
rect 16945 20281 16957 20284
rect 16991 20281 17003 20315
rect 16945 20275 17003 20281
rect 17405 20315 17463 20321
rect 17405 20281 17417 20315
rect 17451 20281 17463 20315
rect 17862 20312 17868 20324
rect 17823 20284 17868 20312
rect 17405 20275 17463 20281
rect 8570 20244 8576 20256
rect 7708 20216 7972 20244
rect 8531 20216 8576 20244
rect 7708 20204 7714 20216
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 9214 20244 9220 20256
rect 9175 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 9585 20247 9643 20253
rect 9585 20244 9597 20247
rect 9456 20216 9597 20244
rect 9456 20204 9462 20216
rect 9585 20213 9597 20216
rect 9631 20213 9643 20247
rect 9585 20207 9643 20213
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 9824 20216 10149 20244
rect 9824 20204 9830 20216
rect 10137 20213 10149 20216
rect 10183 20213 10195 20247
rect 10137 20207 10195 20213
rect 10410 20204 10416 20256
rect 10468 20244 10474 20256
rect 10505 20247 10563 20253
rect 10505 20244 10517 20247
rect 10468 20216 10517 20244
rect 10468 20204 10474 20216
rect 10505 20213 10517 20216
rect 10551 20213 10563 20247
rect 10505 20207 10563 20213
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 11333 20247 11391 20253
rect 11333 20244 11345 20247
rect 11296 20216 11345 20244
rect 11296 20204 11302 20216
rect 11333 20213 11345 20216
rect 11379 20213 11391 20247
rect 11333 20207 11391 20213
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11940 20216 11989 20244
rect 11940 20204 11946 20216
rect 11977 20213 11989 20216
rect 12023 20213 12035 20247
rect 11977 20207 12035 20213
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 12345 20247 12403 20253
rect 12345 20244 12357 20247
rect 12216 20216 12357 20244
rect 12216 20204 12222 20216
rect 12345 20213 12357 20216
rect 12391 20213 12403 20247
rect 12345 20207 12403 20213
rect 12434 20204 12440 20256
rect 12492 20244 12498 20256
rect 13538 20244 13544 20256
rect 12492 20216 13544 20244
rect 12492 20204 12498 20216
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 17420 20244 17448 20275
rect 17862 20272 17868 20284
rect 17920 20272 17926 20324
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 18325 20315 18383 20321
rect 18325 20312 18337 20315
rect 18196 20284 18337 20312
rect 18196 20272 18202 20284
rect 18325 20281 18337 20284
rect 18371 20281 18383 20315
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 18325 20275 18383 20281
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 18874 20272 18880 20324
rect 18932 20312 18938 20324
rect 19245 20315 19303 20321
rect 19245 20312 19257 20315
rect 18932 20284 19257 20312
rect 18932 20272 18938 20284
rect 19245 20281 19257 20284
rect 19291 20281 19303 20315
rect 19518 20312 19524 20324
rect 19479 20284 19524 20312
rect 19245 20275 19303 20281
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 20070 20312 20076 20324
rect 20031 20284 20076 20312
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 20438 20312 20444 20324
rect 20399 20284 20444 20312
rect 20438 20272 20444 20284
rect 20496 20272 20502 20324
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 20809 20315 20867 20321
rect 20809 20312 20821 20315
rect 20588 20284 20821 20312
rect 20588 20272 20594 20284
rect 20809 20281 20821 20284
rect 20855 20281 20867 20315
rect 20809 20275 20867 20281
rect 21358 20244 21364 20256
rect 13872 20216 17448 20244
rect 21319 20216 21364 20244
rect 13872 20204 13878 20216
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1762 20000 1768 20052
rect 1820 20040 1826 20052
rect 1857 20043 1915 20049
rect 1857 20040 1869 20043
rect 1820 20012 1869 20040
rect 1820 20000 1826 20012
rect 1857 20009 1869 20012
rect 1903 20009 1915 20043
rect 2133 20043 2191 20049
rect 2133 20040 2145 20043
rect 1857 20003 1915 20009
rect 1964 20012 2145 20040
rect 1964 19981 1992 20012
rect 2133 20009 2145 20012
rect 2179 20009 2191 20043
rect 2133 20003 2191 20009
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 2682 20040 2688 20052
rect 2639 20012 2688 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20009 3203 20043
rect 3145 20003 3203 20009
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 6454 20040 6460 20052
rect 4387 20012 6460 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 1949 19975 2007 19981
rect 1949 19941 1961 19975
rect 1995 19941 2007 19975
rect 3160 19972 3188 20003
rect 6454 20000 6460 20012
rect 6512 20000 6518 20052
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20009 6975 20043
rect 6917 20003 6975 20009
rect 5166 19972 5172 19984
rect 1949 19935 2007 19941
rect 2240 19944 3004 19972
rect 3160 19944 5172 19972
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19904 1639 19907
rect 2038 19904 2044 19916
rect 1627 19876 2044 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 658 19796 664 19848
rect 716 19836 722 19848
rect 2240 19836 2268 19944
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 716 19808 2268 19836
rect 2332 19836 2360 19867
rect 2406 19864 2412 19916
rect 2464 19904 2470 19916
rect 2866 19904 2872 19916
rect 2464 19876 2509 19904
rect 2827 19876 2872 19904
rect 2464 19864 2470 19876
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 2976 19913 3004 19944
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 6932 19972 6960 20003
rect 8478 20000 8484 20052
rect 8536 20040 8542 20052
rect 8849 20043 8907 20049
rect 8849 20040 8861 20043
rect 8536 20012 8861 20040
rect 8536 20000 8542 20012
rect 8849 20009 8861 20012
rect 8895 20009 8907 20043
rect 8849 20003 8907 20009
rect 8938 20000 8944 20052
rect 8996 20040 9002 20052
rect 11790 20040 11796 20052
rect 8996 20012 11796 20040
rect 8996 20000 9002 20012
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12618 20000 12624 20052
rect 12676 20000 12682 20052
rect 12894 20000 12900 20052
rect 12952 20040 12958 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 12952 20012 13461 20040
rect 12952 20000 12958 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13596 20012 13645 20040
rect 13596 20000 13602 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 17862 20040 17868 20052
rect 16991 20012 17868 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 21542 20040 21548 20052
rect 21503 20012 21548 20040
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 5368 19944 6960 19972
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19904 3019 19907
rect 3142 19904 3148 19916
rect 3007 19876 3148 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 3142 19864 3148 19876
rect 3200 19864 3206 19916
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19904 3295 19907
rect 3418 19904 3424 19916
rect 3283 19876 3424 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 3418 19864 3424 19876
rect 3476 19904 3482 19916
rect 3694 19904 3700 19916
rect 3476 19876 3700 19904
rect 3476 19864 3482 19876
rect 3694 19864 3700 19876
rect 3752 19864 3758 19916
rect 4249 19907 4307 19913
rect 4249 19873 4261 19907
rect 4295 19904 4307 19907
rect 4890 19904 4896 19916
rect 4295 19876 4896 19904
rect 4295 19873 4307 19876
rect 4249 19867 4307 19873
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19904 5043 19907
rect 5258 19904 5264 19916
rect 5031 19876 5264 19904
rect 5031 19873 5043 19876
rect 4985 19867 5043 19873
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 3510 19836 3516 19848
rect 2332 19808 2728 19836
rect 3471 19808 3516 19836
rect 716 19796 722 19808
rect 1394 19768 1400 19780
rect 1355 19740 1400 19768
rect 1394 19728 1400 19740
rect 1452 19728 1458 19780
rect 2700 19777 2728 19808
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 4525 19839 4583 19845
rect 4525 19805 4537 19839
rect 4571 19836 4583 19839
rect 5368 19836 5396 19944
rect 8294 19932 8300 19984
rect 8352 19972 8358 19984
rect 8573 19975 8631 19981
rect 8573 19972 8585 19975
rect 8352 19944 8585 19972
rect 8352 19932 8358 19944
rect 8573 19941 8585 19944
rect 8619 19941 8631 19975
rect 8573 19935 8631 19941
rect 10864 19975 10922 19981
rect 10864 19941 10876 19975
rect 10910 19972 10922 19975
rect 11054 19972 11060 19984
rect 10910 19944 11060 19972
rect 10910 19941 10922 19944
rect 10864 19935 10922 19941
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 12636 19972 12664 20000
rect 13817 19975 13875 19981
rect 13817 19972 13829 19975
rect 12636 19944 13829 19972
rect 6201 19907 6259 19913
rect 6201 19873 6213 19907
rect 6247 19904 6259 19907
rect 6546 19904 6552 19916
rect 6247 19876 6552 19904
rect 6247 19873 6259 19876
rect 6201 19867 6259 19873
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 7098 19904 7104 19916
rect 6687 19876 7104 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7466 19864 7472 19916
rect 7524 19904 7530 19916
rect 8030 19907 8088 19913
rect 8030 19904 8042 19907
rect 7524 19876 8042 19904
rect 7524 19864 7530 19876
rect 8030 19873 8042 19876
rect 8076 19873 8088 19907
rect 8030 19867 8088 19873
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 10238 19907 10296 19913
rect 10238 19904 10250 19907
rect 9180 19876 10250 19904
rect 9180 19864 9186 19876
rect 10238 19873 10250 19876
rect 10284 19873 10296 19907
rect 12066 19904 12072 19916
rect 12027 19876 12072 19904
rect 10238 19867 10296 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19904 12495 19907
rect 12618 19904 12624 19916
rect 12483 19876 12624 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13372 19913 13400 19944
rect 13817 19941 13829 19944
rect 13863 19941 13875 19975
rect 17218 19972 17224 19984
rect 17179 19944 17224 19972
rect 13817 19935 13875 19941
rect 17218 19932 17224 19944
rect 17276 19932 17282 19984
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19873 12955 19907
rect 12897 19867 12955 19873
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19873 13415 19907
rect 13357 19867 13415 19873
rect 6454 19836 6460 19848
rect 4571 19808 5396 19836
rect 6415 19808 6460 19836
rect 4571 19805 4583 19808
rect 4525 19799 4583 19805
rect 2685 19771 2743 19777
rect 2685 19737 2697 19771
rect 2731 19737 2743 19771
rect 2685 19731 2743 19737
rect 3050 19728 3056 19780
rect 3108 19768 3114 19780
rect 3881 19771 3939 19777
rect 3881 19768 3893 19771
rect 3108 19740 3893 19768
rect 3108 19728 3114 19740
rect 3881 19737 3893 19740
rect 3927 19737 3939 19771
rect 3881 19731 3939 19737
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 4540 19768 4568 19799
rect 6454 19796 6460 19808
rect 6512 19796 6518 19848
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 10502 19836 10508 19848
rect 10463 19808 10508 19836
rect 8297 19799 8355 19805
rect 5350 19768 5356 19780
rect 4304 19740 4568 19768
rect 4632 19740 5356 19768
rect 4304 19728 4310 19740
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 4632 19700 4660 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 4798 19700 4804 19712
rect 3467 19672 4660 19700
rect 4759 19672 4804 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5810 19700 5816 19712
rect 5123 19672 5816 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 6472 19700 6500 19796
rect 6825 19771 6883 19777
rect 6825 19737 6837 19771
rect 6871 19768 6883 19771
rect 7006 19768 7012 19780
rect 6871 19740 7012 19768
rect 6871 19737 6883 19740
rect 6825 19731 6883 19737
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 8312 19700 8340 19799
rect 10502 19796 10508 19808
rect 10560 19836 10566 19848
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 10560 19808 10609 19836
rect 10560 19796 10566 19808
rect 10597 19805 10609 19808
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12400 19808 12725 19836
rect 12400 19796 12406 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 12912 19836 12940 19867
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 16761 19907 16819 19913
rect 16761 19904 16773 19907
rect 16632 19876 16773 19904
rect 16632 19864 16638 19876
rect 16761 19873 16773 19876
rect 16807 19873 16819 19907
rect 17402 19904 17408 19916
rect 17363 19876 17408 19904
rect 16761 19867 16819 19873
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 12860 19808 12940 19836
rect 12860 19796 12866 19808
rect 8389 19771 8447 19777
rect 8389 19737 8401 19771
rect 8435 19768 8447 19771
rect 8754 19768 8760 19780
rect 8435 19740 8760 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 8754 19728 8760 19740
rect 8812 19728 8818 19780
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 13173 19771 13231 19777
rect 13173 19768 13185 19771
rect 11848 19740 13185 19768
rect 11848 19728 11854 19740
rect 13173 19737 13185 19740
rect 13219 19737 13231 19771
rect 13173 19731 13231 19737
rect 8478 19700 8484 19712
rect 6472 19672 8484 19700
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 9125 19703 9183 19709
rect 9125 19700 9137 19703
rect 8720 19672 9137 19700
rect 8720 19660 8726 19672
rect 9125 19669 9137 19672
rect 9171 19669 9183 19703
rect 11974 19700 11980 19712
rect 11935 19672 11980 19700
rect 9125 19663 9183 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 12526 19700 12532 19712
rect 12299 19672 12532 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 12621 19703 12679 19709
rect 12621 19669 12633 19703
rect 12667 19700 12679 19703
rect 12986 19700 12992 19712
rect 12667 19672 12992 19700
rect 12667 19669 12679 19672
rect 12621 19663 12679 19669
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13814 19700 13820 19712
rect 13127 19672 13820 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 14274 19660 14280 19712
rect 14332 19700 14338 19712
rect 14369 19703 14427 19709
rect 14369 19700 14381 19703
rect 14332 19672 14381 19700
rect 14332 19660 14338 19672
rect 14369 19669 14381 19672
rect 14415 19669 14427 19703
rect 16574 19700 16580 19712
rect 16535 19672 16580 19700
rect 14369 19663 14427 19669
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1765 19499 1823 19505
rect 1765 19465 1777 19499
rect 1811 19496 1823 19499
rect 1946 19496 1952 19508
rect 1811 19468 1952 19496
rect 1811 19465 1823 19468
rect 1765 19459 1823 19465
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2041 19499 2099 19505
rect 2041 19465 2053 19499
rect 2087 19496 2099 19499
rect 2314 19496 2320 19508
rect 2087 19468 2320 19496
rect 2087 19465 2099 19468
rect 2041 19459 2099 19465
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 2866 19456 2872 19508
rect 2924 19496 2930 19508
rect 3053 19499 3111 19505
rect 3053 19496 3065 19499
rect 2924 19468 3065 19496
rect 2924 19456 2930 19468
rect 3053 19465 3065 19468
rect 3099 19465 3111 19499
rect 3053 19459 3111 19465
rect 3344 19468 4660 19496
rect 3344 19428 3372 19468
rect 2424 19400 3372 19428
rect 1946 19292 1952 19304
rect 1907 19264 1952 19292
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19292 2283 19295
rect 2424 19292 2452 19400
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 4632 19360 4660 19468
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 7101 19499 7159 19505
rect 5408 19468 7052 19496
rect 5408 19456 5414 19468
rect 7024 19428 7052 19468
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7466 19496 7472 19508
rect 7147 19468 7472 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7466 19456 7472 19468
rect 7524 19456 7530 19508
rect 9122 19496 9128 19508
rect 7576 19468 8984 19496
rect 9083 19468 9128 19496
rect 7576 19428 7604 19468
rect 7024 19400 7604 19428
rect 8956 19428 8984 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 10226 19456 10232 19508
rect 10284 19496 10290 19508
rect 10597 19499 10655 19505
rect 10597 19496 10609 19499
rect 10284 19468 10609 19496
rect 10284 19456 10290 19468
rect 10597 19465 10609 19468
rect 10643 19465 10655 19499
rect 10597 19459 10655 19465
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13357 19499 13415 19505
rect 13357 19496 13369 19499
rect 13320 19468 13369 19496
rect 13320 19456 13326 19468
rect 13357 19465 13369 19468
rect 13403 19465 13415 19499
rect 13357 19459 13415 19465
rect 13633 19499 13691 19505
rect 13633 19465 13645 19499
rect 13679 19496 13691 19499
rect 13722 19496 13728 19508
rect 13679 19468 13728 19496
rect 13679 19465 13691 19468
rect 13633 19459 13691 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 13909 19499 13967 19505
rect 13909 19465 13921 19499
rect 13955 19496 13967 19499
rect 14366 19496 14372 19508
rect 13955 19468 14372 19496
rect 13955 19465 13967 19468
rect 13909 19459 13967 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 15654 19496 15660 19508
rect 15335 19468 15660 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 16206 19496 16212 19508
rect 15887 19468 16212 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 17402 19496 17408 19508
rect 16531 19468 17408 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 18196 19468 18245 19496
rect 18196 19456 18202 19468
rect 18233 19465 18245 19468
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 18509 19499 18567 19505
rect 18509 19465 18521 19499
rect 18555 19496 18567 19499
rect 18782 19496 18788 19508
rect 18555 19468 18788 19496
rect 18555 19465 18567 19468
rect 18509 19459 18567 19465
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20530 19496 20536 19508
rect 19843 19468 20536 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 9490 19428 9496 19440
rect 8956 19400 9496 19428
rect 9490 19388 9496 19400
rect 9548 19388 9554 19440
rect 15013 19431 15071 19437
rect 15013 19397 15025 19431
rect 15059 19428 15071 19431
rect 15378 19428 15384 19440
rect 15059 19400 15384 19428
rect 15059 19397 15071 19400
rect 15013 19391 15071 19397
rect 15378 19388 15384 19400
rect 15436 19388 15442 19440
rect 19245 19431 19303 19437
rect 19245 19397 19257 19431
rect 19291 19428 19303 19431
rect 20438 19428 20444 19440
rect 19291 19400 20444 19428
rect 19291 19397 19303 19400
rect 19245 19391 19303 19397
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 2547 19332 2636 19360
rect 4632 19332 4752 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 2271 19264 2452 19292
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 1394 19224 1400 19236
rect 1355 19196 1400 19224
rect 1394 19184 1400 19196
rect 1452 19184 1458 19236
rect 1578 19224 1584 19236
rect 1539 19196 1584 19224
rect 1578 19184 1584 19196
rect 1636 19184 1642 19236
rect 2608 19224 2636 19332
rect 2685 19295 2743 19301
rect 2685 19261 2697 19295
rect 2731 19292 2743 19295
rect 3510 19292 3516 19304
rect 2731 19264 3516 19292
rect 2731 19261 2743 19264
rect 2685 19255 2743 19261
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 4246 19292 4252 19304
rect 4304 19301 4310 19304
rect 4216 19264 4252 19292
rect 4246 19252 4252 19264
rect 4304 19255 4316 19301
rect 4525 19295 4583 19301
rect 4525 19292 4537 19295
rect 4356 19264 4537 19292
rect 4304 19252 4310 19255
rect 2608 19196 3188 19224
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 3050 19156 3056 19168
rect 2639 19128 3056 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3160 19165 3188 19196
rect 3786 19184 3792 19236
rect 3844 19224 3850 19236
rect 4356 19224 4384 19264
rect 4525 19261 4537 19264
rect 4571 19292 4583 19295
rect 4617 19295 4675 19301
rect 4617 19292 4629 19295
rect 4571 19264 4629 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 4617 19261 4629 19264
rect 4663 19261 4675 19295
rect 4724 19292 4752 19332
rect 5902 19320 5908 19372
rect 5960 19360 5966 19372
rect 7009 19363 7067 19369
rect 5960 19332 6132 19360
rect 5960 19320 5966 19332
rect 6104 19301 6132 19332
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7282 19360 7288 19372
rect 7055 19332 7288 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 8478 19360 8484 19372
rect 8439 19332 8484 19360
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 8662 19360 8668 19372
rect 8588 19332 8668 19360
rect 6089 19295 6147 19301
rect 4724 19264 5939 19292
rect 4617 19255 4675 19261
rect 4862 19227 4920 19233
rect 4862 19224 4874 19227
rect 3844 19196 4384 19224
rect 4428 19196 4874 19224
rect 3844 19184 3850 19196
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 4428 19156 4456 19196
rect 4862 19193 4874 19196
rect 4908 19193 4920 19227
rect 5911 19224 5939 19264
rect 6089 19261 6101 19295
rect 6135 19261 6147 19295
rect 6089 19255 6147 19261
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19292 6791 19295
rect 6914 19292 6920 19304
rect 6779 19264 6920 19292
rect 6779 19261 6791 19264
rect 6733 19255 6791 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 8236 19227 8294 19233
rect 5911 19196 6592 19224
rect 4862 19187 4920 19193
rect 3191 19128 4456 19156
rect 5997 19159 6055 19165
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 5997 19125 6009 19159
rect 6043 19156 6055 19159
rect 6454 19156 6460 19168
rect 6043 19128 6460 19156
rect 6043 19125 6055 19128
rect 5997 19119 6055 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6564 19165 6592 19196
rect 8236 19193 8248 19227
rect 8282 19224 8294 19227
rect 8588 19224 8616 19332
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 9033 19363 9091 19369
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9398 19360 9404 19372
rect 9079 19332 9404 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 11425 19363 11483 19369
rect 11425 19329 11437 19363
rect 11471 19360 11483 19363
rect 11471 19332 11836 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19292 8815 19295
rect 9214 19292 9220 19304
rect 8803 19264 9220 19292
rect 8803 19261 8815 19264
rect 8757 19255 8815 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 10502 19292 10508 19304
rect 10463 19264 10508 19292
rect 10502 19252 10508 19264
rect 10560 19292 10566 19304
rect 11701 19295 11759 19301
rect 11701 19292 11713 19295
rect 10560 19264 11713 19292
rect 10560 19252 10566 19264
rect 11701 19261 11713 19264
rect 11747 19261 11759 19295
rect 11808 19292 11836 19332
rect 12986 19320 12992 19372
rect 13044 19360 13050 19372
rect 20070 19360 20076 19372
rect 13044 19332 13492 19360
rect 13044 19320 13050 19332
rect 11974 19301 11980 19304
rect 11968 19292 11980 19301
rect 11808 19264 11980 19292
rect 11701 19255 11759 19261
rect 11968 19255 11980 19264
rect 11974 19252 11980 19255
rect 12032 19252 12038 19304
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 13464 19301 13492 19332
rect 17880 19332 20076 19360
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12584 19264 13185 19292
rect 12584 19252 12590 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13722 19292 13728 19304
rect 13683 19264 13728 19292
rect 13449 19255 13507 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13872 19264 14013 19292
rect 13872 19252 13878 19264
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 8282 19196 8616 19224
rect 8282 19193 8294 19196
rect 8236 19187 8294 19193
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10260 19227 10318 19233
rect 10260 19224 10272 19227
rect 10008 19196 10272 19224
rect 10008 19184 10014 19196
rect 10260 19193 10272 19196
rect 10306 19224 10318 19227
rect 14016 19224 14044 19255
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14332 19264 14473 19292
rect 14332 19252 14338 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 14550 19252 14556 19304
rect 14608 19292 14614 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14608 19264 14841 19292
rect 14608 19252 14614 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15286 19292 15292 19304
rect 15151 19264 15292 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15286 19252 15292 19264
rect 15344 19292 15350 19304
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 15344 19264 15393 19292
rect 15344 19252 15350 19264
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15620 19264 15669 19292
rect 15620 19252 15626 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 15930 19292 15936 19304
rect 15891 19264 15936 19292
rect 15657 19255 15715 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 16301 19295 16359 19301
rect 16301 19292 16313 19295
rect 16172 19264 16313 19292
rect 16172 19252 16178 19264
rect 16301 19261 16313 19264
rect 16347 19261 16359 19295
rect 16301 19255 16359 19261
rect 16390 19252 16396 19304
rect 16448 19292 16454 19304
rect 16577 19295 16635 19301
rect 16577 19292 16589 19295
rect 16448 19264 16589 19292
rect 16448 19252 16454 19264
rect 16577 19261 16589 19264
rect 16623 19261 16635 19295
rect 17880 19292 17908 19332
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 16577 19255 16635 19261
rect 16960 19264 17908 19292
rect 17957 19295 18015 19301
rect 14369 19227 14427 19233
rect 14369 19224 14381 19227
rect 10306 19196 12434 19224
rect 14016 19196 14381 19224
rect 10306 19193 10318 19196
rect 10260 19187 10318 19193
rect 6549 19159 6607 19165
rect 6549 19125 6561 19159
rect 6595 19125 6607 19159
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 6549 19119 6607 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 11698 19156 11704 19168
rect 11287 19128 11704 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12406 19156 12434 19196
rect 14369 19193 14381 19196
rect 14415 19193 14427 19227
rect 16960 19224 16988 19264
rect 17957 19261 17969 19295
rect 18003 19261 18015 19295
rect 17957 19255 18015 19261
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18138 19292 18144 19304
rect 18095 19264 18144 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 17126 19224 17132 19236
rect 14369 19187 14427 19193
rect 14568 19196 16988 19224
rect 17087 19196 17132 19224
rect 13081 19159 13139 19165
rect 13081 19156 13093 19159
rect 12406 19128 13093 19156
rect 13081 19125 13093 19128
rect 13127 19125 13139 19159
rect 13081 19119 13139 19125
rect 14185 19159 14243 19165
rect 14185 19125 14197 19159
rect 14231 19156 14243 19159
rect 14568 19156 14596 19196
rect 17126 19184 17132 19196
rect 17184 19184 17190 19236
rect 17972 19224 18000 19255
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 18322 19292 18328 19304
rect 18283 19264 18328 19292
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 18598 19292 18604 19304
rect 18559 19264 18604 19292
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 19058 19292 19064 19304
rect 18971 19264 19064 19292
rect 19058 19252 19064 19264
rect 19116 19292 19122 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19116 19264 19349 19292
rect 19116 19252 19122 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19610 19292 19616 19304
rect 19571 19264 19616 19292
rect 19337 19255 19395 19261
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 18969 19227 19027 19233
rect 18969 19224 18981 19227
rect 17972 19196 18981 19224
rect 18969 19193 18981 19196
rect 19015 19224 19027 19227
rect 22278 19224 22284 19236
rect 19015 19196 22284 19224
rect 19015 19193 19027 19196
rect 18969 19187 19027 19193
rect 22278 19184 22284 19196
rect 22336 19184 22342 19236
rect 14231 19128 14596 19156
rect 14645 19159 14703 19165
rect 14231 19125 14243 19128
rect 14185 19119 14243 19125
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 15194 19156 15200 19168
rect 14691 19128 15200 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16666 19156 16672 19168
rect 16163 19128 16672 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17954 19156 17960 19168
rect 16807 19128 17960 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18782 19156 18788 19168
rect 18743 19128 18788 19156
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 1765 18955 1823 18961
rect 1765 18952 1777 18955
rect 1636 18924 1777 18952
rect 1636 18912 1642 18924
rect 1765 18921 1777 18924
rect 1811 18921 1823 18955
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 1765 18915 1823 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 2593 18955 2651 18961
rect 2593 18952 2605 18955
rect 2464 18924 2605 18952
rect 2464 18912 2470 18924
rect 2593 18921 2605 18924
rect 2639 18921 2651 18955
rect 2869 18955 2927 18961
rect 2869 18952 2881 18955
rect 2593 18915 2651 18921
rect 2746 18924 2881 18952
rect 2746 18884 2774 18924
rect 2869 18921 2881 18924
rect 2915 18921 2927 18955
rect 2869 18915 2927 18921
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3510 18952 3516 18964
rect 3292 18924 3516 18952
rect 3292 18912 3298 18924
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 3660 18924 4752 18952
rect 3660 18912 3666 18924
rect 4246 18884 4252 18896
rect 2332 18856 2774 18884
rect 4207 18856 4252 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 1762 18816 1768 18828
rect 1627 18788 1768 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2038 18816 2044 18828
rect 1995 18788 2044 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 2332 18825 2360 18856
rect 4246 18844 4252 18856
rect 4304 18844 4310 18896
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18785 2283 18819
rect 2225 18779 2283 18785
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18785 2375 18819
rect 2317 18779 2375 18785
rect 2240 18748 2268 18779
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 3053 18819 3111 18825
rect 2832 18788 2877 18816
rect 2832 18776 2838 18788
rect 3053 18785 3065 18819
rect 3099 18785 3111 18819
rect 3053 18779 3111 18785
rect 3145 18819 3203 18825
rect 3145 18785 3157 18819
rect 3191 18816 3203 18819
rect 3234 18816 3240 18828
rect 3191 18788 3240 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 2406 18748 2412 18760
rect 2240 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 3068 18748 3096 18779
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18816 3479 18819
rect 3510 18816 3516 18828
rect 3467 18788 3516 18816
rect 3467 18785 3479 18788
rect 3421 18779 3479 18785
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 4724 18825 4752 18924
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 5592 18924 6561 18952
rect 5592 18912 5598 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 7006 18952 7012 18964
rect 6967 18924 7012 18952
rect 6549 18915 6607 18921
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7374 18952 7380 18964
rect 7335 18924 7380 18952
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8205 18955 8263 18961
rect 8205 18952 8217 18955
rect 7708 18924 8217 18952
rect 7708 18912 7714 18924
rect 8205 18921 8217 18924
rect 8251 18921 8263 18955
rect 8386 18952 8392 18964
rect 8347 18924 8392 18952
rect 8205 18915 8263 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9306 18952 9312 18964
rect 9267 18924 9312 18952
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 10318 18912 10324 18964
rect 10376 18952 10382 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10376 18924 10609 18952
rect 10376 18912 10382 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10744 18924 11069 18952
rect 10744 18912 10750 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 11204 18924 11529 18952
rect 11204 18912 11210 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 11698 18952 11704 18964
rect 11659 18924 11704 18952
rect 11517 18915 11575 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 12158 18952 12164 18964
rect 12119 18924 12164 18952
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 12529 18955 12587 18961
rect 12529 18952 12541 18955
rect 12308 18924 12541 18952
rect 12308 18912 12314 18924
rect 12529 18921 12541 18924
rect 12575 18921 12587 18955
rect 12529 18915 12587 18921
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13722 18952 13728 18964
rect 13679 18924 13728 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18952 14243 18955
rect 14550 18952 14556 18964
rect 14231 18924 14556 18952
rect 14231 18921 14243 18924
rect 14185 18915 14243 18921
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 15013 18955 15071 18961
rect 15013 18921 15025 18955
rect 15059 18952 15071 18955
rect 15930 18952 15936 18964
rect 15059 18924 15936 18952
rect 15059 18921 15071 18924
rect 15013 18915 15071 18921
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18952 16911 18955
rect 18322 18952 18328 18964
rect 16899 18924 18328 18952
rect 16899 18921 16911 18924
rect 16853 18915 16911 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 18877 18955 18935 18961
rect 18877 18921 18889 18955
rect 18923 18952 18935 18955
rect 19610 18952 19616 18964
rect 18923 18924 19616 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6190 18887 6248 18893
rect 6190 18884 6202 18887
rect 5868 18856 6202 18884
rect 5868 18844 5874 18856
rect 6190 18853 6202 18856
rect 6236 18853 6248 18887
rect 6190 18847 6248 18853
rect 6454 18844 6460 18896
rect 6512 18884 6518 18896
rect 6917 18887 6975 18893
rect 6917 18884 6929 18887
rect 6512 18856 6929 18884
rect 6512 18844 6518 18856
rect 6917 18853 6929 18856
rect 6963 18853 6975 18887
rect 6917 18847 6975 18853
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 8573 18887 8631 18893
rect 8573 18884 8585 18887
rect 8352 18856 8585 18884
rect 8352 18844 8358 18856
rect 8573 18853 8585 18856
rect 8619 18853 8631 18887
rect 8573 18847 8631 18853
rect 9769 18887 9827 18893
rect 9769 18853 9781 18887
rect 9815 18884 9827 18887
rect 11790 18884 11796 18896
rect 9815 18856 11796 18884
rect 9815 18853 9827 18856
rect 9769 18847 9827 18853
rect 11790 18844 11796 18856
rect 11848 18844 11854 18896
rect 12176 18884 12204 18912
rect 12805 18887 12863 18893
rect 12805 18884 12817 18887
rect 12176 18856 12817 18884
rect 12805 18853 12817 18856
rect 12851 18884 12863 18887
rect 15562 18884 15568 18896
rect 12851 18856 14688 18884
rect 15523 18856 15568 18884
rect 12851 18853 12863 18856
rect 12805 18847 12863 18853
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 4982 18816 4988 18828
rect 4755 18788 4988 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 4982 18776 4988 18788
rect 5040 18776 5046 18828
rect 6362 18776 6368 18828
rect 6420 18776 6426 18828
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7340 18788 7757 18816
rect 7340 18776 7346 18788
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8938 18816 8944 18828
rect 7883 18788 8944 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 9214 18816 9220 18828
rect 9127 18788 9220 18816
rect 9214 18776 9220 18788
rect 9272 18816 9278 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9272 18788 9689 18816
rect 9272 18776 9278 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 10321 18819 10379 18825
rect 10321 18785 10333 18819
rect 10367 18816 10379 18819
rect 10778 18816 10784 18828
rect 10367 18788 10784 18816
rect 10367 18785 10379 18788
rect 10321 18779 10379 18785
rect 10778 18776 10784 18788
rect 10836 18776 10842 18828
rect 11146 18816 11152 18828
rect 11107 18788 11152 18816
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18816 12127 18819
rect 12710 18816 12716 18828
rect 12115 18788 12716 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 13998 18816 14004 18828
rect 13959 18788 14004 18816
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 14458 18816 14464 18828
rect 14371 18788 14464 18816
rect 14458 18776 14464 18788
rect 14516 18816 14522 18828
rect 14553 18819 14611 18825
rect 14553 18816 14565 18819
rect 14516 18788 14565 18816
rect 14516 18776 14522 18788
rect 14553 18785 14565 18788
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 3068 18720 3924 18748
rect 2501 18683 2559 18689
rect 2501 18649 2513 18683
rect 2547 18680 2559 18683
rect 2958 18680 2964 18692
rect 2547 18652 2964 18680
rect 2547 18649 2559 18652
rect 2501 18643 2559 18649
rect 2958 18640 2964 18652
rect 3016 18640 3022 18692
rect 3329 18683 3387 18689
rect 3329 18649 3341 18683
rect 3375 18680 3387 18683
rect 3510 18680 3516 18692
rect 3375 18652 3516 18680
rect 3375 18649 3387 18652
rect 3329 18643 3387 18649
rect 3510 18640 3516 18652
rect 3568 18640 3574 18692
rect 3896 18689 3924 18720
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 4525 18751 4583 18757
rect 4396 18720 4441 18748
rect 4396 18708 4402 18720
rect 4525 18717 4537 18751
rect 4571 18717 4583 18751
rect 5166 18748 5172 18760
rect 4525 18711 4583 18717
rect 4816 18720 5172 18748
rect 3881 18683 3939 18689
rect 3881 18649 3893 18683
rect 3927 18649 3939 18683
rect 3881 18643 3939 18649
rect 3970 18640 3976 18692
rect 4028 18680 4034 18692
rect 4540 18680 4568 18711
rect 4028 18652 4568 18680
rect 4028 18640 4034 18652
rect 2590 18572 2596 18624
rect 2648 18612 2654 18624
rect 3234 18612 3240 18624
rect 2648 18584 3240 18612
rect 2648 18572 2654 18584
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 3605 18615 3663 18621
rect 3605 18581 3617 18615
rect 3651 18612 3663 18615
rect 4816 18612 4844 18720
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 6380 18748 6408 18776
rect 6457 18751 6515 18757
rect 6457 18748 6469 18751
rect 6380 18720 6469 18748
rect 6457 18717 6469 18720
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 6546 18708 6552 18760
rect 6604 18748 6610 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 6604 18720 7113 18748
rect 6604 18708 6610 18720
rect 7101 18717 7113 18720
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 8021 18751 8079 18757
rect 8021 18717 8033 18751
rect 8067 18748 8079 18751
rect 8662 18748 8668 18760
rect 8067 18720 8668 18748
rect 8067 18717 8079 18720
rect 8021 18711 8079 18717
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 9950 18748 9956 18760
rect 9911 18720 9956 18748
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 10686 18748 10692 18760
rect 10551 18720 10692 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 4893 18683 4951 18689
rect 4893 18649 4905 18683
rect 4939 18680 4951 18683
rect 5350 18680 5356 18692
rect 4939 18652 5356 18680
rect 4939 18649 4951 18652
rect 4893 18643 4951 18649
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 6638 18640 6644 18692
rect 6696 18680 6702 18692
rect 10137 18683 10195 18689
rect 10137 18680 10149 18683
rect 6696 18652 10149 18680
rect 6696 18640 6702 18652
rect 10137 18649 10149 18652
rect 10183 18649 10195 18683
rect 10137 18643 10195 18649
rect 5074 18612 5080 18624
rect 3651 18584 4844 18612
rect 5035 18584 5080 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 10520 18612 10548 18711
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 12342 18748 12348 18760
rect 12303 18720 12348 18748
rect 10965 18711 11023 18717
rect 10980 18680 11008 18711
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 14660 18748 14688 18856
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 14826 18816 14832 18828
rect 14787 18788 14832 18816
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 16666 18816 16672 18828
rect 16627 18788 16672 18816
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 18690 18816 18696 18828
rect 18651 18788 18696 18816
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 17310 18748 17316 18760
rect 14660 18720 17316 18748
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 12360 18680 12388 18708
rect 10980 18652 12388 18680
rect 14737 18683 14795 18689
rect 11072 18624 11100 18652
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 19518 18680 19524 18692
rect 14783 18652 19524 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 6604 18584 10548 18612
rect 6604 18572 6610 18584
rect 11054 18572 11060 18624
rect 11112 18572 11118 18624
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 17954 18612 17960 18624
rect 17915 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 18417 18615 18475 18621
rect 18417 18612 18429 18615
rect 18196 18584 18429 18612
rect 18196 18572 18202 18584
rect 18417 18581 18429 18584
rect 18463 18612 18475 18615
rect 18598 18612 18604 18624
rect 18463 18584 18604 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2958 18408 2964 18420
rect 2004 18380 2964 18408
rect 2004 18368 2010 18380
rect 2958 18368 2964 18380
rect 3016 18368 3022 18420
rect 3234 18368 3240 18420
rect 3292 18408 3298 18420
rect 3970 18408 3976 18420
rect 3292 18380 3556 18408
rect 3931 18380 3976 18408
rect 3292 18368 3298 18380
rect 2498 18340 2504 18352
rect 2459 18312 2504 18340
rect 2498 18300 2504 18312
rect 2556 18300 2562 18352
rect 3528 18340 3556 18380
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4338 18408 4344 18420
rect 4299 18380 4344 18408
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 5258 18408 5264 18420
rect 5219 18380 5264 18408
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5718 18408 5724 18420
rect 5679 18380 5724 18408
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6457 18411 6515 18417
rect 6457 18408 6469 18411
rect 6236 18380 6469 18408
rect 6236 18368 6242 18380
rect 6457 18377 6469 18380
rect 6503 18377 6515 18411
rect 6457 18371 6515 18377
rect 7009 18411 7067 18417
rect 7009 18377 7021 18411
rect 7055 18408 7067 18411
rect 7098 18408 7104 18420
rect 7055 18380 7104 18408
rect 7055 18377 7067 18380
rect 7009 18371 7067 18377
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 9214 18408 9220 18420
rect 7616 18380 9220 18408
rect 7616 18368 7622 18380
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 12066 18408 12072 18420
rect 10376 18380 12072 18408
rect 10376 18368 10382 18380
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 5353 18343 5411 18349
rect 5353 18340 5365 18343
rect 3528 18312 5365 18340
rect 5353 18309 5365 18312
rect 5399 18309 5411 18343
rect 5353 18303 5411 18309
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 9674 18340 9680 18352
rect 5500 18312 9680 18340
rect 5500 18300 5506 18312
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18232 1458 18284
rect 1486 18232 1492 18284
rect 1544 18272 1550 18284
rect 4246 18272 4252 18284
rect 1544 18244 2728 18272
rect 4207 18244 4252 18272
rect 1544 18232 1550 18244
rect 2056 18213 2084 18244
rect 1949 18207 2007 18213
rect 1949 18173 1961 18207
rect 1995 18173 2007 18207
rect 1949 18167 2007 18173
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 1578 18136 1584 18148
rect 1539 18108 1584 18136
rect 1578 18096 1584 18108
rect 1636 18096 1642 18148
rect 1964 18136 1992 18167
rect 2130 18164 2136 18216
rect 2188 18204 2194 18216
rect 2314 18204 2320 18216
rect 2188 18176 2320 18204
rect 2188 18164 2194 18176
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 2498 18136 2504 18148
rect 1964 18108 2504 18136
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 2222 18068 2228 18080
rect 2183 18040 2228 18068
rect 2222 18028 2228 18040
rect 2280 18028 2286 18080
rect 2608 18068 2636 18167
rect 2700 18136 2728 18244
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 4798 18272 4804 18284
rect 4759 18244 4804 18272
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5074 18272 5080 18284
rect 4939 18244 5080 18272
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 2860 18207 2918 18213
rect 2860 18173 2872 18207
rect 2906 18204 2918 18207
rect 4908 18204 4936 18235
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 9122 18272 9128 18284
rect 5316 18244 9128 18272
rect 5316 18232 5322 18244
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9401 18275 9459 18281
rect 9401 18272 9413 18275
rect 9364 18244 9413 18272
rect 9364 18232 9370 18244
rect 9401 18241 9413 18244
rect 9447 18241 9459 18275
rect 11146 18272 11152 18284
rect 11107 18244 11152 18272
rect 9401 18235 9459 18241
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 12124 18244 12265 18272
rect 12124 18232 12130 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 5994 18204 6000 18216
rect 2906 18176 4936 18204
rect 5907 18176 6000 18204
rect 2906 18173 2918 18176
rect 2860 18167 2918 18173
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 6052 18176 8800 18204
rect 6052 18164 6058 18176
rect 3510 18136 3516 18148
rect 2700 18108 3516 18136
rect 3510 18096 3516 18108
rect 3568 18096 3574 18148
rect 8570 18136 8576 18148
rect 3620 18108 8576 18136
rect 2866 18068 2872 18080
rect 2608 18040 2872 18068
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3620 18068 3648 18108
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8772 18145 8800 18176
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 16666 18204 16672 18216
rect 10744 18176 16672 18204
rect 10744 18164 10750 18176
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 9309 18139 9367 18145
rect 9309 18136 9321 18139
rect 8803 18108 9321 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 9309 18105 9321 18108
rect 9355 18105 9367 18139
rect 9309 18099 9367 18105
rect 13906 18096 13912 18148
rect 13964 18136 13970 18148
rect 14826 18136 14832 18148
rect 13964 18108 14832 18136
rect 13964 18096 13970 18108
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 3016 18040 3648 18068
rect 3016 18028 3022 18040
rect 3694 18028 3700 18080
rect 3752 18068 3758 18080
rect 4614 18068 4620 18080
rect 3752 18040 4620 18068
rect 3752 18028 3758 18040
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 4706 18028 4712 18080
rect 4764 18068 4770 18080
rect 4764 18040 4809 18068
rect 4764 18028 4770 18040
rect 4890 18028 4896 18080
rect 4948 18068 4954 18080
rect 5166 18068 5172 18080
rect 4948 18040 5172 18068
rect 4948 18028 4954 18040
rect 5166 18028 5172 18040
rect 5224 18068 5230 18080
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 5224 18040 5549 18068
rect 5224 18028 5230 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 5537 18031 5595 18037
rect 6454 18028 6460 18080
rect 6512 18068 6518 18080
rect 6641 18071 6699 18077
rect 6641 18068 6653 18071
rect 6512 18040 6653 18068
rect 6512 18028 6518 18040
rect 6641 18037 6653 18040
rect 6687 18037 6699 18071
rect 7282 18068 7288 18080
rect 7243 18040 7288 18068
rect 6641 18031 6699 18037
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 8846 18068 8852 18080
rect 8807 18040 8852 18068
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11112 18040 11713 18068
rect 11112 18028 11118 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 11790 18028 11796 18080
rect 11848 18068 11854 18080
rect 12069 18071 12127 18077
rect 12069 18068 12081 18071
rect 11848 18040 12081 18068
rect 11848 18028 11854 18040
rect 12069 18037 12081 18040
rect 12115 18037 12127 18071
rect 12069 18031 12127 18037
rect 12158 18028 12164 18080
rect 12216 18068 12222 18080
rect 12216 18040 12261 18068
rect 12216 18028 12222 18040
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1486 17864 1492 17876
rect 1447 17836 1492 17864
rect 1486 17824 1492 17836
rect 1544 17824 1550 17876
rect 1578 17824 1584 17876
rect 1636 17864 1642 17876
rect 1765 17867 1823 17873
rect 1765 17864 1777 17867
rect 1636 17836 1777 17864
rect 1636 17824 1642 17836
rect 1765 17833 1777 17836
rect 1811 17833 1823 17867
rect 1765 17827 1823 17833
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 2332 17796 2360 17827
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 2593 17867 2651 17873
rect 2593 17864 2605 17867
rect 2556 17836 2605 17864
rect 2556 17824 2562 17836
rect 2593 17833 2605 17836
rect 2639 17833 2651 17867
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 2593 17827 2651 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 3510 17864 3516 17876
rect 3471 17836 3516 17864
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4433 17867 4491 17873
rect 4433 17864 4445 17867
rect 4212 17836 4445 17864
rect 4212 17824 4218 17836
rect 4433 17833 4445 17836
rect 4479 17833 4491 17867
rect 4433 17827 4491 17833
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4672 17836 4813 17864
rect 4672 17824 4678 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 4801 17827 4859 17833
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4948 17836 4997 17864
rect 4948 17824 4954 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 4985 17827 5043 17833
rect 5460 17836 8217 17864
rect 5460 17796 5488 17836
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 8205 17827 8263 17833
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 8846 17864 8852 17876
rect 8619 17836 8852 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 8846 17824 8852 17836
rect 8904 17824 8910 17876
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9858 17864 9864 17876
rect 9416 17836 9864 17864
rect 1964 17768 2360 17796
rect 2516 17768 5488 17796
rect 7193 17799 7251 17805
rect 1964 17737 1992 17768
rect 2516 17737 2544 17768
rect 7193 17765 7205 17799
rect 7239 17796 7251 17799
rect 7650 17796 7656 17808
rect 7239 17768 7656 17796
rect 7239 17765 7251 17768
rect 7193 17759 7251 17765
rect 7650 17756 7656 17768
rect 7708 17756 7714 17808
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17697 1639 17731
rect 1581 17691 1639 17697
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17697 2007 17731
rect 1949 17691 2007 17697
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17697 2559 17731
rect 2501 17691 2559 17697
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 3053 17731 3111 17737
rect 2823 17700 3004 17728
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 1596 17592 1624 17691
rect 2056 17660 2084 17691
rect 2976 17660 3004 17700
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 3326 17728 3332 17740
rect 3099 17700 3332 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 3476 17700 3521 17728
rect 3476 17688 3482 17700
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 4341 17731 4399 17737
rect 4341 17728 4353 17731
rect 4304 17700 4353 17728
rect 4304 17688 4310 17700
rect 4341 17697 4353 17700
rect 4387 17697 4399 17731
rect 7101 17731 7159 17737
rect 4341 17691 4399 17697
rect 4428 17700 6960 17728
rect 4428 17660 4456 17700
rect 2056 17632 2912 17660
rect 2976 17632 4456 17660
rect 4617 17663 4675 17669
rect 2130 17592 2136 17604
rect 1596 17564 2136 17592
rect 2130 17552 2136 17564
rect 2188 17552 2194 17604
rect 2884 17601 2912 17632
rect 4617 17629 4629 17663
rect 4663 17660 4675 17663
rect 4798 17660 4804 17672
rect 4663 17632 4804 17660
rect 4663 17629 4675 17632
rect 4617 17623 4675 17629
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 5350 17620 5356 17672
rect 5408 17660 5414 17672
rect 6546 17660 6552 17672
rect 5408 17632 6552 17660
rect 5408 17620 5414 17632
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 2225 17595 2283 17601
rect 2225 17561 2237 17595
rect 2271 17592 2283 17595
rect 2869 17595 2927 17601
rect 2271 17564 2774 17592
rect 2271 17561 2283 17564
rect 2225 17555 2283 17561
rect 2746 17524 2774 17564
rect 2869 17561 2881 17595
rect 2915 17561 2927 17595
rect 2869 17555 2927 17561
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 3973 17595 4031 17601
rect 3973 17592 3985 17595
rect 3016 17564 3985 17592
rect 3016 17552 3022 17564
rect 3973 17561 3985 17564
rect 4019 17561 4031 17595
rect 3973 17555 4031 17561
rect 4338 17552 4344 17604
rect 4396 17592 4402 17604
rect 6733 17595 6791 17601
rect 6733 17592 6745 17595
rect 4396 17564 6745 17592
rect 4396 17552 4402 17564
rect 6733 17561 6745 17564
rect 6779 17561 6791 17595
rect 6733 17555 6791 17561
rect 3234 17524 3240 17536
rect 2746 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 5261 17527 5319 17533
rect 5261 17524 5273 17527
rect 4304 17496 5273 17524
rect 4304 17484 4310 17496
rect 5261 17493 5273 17496
rect 5307 17524 5319 17527
rect 5442 17524 5448 17536
rect 5307 17496 5448 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 6932 17524 6960 17700
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7374 17728 7380 17740
rect 7147 17700 7380 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17660 7343 17663
rect 7466 17660 7472 17672
rect 7331 17632 7472 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17629 7619 17663
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 7561 17623 7619 17629
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 7576 17592 7604 17623
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 8849 17663 8907 17669
rect 8849 17629 8861 17663
rect 8895 17660 8907 17663
rect 9416 17660 9444 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 12400 17836 13185 17864
rect 12400 17824 12406 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 13630 17824 13636 17876
rect 13688 17864 13694 17876
rect 13725 17867 13783 17873
rect 13725 17864 13737 17867
rect 13688 17836 13737 17864
rect 13688 17824 13694 17836
rect 13725 17833 13737 17836
rect 13771 17833 13783 17867
rect 13725 17827 13783 17833
rect 9784 17768 10180 17796
rect 9784 17669 9812 17768
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10025 17731 10083 17737
rect 10025 17728 10037 17731
rect 9916 17700 10037 17728
rect 9916 17688 9922 17700
rect 10025 17697 10037 17700
rect 10071 17697 10083 17731
rect 10152 17728 10180 17768
rect 10962 17756 10968 17808
rect 11020 17796 11026 17808
rect 15470 17796 15476 17808
rect 11020 17768 15476 17796
rect 11020 17756 11026 17768
rect 15470 17756 15476 17768
rect 15528 17796 15534 17808
rect 16390 17796 16396 17808
rect 15528 17768 16396 17796
rect 15528 17756 15534 17768
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 10502 17728 10508 17740
rect 10152 17700 10508 17728
rect 10025 17691 10083 17697
rect 10502 17688 10508 17700
rect 10560 17728 10566 17740
rect 12066 17737 12072 17740
rect 12060 17728 12072 17737
rect 10560 17700 11744 17728
rect 12027 17700 12072 17728
rect 10560 17688 10566 17700
rect 11716 17672 11744 17700
rect 12060 17691 12072 17700
rect 12066 17688 12072 17691
rect 12124 17688 12130 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 13412 17700 13553 17728
rect 13412 17688 13418 17700
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 8895 17632 9444 17660
rect 9769 17663 9827 17669
rect 8895 17629 8907 17632
rect 8849 17623 8907 17629
rect 9769 17629 9781 17663
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11756 17632 11805 17660
rect 11756 17620 11762 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 7064 17564 7604 17592
rect 7064 17552 7070 17564
rect 11054 17524 11060 17536
rect 6932 17496 11060 17524
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11974 17524 11980 17536
rect 11195 17496 11980 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1854 17320 1860 17332
rect 1815 17292 1860 17320
rect 1854 17280 1860 17292
rect 1912 17280 1918 17332
rect 2130 17320 2136 17332
rect 2091 17292 2136 17320
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 3326 17320 3332 17332
rect 3287 17292 3332 17320
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 4338 17320 4344 17332
rect 3436 17292 4344 17320
rect 2038 17212 2044 17264
rect 2096 17252 2102 17264
rect 3436 17252 3464 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4798 17320 4804 17332
rect 4759 17292 4804 17320
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7524 17292 7849 17320
rect 7524 17280 7530 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 9858 17320 9864 17332
rect 9447 17292 9864 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 2096 17224 3464 17252
rect 2096 17212 2102 17224
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 1728 17156 2421 17184
rect 1728 17144 1734 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17184 2927 17187
rect 2958 17184 2964 17196
rect 2915 17156 2964 17184
rect 2915 17153 2927 17156
rect 2869 17147 2927 17153
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 2280 17088 2329 17116
rect 2280 17076 2286 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2792 17116 2820 17147
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 4816 17184 4844 17280
rect 7852 17184 7880 17283
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10962 17320 10968 17332
rect 10923 17292 10968 17320
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 12066 17280 12072 17332
rect 12124 17320 12130 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 12124 17292 13093 17320
rect 12124 17280 12130 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 13081 17283 13139 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 9306 17252 9312 17264
rect 9267 17224 9312 17252
rect 9306 17212 9312 17224
rect 9364 17212 9370 17264
rect 4816 17156 5028 17184
rect 7852 17156 8064 17184
rect 2792 17088 2912 17116
rect 2317 17079 2375 17085
rect 1578 17048 1584 17060
rect 1539 17020 1584 17048
rect 1578 17008 1584 17020
rect 1636 17008 1642 17060
rect 1946 17048 1952 17060
rect 1907 17020 1952 17048
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 2884 17048 2912 17088
rect 3050 17076 3056 17128
rect 3108 17116 3114 17128
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 3108 17088 3433 17116
rect 3108 17076 3114 17088
rect 3421 17085 3433 17088
rect 3467 17116 3479 17119
rect 3688 17119 3746 17125
rect 3467 17088 3648 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 3620 17048 3648 17088
rect 3688 17085 3700 17119
rect 3734 17116 3746 17119
rect 3970 17116 3976 17128
rect 3734 17088 3976 17116
rect 3734 17085 3746 17088
rect 3688 17079 3746 17085
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17085 4951 17119
rect 5000 17116 5028 17156
rect 5149 17119 5207 17125
rect 5149 17116 5161 17119
rect 5000 17088 5161 17116
rect 4893 17079 4951 17085
rect 5149 17085 5161 17088
rect 5195 17085 5207 17119
rect 5149 17079 5207 17085
rect 6457 17119 6515 17125
rect 6457 17085 6469 17119
rect 6503 17116 6515 17119
rect 7929 17119 7987 17125
rect 7929 17116 7941 17119
rect 6503 17088 7941 17116
rect 6503 17085 6515 17088
rect 6457 17079 6515 17085
rect 7929 17085 7941 17088
rect 7975 17085 7987 17119
rect 8036 17116 8064 17156
rect 8185 17119 8243 17125
rect 8185 17116 8197 17119
rect 8036 17088 8197 17116
rect 7929 17079 7987 17085
rect 8185 17085 8197 17088
rect 8231 17085 8243 17119
rect 9324 17116 9352 17212
rect 11698 17184 11704 17196
rect 11072 17156 11704 17184
rect 11072 17128 11100 17156
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 21542 17184 21548 17196
rect 21503 17156 21548 17184
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 10502 17116 10508 17128
rect 10560 17125 10566 17128
rect 9324 17088 10508 17116
rect 8185 17079 8243 17085
rect 3786 17048 3792 17060
rect 2884 17020 3464 17048
rect 3620 17020 3792 17048
rect 3436 16992 3464 17020
rect 3786 17008 3792 17020
rect 3844 17048 3850 17060
rect 4908 17048 4936 17079
rect 6362 17048 6368 17060
rect 3844 17020 6368 17048
rect 3844 17008 3850 17020
rect 6362 17008 6368 17020
rect 6420 17048 6426 17060
rect 6472 17048 6500 17079
rect 10502 17076 10508 17088
rect 10560 17079 10572 17125
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 11054 17116 11060 17128
rect 10827 17088 11060 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10560 17076 10566 17079
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11974 17125 11980 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11204 17088 11253 17116
rect 11204 17076 11210 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 11968 17116 11980 17125
rect 11935 17088 11980 17116
rect 11241 17079 11299 17085
rect 11968 17079 11980 17088
rect 11974 17076 11980 17079
rect 12032 17076 12038 17128
rect 13170 17116 13176 17128
rect 13131 17088 13176 17116
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 6420 17020 6500 17048
rect 6724 17051 6782 17057
rect 6420 17008 6426 17020
rect 6724 17017 6736 17051
rect 6770 17048 6782 17051
rect 7098 17048 7104 17060
rect 6770 17020 7104 17048
rect 6770 17017 6782 17020
rect 6724 17011 6782 17017
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 21085 17051 21143 17057
rect 21085 17048 21097 17051
rect 7208 17020 21097 17048
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3016 16952 3061 16980
rect 3016 16940 3022 16952
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 6273 16983 6331 16989
rect 6273 16980 6285 16983
rect 3476 16952 6285 16980
rect 3476 16940 3482 16952
rect 6273 16949 6285 16952
rect 6319 16980 6331 16983
rect 7208 16980 7236 17020
rect 21085 17017 21097 17020
rect 21131 17048 21143 17051
rect 21361 17051 21419 17057
rect 21361 17048 21373 17051
rect 21131 17020 21373 17048
rect 21131 17017 21143 17020
rect 21085 17011 21143 17017
rect 21361 17017 21373 17020
rect 21407 17017 21419 17051
rect 21361 17011 21419 17017
rect 11054 16980 11060 16992
rect 6319 16952 7236 16980
rect 11015 16952 11060 16980
rect 6319 16949 6331 16952
rect 6273 16943 6331 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11330 16980 11336 16992
rect 11291 16952 11336 16980
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 18138 16980 18144 16992
rect 12124 16952 18144 16980
rect 12124 16940 12130 16952
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2222 16776 2228 16788
rect 2183 16748 2228 16776
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2372 16748 2417 16776
rect 2372 16736 2378 16748
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3513 16779 3571 16785
rect 3513 16776 3525 16779
rect 3016 16748 3525 16776
rect 3016 16736 3022 16748
rect 3513 16745 3525 16748
rect 3559 16745 3571 16779
rect 3513 16739 3571 16745
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 7374 16776 7380 16788
rect 5500 16748 7144 16776
rect 7335 16748 7380 16776
rect 5500 16736 5506 16748
rect 2406 16668 2412 16720
rect 2464 16708 2470 16720
rect 2501 16711 2559 16717
rect 2501 16708 2513 16711
rect 2464 16680 2513 16708
rect 2464 16668 2470 16680
rect 2501 16677 2513 16680
rect 2547 16677 2559 16711
rect 3418 16708 3424 16720
rect 3379 16680 3424 16708
rect 2501 16671 2559 16677
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 1670 16640 1676 16652
rect 1627 16612 1676 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 1854 16640 1860 16652
rect 1811 16612 1860 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2038 16640 2044 16652
rect 1999 16612 2044 16640
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2516 16640 2544 16671
rect 3418 16668 3424 16680
rect 3476 16668 3482 16720
rect 4433 16711 4491 16717
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 6822 16708 6828 16720
rect 4479 16680 6828 16708
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 7116 16708 7144 16748
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 7650 16776 7656 16788
rect 7611 16748 7656 16776
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 7760 16748 8524 16776
rect 7760 16708 7788 16748
rect 7116 16680 7788 16708
rect 8021 16711 8079 16717
rect 8021 16677 8033 16711
rect 8067 16708 8079 16711
rect 8067 16680 8432 16708
rect 8067 16677 8079 16680
rect 8021 16671 8079 16677
rect 2958 16640 2964 16652
rect 2516 16612 2964 16640
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 4338 16640 4344 16652
rect 4299 16612 4344 16640
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 5258 16640 5264 16652
rect 4632 16612 5264 16640
rect 4632 16581 4660 16612
rect 5258 16600 5264 16612
rect 5316 16640 5322 16652
rect 5425 16643 5483 16649
rect 5425 16640 5437 16643
rect 5316 16612 5437 16640
rect 5316 16600 5322 16612
rect 5425 16609 5437 16612
rect 5471 16609 5483 16643
rect 6917 16643 6975 16649
rect 6917 16640 6929 16643
rect 5425 16603 5483 16609
rect 6748 16612 6929 16640
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 5184 16504 5212 16535
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 6748 16572 6776 16612
rect 6917 16609 6929 16612
rect 6963 16609 6975 16643
rect 6917 16603 6975 16609
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 8113 16643 8171 16649
rect 7064 16612 7109 16640
rect 7064 16600 7070 16612
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8159 16612 8340 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 6512 16544 6776 16572
rect 6825 16575 6883 16581
rect 6512 16532 6518 16544
rect 6825 16541 6837 16575
rect 6871 16541 6883 16575
rect 6825 16535 6883 16541
rect 8205 16575 8263 16581
rect 8205 16541 8217 16575
rect 8251 16541 8263 16575
rect 8205 16535 8263 16541
rect 3844 16476 5212 16504
rect 6549 16507 6607 16513
rect 3844 16464 3850 16476
rect 6549 16473 6561 16507
rect 6595 16504 6607 16507
rect 6840 16504 6868 16535
rect 7098 16504 7104 16516
rect 6595 16476 7104 16504
rect 6595 16473 6607 16476
rect 6549 16467 6607 16473
rect 7098 16464 7104 16476
rect 7156 16504 7162 16516
rect 8220 16504 8248 16535
rect 7156 16476 8248 16504
rect 7156 16464 7162 16476
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3476 16408 3985 16436
rect 3476 16396 3482 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 8312 16436 8340 16612
rect 8404 16572 8432 16680
rect 8496 16640 8524 16748
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 8720 16748 9781 16776
rect 8720 16736 8726 16748
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 9769 16739 9827 16745
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10962 16776 10968 16788
rect 10183 16748 10968 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 11057 16779 11115 16785
rect 11057 16745 11069 16779
rect 11103 16776 11115 16779
rect 11330 16776 11336 16788
rect 11103 16748 11336 16776
rect 11103 16745 11115 16748
rect 11057 16739 11115 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 11790 16776 11796 16788
rect 11471 16748 11796 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 12253 16779 12311 16785
rect 12253 16776 12265 16779
rect 12216 16748 12265 16776
rect 12216 16736 12222 16748
rect 12253 16745 12265 16748
rect 12299 16745 12311 16779
rect 12253 16739 12311 16745
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 13446 16776 13452 16788
rect 12483 16748 13452 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 8849 16711 8907 16717
rect 8849 16677 8861 16711
rect 8895 16708 8907 16711
rect 11698 16708 11704 16720
rect 8895 16680 11704 16708
rect 8895 16677 8907 16680
rect 8849 16671 8907 16677
rect 11698 16668 11704 16680
rect 11756 16668 11762 16720
rect 11885 16711 11943 16717
rect 11885 16677 11897 16711
rect 11931 16708 11943 16711
rect 12452 16708 12480 16739
rect 13446 16736 13452 16748
rect 13504 16776 13510 16788
rect 14458 16776 14464 16788
rect 13504 16748 14464 16776
rect 13504 16736 13510 16748
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 11931 16680 12480 16708
rect 11931 16677 11943 16680
rect 11885 16671 11943 16677
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 8496 16612 9689 16640
rect 9677 16609 9689 16612
rect 9723 16640 9735 16643
rect 10229 16643 10287 16649
rect 9723 16612 10180 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 8404 16544 8616 16572
rect 8588 16513 8616 16544
rect 8573 16507 8631 16513
rect 8573 16473 8585 16507
rect 8619 16504 8631 16507
rect 8849 16507 8907 16513
rect 8849 16504 8861 16507
rect 8619 16476 8861 16504
rect 8619 16473 8631 16476
rect 8573 16467 8631 16473
rect 8849 16473 8861 16476
rect 8895 16473 8907 16507
rect 10152 16504 10180 16612
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 10778 16640 10784 16652
rect 10275 16612 10784 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 11974 16640 11980 16652
rect 10888 16612 11980 16640
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16572 10471 16575
rect 10502 16572 10508 16584
rect 10459 16544 10508 16572
rect 10459 16541 10471 16544
rect 10413 16535 10471 16541
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 10888 16581 10916 16612
rect 11716 16581 11744 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12084 16612 12633 16640
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16541 10931 16575
rect 10873 16535 10931 16541
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 10965 16535 11023 16541
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16572 11851 16575
rect 11882 16572 11888 16584
rect 11839 16544 11888 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 10980 16504 11008 16535
rect 11882 16532 11888 16544
rect 11940 16572 11946 16584
rect 12084 16572 12112 16612
rect 12621 16609 12633 16612
rect 12667 16640 12679 16643
rect 14550 16640 14556 16652
rect 12667 16612 14556 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 11940 16544 12112 16572
rect 11940 16532 11946 16544
rect 10152 16476 11008 16504
rect 8849 16467 8907 16473
rect 8757 16439 8815 16445
rect 8757 16436 8769 16439
rect 8312 16408 8769 16436
rect 3973 16399 4031 16405
rect 8757 16405 8769 16408
rect 8803 16436 8815 16439
rect 10870 16436 10876 16448
rect 8803 16408 10876 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 13078 16436 13084 16448
rect 11756 16408 13084 16436
rect 11756 16396 11762 16408
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1765 16235 1823 16241
rect 1765 16232 1777 16235
rect 1636 16204 1777 16232
rect 1636 16192 1642 16204
rect 1765 16201 1777 16204
rect 1811 16201 1823 16235
rect 1765 16195 1823 16201
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 2133 16235 2191 16241
rect 2133 16232 2145 16235
rect 1912 16204 2145 16232
rect 1912 16192 1918 16204
rect 2133 16201 2145 16204
rect 2179 16201 2191 16235
rect 5258 16232 5264 16244
rect 5219 16204 5264 16232
rect 2133 16195 2191 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 6420 16204 6745 16232
rect 6420 16192 6426 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 6733 16195 6791 16201
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6880 16204 7941 16232
rect 6880 16192 6886 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9858 16232 9864 16244
rect 9079 16204 9864 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 8478 16096 8484 16108
rect 6196 16068 8484 16096
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 16028 2375 16031
rect 3418 16028 3424 16040
rect 2363 16000 3424 16028
rect 2363 15997 2375 16000
rect 2317 15991 2375 15997
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3786 15988 3792 16040
rect 3844 16028 3850 16040
rect 4154 16037 4160 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3844 16000 3893 16028
rect 3844 15988 3850 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 4148 16028 4160 16037
rect 4067 16000 4160 16028
rect 3881 15991 3939 15997
rect 4148 15991 4160 16000
rect 4212 16028 4218 16040
rect 6196 16028 6224 16068
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 4212 16000 6224 16028
rect 6917 16031 6975 16037
rect 4154 15988 4160 15991
rect 4212 15988 4218 16000
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 7006 16028 7012 16040
rect 6963 16000 7012 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 8389 16031 8447 16037
rect 8389 15997 8401 16031
rect 8435 16028 8447 16031
rect 9048 16028 9076 16195
rect 9858 16192 9864 16204
rect 9916 16232 9922 16244
rect 10410 16232 10416 16244
rect 9916 16204 10416 16232
rect 9916 16192 9922 16204
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 10836 16204 11161 16232
rect 10836 16192 10842 16204
rect 11149 16201 11161 16204
rect 11195 16232 11207 16235
rect 11238 16232 11244 16244
rect 11195 16204 11244 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 13449 16235 13507 16241
rect 13449 16232 13461 16235
rect 13228 16204 13461 16232
rect 13228 16192 13234 16204
rect 13449 16201 13461 16204
rect 13495 16201 13507 16235
rect 13449 16195 13507 16201
rect 11698 16124 11704 16176
rect 11756 16164 11762 16176
rect 13814 16164 13820 16176
rect 11756 16136 13820 16164
rect 11756 16124 11762 16136
rect 13814 16124 13820 16136
rect 13872 16124 13878 16176
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 11422 16096 11428 16108
rect 10459 16068 11428 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 12526 16096 12532 16108
rect 11931 16068 12532 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12526 16056 12532 16068
rect 12584 16056 12590 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 14090 16096 14096 16108
rect 12943 16068 14096 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 11698 16028 11704 16040
rect 8435 16000 9076 16028
rect 10152 16000 11704 16028
rect 8435 15997 8447 16000
rect 8389 15991 8447 15997
rect 1394 15960 1400 15972
rect 1355 15932 1400 15960
rect 1394 15920 1400 15932
rect 1452 15920 1458 15972
rect 1578 15960 1584 15972
rect 1539 15932 1584 15960
rect 1578 15920 1584 15932
rect 1636 15920 1642 15972
rect 8297 15963 8355 15969
rect 8297 15929 8309 15963
rect 8343 15960 8355 15963
rect 8849 15963 8907 15969
rect 8849 15960 8861 15963
rect 8343 15932 8861 15960
rect 8343 15929 8355 15932
rect 8297 15923 8355 15929
rect 8849 15929 8861 15932
rect 8895 15960 8907 15963
rect 10152 15960 10180 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12434 16028 12440 16040
rect 12023 16000 12440 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 13078 16028 13084 16040
rect 13039 16000 13084 16028
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 12069 15963 12127 15969
rect 12069 15960 12081 15963
rect 8895 15932 10180 15960
rect 10980 15932 12081 15960
rect 8895 15929 8907 15932
rect 8849 15923 8907 15929
rect 5718 15852 5724 15904
rect 5776 15892 5782 15904
rect 6454 15892 6460 15904
rect 5776 15864 6460 15892
rect 5776 15852 5782 15864
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 10502 15892 10508 15904
rect 10463 15864 10508 15892
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 10980 15901 11008 15932
rect 12069 15929 12081 15932
rect 12115 15929 12127 15963
rect 14182 15960 14188 15972
rect 12069 15923 12127 15929
rect 12176 15932 14188 15960
rect 10965 15895 11023 15901
rect 10652 15864 10697 15892
rect 10652 15852 10658 15864
rect 10965 15861 10977 15895
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 12176 15892 12204 15932
rect 14182 15920 14188 15932
rect 14240 15920 14246 15972
rect 11296 15864 12204 15892
rect 12437 15895 12495 15901
rect 11296 15852 11302 15864
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12483 15864 13001 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12989 15861 13001 15864
rect 13035 15861 13047 15895
rect 12989 15855 13047 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1578 15648 1584 15700
rect 1636 15688 1642 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1636 15660 1777 15688
rect 1636 15648 1642 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2004 15660 2329 15688
rect 2004 15648 2010 15660
rect 2317 15657 2329 15660
rect 2363 15657 2375 15691
rect 2317 15651 2375 15657
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4396 15660 4721 15688
rect 4396 15648 4402 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 5534 15688 5540 15700
rect 4856 15660 5540 15688
rect 4856 15648 4862 15660
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8478 15688 8484 15700
rect 8159 15660 8484 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 9088 15660 9321 15688
rect 9088 15648 9094 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 3602 15580 3608 15632
rect 3660 15620 3666 15632
rect 4249 15623 4307 15629
rect 4249 15620 4261 15623
rect 3660 15592 4261 15620
rect 3660 15580 3666 15592
rect 4249 15589 4261 15592
rect 4295 15620 4307 15623
rect 5166 15620 5172 15632
rect 4295 15592 5172 15620
rect 4295 15589 4307 15592
rect 4249 15583 4307 15589
rect 5166 15580 5172 15592
rect 5224 15580 5230 15632
rect 6914 15580 6920 15632
rect 6972 15629 6978 15632
rect 6972 15623 7036 15629
rect 6972 15589 6990 15623
rect 7024 15589 7036 15623
rect 9324 15620 9352 15651
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9769 15691 9827 15697
rect 9769 15688 9781 15691
rect 9548 15660 9781 15688
rect 9548 15648 9554 15660
rect 9769 15657 9781 15660
rect 9815 15657 9827 15691
rect 9769 15651 9827 15657
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 9950 15688 9956 15700
rect 9907 15660 9956 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10410 15688 10416 15700
rect 10192 15660 10416 15688
rect 10192 15648 10198 15660
rect 10410 15648 10416 15660
rect 10468 15688 10474 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10468 15660 10793 15688
rect 10468 15648 10474 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 13538 15688 13544 15700
rect 10781 15651 10839 15657
rect 11348 15660 13544 15688
rect 10689 15623 10747 15629
rect 10689 15620 10701 15623
rect 9324 15592 10701 15620
rect 6972 15583 7036 15589
rect 10689 15589 10701 15592
rect 10735 15620 10747 15623
rect 11348 15620 11376 15660
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 10735 15592 11376 15620
rect 10735 15589 10747 15592
rect 10689 15583 10747 15589
rect 6972 15580 6978 15583
rect 11422 15580 11428 15632
rect 11480 15629 11486 15632
rect 11480 15623 11544 15629
rect 11480 15589 11498 15623
rect 11532 15589 11544 15623
rect 14108 15620 14136 15648
rect 14614 15623 14672 15629
rect 14614 15620 14626 15623
rect 11480 15583 11544 15589
rect 12728 15592 13124 15620
rect 14108 15592 14626 15620
rect 11480 15580 11486 15583
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15521 1639 15555
rect 1946 15552 1952 15564
rect 1907 15524 1952 15552
rect 1581 15515 1639 15521
rect 1596 15484 1624 15515
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2222 15552 2228 15564
rect 2183 15524 2228 15552
rect 2222 15512 2228 15524
rect 2280 15512 2286 15564
rect 2501 15555 2559 15561
rect 2501 15521 2513 15555
rect 2547 15552 2559 15555
rect 4154 15552 4160 15564
rect 2547 15524 2774 15552
rect 2547 15521 2559 15524
rect 2501 15515 2559 15521
rect 2038 15484 2044 15496
rect 1596 15456 2044 15484
rect 2038 15444 2044 15456
rect 2096 15444 2102 15496
rect 1394 15416 1400 15428
rect 1355 15388 1400 15416
rect 1394 15376 1400 15388
rect 1452 15376 1458 15428
rect 2746 15416 2774 15524
rect 4080 15524 4160 15552
rect 4080 15493 4108 15524
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4387 15524 4813 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6420 15524 6745 15552
rect 6420 15512 6426 15524
rect 6733 15521 6745 15524
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11112 15524 11253 15552
rect 11112 15512 11118 15524
rect 11241 15521 11253 15524
rect 11287 15552 11299 15555
rect 11790 15552 11796 15564
rect 11287 15524 11796 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 12728 15561 12756 15592
rect 12986 15561 12992 15564
rect 12713 15555 12771 15561
rect 12584 15524 12664 15552
rect 12584 15512 12590 15524
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 9723 15456 10609 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 10597 15453 10609 15456
rect 10643 15484 10655 15487
rect 10962 15484 10968 15496
rect 10643 15456 10968 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 5534 15416 5540 15428
rect 2746 15388 5540 15416
rect 5534 15376 5540 15388
rect 5592 15376 5598 15428
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 2041 15351 2099 15357
rect 2041 15348 2053 15351
rect 1728 15320 2053 15348
rect 1728 15308 1734 15320
rect 2041 15317 2053 15320
rect 2087 15317 2099 15351
rect 2041 15311 2099 15317
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 7374 15348 7380 15360
rect 6236 15320 7380 15348
rect 6236 15308 6242 15320
rect 7374 15308 7380 15320
rect 7432 15348 7438 15360
rect 8202 15348 8208 15360
rect 7432 15320 8208 15348
rect 7432 15308 7438 15320
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 10229 15351 10287 15357
rect 10229 15317 10241 15351
rect 10275 15348 10287 15351
rect 11054 15348 11060 15360
rect 10275 15320 11060 15348
rect 10275 15317 10287 15320
rect 10229 15311 10287 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11149 15351 11207 15357
rect 11149 15317 11161 15351
rect 11195 15348 11207 15351
rect 11974 15348 11980 15360
rect 11195 15320 11980 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12636 15357 12664 15524
rect 12713 15521 12725 15555
rect 12759 15521 12771 15555
rect 12980 15552 12992 15561
rect 12947 15524 12992 15552
rect 12713 15515 12771 15521
rect 12980 15515 12992 15524
rect 12986 15512 12992 15515
rect 13044 15512 13050 15564
rect 13096 15552 13124 15592
rect 14614 15589 14626 15592
rect 14660 15589 14672 15623
rect 14614 15583 14672 15589
rect 13096 15524 14412 15552
rect 14384 15496 14412 15524
rect 14366 15484 14372 15496
rect 14327 15456 14372 15484
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 12621 15351 12679 15357
rect 12621 15317 12633 15351
rect 12667 15348 12679 15351
rect 12986 15348 12992 15360
rect 12667 15320 12992 15348
rect 12667 15317 12679 15320
rect 12621 15311 12679 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 15746 15348 15752 15360
rect 15707 15320 15752 15348
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2041 15147 2099 15153
rect 2041 15144 2053 15147
rect 2004 15116 2053 15144
rect 2004 15104 2010 15116
rect 2041 15113 2053 15116
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 2317 15147 2375 15153
rect 2317 15144 2329 15147
rect 2280 15116 2329 15144
rect 2280 15104 2286 15116
rect 2317 15113 2329 15116
rect 2363 15113 2375 15147
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 2317 15107 2375 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6457 15147 6515 15153
rect 6457 15113 6469 15147
rect 6503 15144 6515 15147
rect 6822 15144 6828 15156
rect 6503 15116 6828 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7558 15144 7564 15156
rect 6932 15116 7564 15144
rect 3694 15036 3700 15088
rect 3752 15076 3758 15088
rect 4249 15079 4307 15085
rect 4249 15076 4261 15079
rect 3752 15048 4261 15076
rect 3752 15036 3758 15048
rect 4249 15045 4261 15048
rect 4295 15076 4307 15079
rect 6932 15076 6960 15116
rect 7558 15104 7564 15116
rect 7616 15104 7622 15156
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 10594 15144 10600 15156
rect 9815 15116 10600 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11238 15144 11244 15156
rect 11199 15116 11244 15144
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12492 15116 12537 15144
rect 12492 15104 12498 15116
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 13136 15116 13369 15144
rect 13136 15104 13142 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 4295 15048 6960 15076
rect 4295 15045 4307 15048
rect 4249 15039 4307 15045
rect 1394 15008 1400 15020
rect 1355 14980 1400 15008
rect 1394 14968 1400 14980
rect 1452 14968 1458 15020
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 15008 6239 15011
rect 6822 15008 6828 15020
rect 6227 14980 6828 15008
rect 6227 14977 6239 14980
rect 6181 14971 6239 14977
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 7944 14980 8493 15008
rect 2225 14943 2283 14949
rect 2225 14909 2237 14943
rect 2271 14909 2283 14943
rect 2225 14903 2283 14909
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14909 2559 14943
rect 2501 14903 2559 14909
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14940 2743 14943
rect 3786 14940 3792 14952
rect 2731 14912 3792 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 1762 14872 1768 14884
rect 1627 14844 1768 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 1762 14832 1768 14844
rect 1820 14832 1826 14884
rect 2240 14804 2268 14903
rect 2516 14872 2544 14903
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 6420 14912 7849 14940
rect 6420 14900 6426 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 2774 14872 2780 14884
rect 2516 14844 2780 14872
rect 2774 14832 2780 14844
rect 2832 14832 2838 14884
rect 2952 14875 3010 14881
rect 2952 14841 2964 14875
rect 2998 14872 3010 14875
rect 3050 14872 3056 14884
rect 2998 14844 3056 14872
rect 2998 14841 3010 14844
rect 2952 14835 3010 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 5905 14875 5963 14881
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 5951 14844 6960 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 3786 14804 3792 14816
rect 2240 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4062 14804 4068 14816
rect 4023 14776 4068 14804
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 5994 14804 6000 14816
rect 5955 14776 6000 14804
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6932 14804 6960 14844
rect 7466 14832 7472 14884
rect 7524 14872 7530 14884
rect 7570 14875 7628 14881
rect 7570 14872 7582 14875
rect 7524 14844 7582 14872
rect 7524 14832 7530 14844
rect 7570 14841 7582 14844
rect 7616 14872 7628 14875
rect 7944 14872 7972 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 15008 9275 15011
rect 11256 15008 11284 15104
rect 12250 15076 12256 15088
rect 11808 15048 12256 15076
rect 11808 15017 11836 15048
rect 12250 15036 12256 15048
rect 12308 15076 12314 15088
rect 12308 15048 12572 15076
rect 12308 15036 12314 15048
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 9263 14980 9996 15008
rect 11256 14980 11805 15008
rect 9263 14977 9275 14980
rect 9217 14971 9275 14977
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 8260 14912 8401 14940
rect 8260 14900 8266 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9180 14912 9321 14940
rect 9180 14900 9186 14912
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 9674 14940 9680 14952
rect 9447 14912 9680 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 7616 14844 7972 14872
rect 9324 14872 9352 14903
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 9968 14940 9996 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11974 15008 11980 15020
rect 11935 14980 11980 15008
rect 11793 14971 11851 14977
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12544 15008 12572 15048
rect 13170 15036 13176 15088
rect 13228 15076 13234 15088
rect 19058 15076 19064 15088
rect 13228 15048 19064 15076
rect 13228 15036 13234 15048
rect 19058 15036 19064 15048
rect 19116 15036 19122 15088
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 12544 14980 12633 15008
rect 12621 14977 12633 14980
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13044 14980 13921 15008
rect 13044 14968 13050 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 14461 15011 14519 15017
rect 14461 14977 14473 15011
rect 14507 15008 14519 15011
rect 15194 15008 15200 15020
rect 14507 14980 15200 15008
rect 14507 14977 14519 14980
rect 14461 14971 14519 14977
rect 15194 14968 15200 14980
rect 15252 15008 15258 15020
rect 15746 15008 15752 15020
rect 15252 14980 15752 15008
rect 15252 14968 15258 14980
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 9968 14912 10171 14940
rect 9861 14903 9919 14909
rect 9582 14872 9588 14884
rect 9324 14844 9588 14872
rect 7616 14841 7628 14844
rect 7570 14835 7628 14841
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 6932 14776 7941 14804
rect 7929 14773 7941 14776
rect 7975 14773 7987 14807
rect 8294 14804 8300 14816
rect 8255 14776 8300 14804
rect 7929 14767 7987 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 9876 14804 9904 14903
rect 10143 14881 10171 14912
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 12069 14943 12127 14949
rect 12069 14940 12081 14943
rect 11112 14912 12081 14940
rect 11112 14900 11118 14912
rect 12069 14909 12081 14912
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 14553 14943 14611 14949
rect 14553 14940 14565 14943
rect 13596 14912 14565 14940
rect 13596 14900 13602 14912
rect 14553 14909 14565 14912
rect 14599 14940 14611 14943
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14599 14912 15117 14940
rect 14599 14909 14611 14912
rect 14553 14903 14611 14909
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15105 14903 15163 14909
rect 10128 14875 10186 14881
rect 10128 14841 10140 14875
rect 10174 14872 10186 14875
rect 10962 14872 10968 14884
rect 10174 14844 10968 14872
rect 10174 14841 10186 14844
rect 10128 14835 10186 14841
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 12802 14872 12808 14884
rect 12763 14844 12808 14872
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 13280 14844 13829 14872
rect 11790 14804 11796 14816
rect 9876 14776 11796 14804
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 13280 14813 13308 14844
rect 13817 14841 13829 14844
rect 13863 14841 13875 14875
rect 13817 14835 13875 14841
rect 13265 14807 13323 14813
rect 12952 14776 12997 14804
rect 12952 14764 12958 14776
rect 13265 14773 13277 14807
rect 13311 14773 13323 14807
rect 13722 14804 13728 14816
rect 13683 14776 13728 14804
rect 13265 14767 13323 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15013 14807 15071 14813
rect 15013 14804 15025 14807
rect 14792 14776 15025 14804
rect 14792 14764 14798 14776
rect 15013 14773 15025 14776
rect 15059 14773 15071 14807
rect 15013 14767 15071 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1762 14600 1768 14612
rect 1723 14572 1768 14600
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 2038 14600 2044 14612
rect 1999 14572 2044 14600
rect 2038 14560 2044 14572
rect 2096 14560 2102 14612
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3200 14572 3249 14600
rect 3200 14560 3206 14572
rect 3237 14569 3249 14572
rect 3283 14600 3295 14603
rect 3694 14600 3700 14612
rect 3283 14572 3700 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 5994 14560 6000 14612
rect 6052 14600 6058 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 6052 14572 7297 14600
rect 6052 14560 6058 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 7745 14603 7803 14609
rect 7745 14569 7757 14603
rect 7791 14600 7803 14603
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7791 14572 8217 14600
rect 7791 14569 7803 14572
rect 7745 14563 7803 14569
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 8665 14603 8723 14609
rect 8665 14569 8677 14603
rect 8711 14600 8723 14603
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 8711 14572 9689 14600
rect 8711 14569 8723 14572
rect 8665 14563 8723 14569
rect 9677 14569 9689 14572
rect 9723 14600 9735 14603
rect 9766 14600 9772 14612
rect 9723 14572 9772 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10502 14600 10508 14612
rect 10459 14572 10508 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10744 14572 10885 14600
rect 10744 14560 10750 14572
rect 10873 14569 10885 14572
rect 10919 14600 10931 14603
rect 11054 14600 11060 14612
rect 10919 14572 11060 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11204 14572 11437 14600
rect 11204 14560 11210 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13081 14603 13139 14609
rect 13081 14600 13093 14603
rect 12860 14572 13093 14600
rect 12860 14560 12866 14572
rect 13081 14569 13093 14572
rect 13127 14569 13139 14603
rect 13081 14563 13139 14569
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13320 14572 13461 14600
rect 13320 14560 13326 14572
rect 13449 14569 13461 14572
rect 13495 14600 13507 14603
rect 15286 14600 15292 14612
rect 13495 14572 15292 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 4062 14492 4068 14544
rect 4120 14541 4126 14544
rect 4120 14535 4184 14541
rect 4120 14501 4138 14535
rect 4172 14501 4184 14535
rect 4120 14495 4184 14501
rect 7101 14535 7159 14541
rect 7101 14501 7113 14535
rect 7147 14532 7159 14535
rect 8294 14532 8300 14544
rect 7147 14504 8300 14532
rect 7147 14501 7159 14504
rect 7101 14495 7159 14501
rect 4120 14492 4126 14495
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 10134 14532 10140 14544
rect 9324 14504 10140 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14433 1639 14467
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1581 14427 1639 14433
rect 1596 14396 1624 14427
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2222 14464 2228 14476
rect 2183 14436 2228 14464
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14464 3387 14467
rect 3694 14464 3700 14476
rect 3375 14436 3700 14464
rect 3375 14433 3387 14436
rect 3329 14427 3387 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14464 3939 14467
rect 5620 14467 5678 14473
rect 5620 14464 5632 14467
rect 3927 14436 5212 14464
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 2314 14396 2320 14408
rect 1596 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3068 14328 3096 14356
rect 3068 14300 3924 14328
rect 2777 14263 2835 14269
rect 2777 14229 2789 14263
rect 2823 14260 2835 14263
rect 2866 14260 2872 14272
rect 2823 14232 2872 14260
rect 2823 14229 2835 14232
rect 2777 14223 2835 14229
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3697 14263 3755 14269
rect 3697 14260 3709 14263
rect 3568 14232 3709 14260
rect 3568 14220 3574 14232
rect 3697 14229 3709 14232
rect 3743 14229 3755 14263
rect 3896 14260 3924 14300
rect 4246 14260 4252 14272
rect 3896 14232 4252 14260
rect 3697 14223 3755 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 5184 14260 5212 14436
rect 5276 14436 5632 14464
rect 5276 14337 5304 14436
rect 5620 14433 5632 14436
rect 5666 14464 5678 14467
rect 5666 14436 6592 14464
rect 5666 14433 5678 14436
rect 5620 14427 5678 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14365 5411 14399
rect 5353 14359 5411 14365
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 5261 14291 5319 14297
rect 5368 14260 5396 14359
rect 6564 14328 6592 14436
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 9324 14473 9352 14504
rect 10134 14492 10140 14504
rect 10192 14532 10198 14544
rect 12621 14535 12679 14541
rect 10192 14504 11284 14532
rect 10192 14492 10198 14504
rect 7653 14467 7711 14473
rect 7653 14464 7665 14467
rect 7616 14436 7665 14464
rect 7616 14424 7622 14436
rect 7653 14433 7665 14436
rect 7699 14433 7711 14467
rect 7653 14427 7711 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 9309 14467 9367 14473
rect 8619 14436 9076 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 7466 14396 7472 14408
rect 7239 14368 7472 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 7466 14356 7472 14368
rect 7524 14396 7530 14408
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 7524 14368 7849 14396
rect 7524 14356 7530 14368
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 8772 14328 8800 14359
rect 6564 14300 8800 14328
rect 9048 14328 9076 14436
rect 9309 14433 9321 14467
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 10042 14464 10048 14476
rect 9732 14436 10048 14464
rect 9732 14424 9738 14436
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10778 14464 10784 14476
rect 10284 14436 10784 14464
rect 10284 14424 10290 14436
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 11256 14473 11284 14504
rect 12621 14501 12633 14535
rect 12667 14532 12679 14535
rect 13909 14535 13967 14541
rect 13909 14532 13921 14535
rect 12667 14504 13921 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 13909 14501 13921 14504
rect 13955 14501 13967 14535
rect 13909 14495 13967 14501
rect 14728 14535 14786 14541
rect 14728 14501 14740 14535
rect 14774 14532 14786 14535
rect 15194 14532 15200 14544
rect 14774 14504 15200 14532
rect 14774 14501 14786 14504
rect 14728 14495 14786 14501
rect 15194 14492 15200 14504
rect 15252 14492 15258 14544
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 13541 14467 13599 14473
rect 11241 14427 11299 14433
rect 11624 14436 13400 14464
rect 9214 14356 9220 14408
rect 9272 14396 9278 14408
rect 10686 14396 10692 14408
rect 9272 14368 10692 14396
rect 9272 14356 9278 14368
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11624 14396 11652 14436
rect 13372 14408 13400 14436
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14090 14464 14096 14476
rect 13587 14436 14096 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 11112 14368 11652 14396
rect 11112 14356 11118 14368
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 12308 14368 12357 14396
rect 12308 14356 12314 14368
rect 12345 14365 12357 14368
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 13078 14396 13084 14408
rect 12575 14368 13084 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13412 14368 13645 14396
rect 13412 14356 13418 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14366 14396 14372 14408
rect 13872 14368 14372 14396
rect 13872 14356 13878 14368
rect 14366 14356 14372 14368
rect 14424 14396 14430 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14424 14368 14473 14396
rect 14424 14356 14430 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 9490 14328 9496 14340
rect 9048 14300 9496 14328
rect 9490 14288 9496 14300
rect 9548 14328 9554 14340
rect 12066 14328 12072 14340
rect 9548 14300 12072 14328
rect 9548 14288 9554 14300
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 12989 14331 13047 14337
rect 12989 14297 13001 14331
rect 13035 14328 13047 14331
rect 13722 14328 13728 14340
rect 13035 14300 13728 14328
rect 13035 14297 13047 14300
rect 12989 14291 13047 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 5534 14260 5540 14272
rect 5184 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6733 14263 6791 14269
rect 6733 14229 6745 14263
rect 6779 14260 6791 14263
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 6779 14232 7205 14260
rect 6779 14229 6791 14232
rect 6733 14223 6791 14229
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 9125 14263 9183 14269
rect 9125 14260 9137 14263
rect 7340 14232 9137 14260
rect 7340 14220 7346 14232
rect 9125 14229 9137 14232
rect 9171 14229 9183 14263
rect 9125 14223 9183 14229
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 11882 14260 11888 14272
rect 9824 14232 11888 14260
rect 9824 14220 9830 14232
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 12161 14263 12219 14269
rect 12161 14229 12173 14263
rect 12207 14260 12219 14263
rect 12342 14260 12348 14272
rect 12207 14232 12348 14260
rect 12207 14229 12219 14232
rect 12161 14223 12219 14229
rect 12342 14220 12348 14232
rect 12400 14260 12406 14272
rect 13262 14260 13268 14272
rect 12400 14232 13268 14260
rect 12400 14220 12406 14232
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 15841 14263 15899 14269
rect 15841 14260 15853 14263
rect 15712 14232 15853 14260
rect 15712 14220 15718 14232
rect 15841 14229 15853 14232
rect 15887 14229 15899 14263
rect 15841 14223 15899 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1486 14056 1492 14068
rect 1447 14028 1492 14056
rect 1486 14016 1492 14028
rect 1544 14016 1550 14068
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2004 14028 2605 14056
rect 2004 14016 2010 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 2832 14028 3157 14056
rect 2832 14016 2838 14028
rect 3145 14025 3157 14028
rect 3191 14025 3203 14059
rect 10962 14056 10968 14068
rect 3145 14019 3203 14025
rect 3528 14028 10968 14056
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13957 2099 13991
rect 2314 13988 2320 14000
rect 2275 13960 2320 13988
rect 2041 13951 2099 13957
rect 2056 13920 2084 13951
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13988 3111 13991
rect 3528 13988 3556 14028
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11793 14059 11851 14065
rect 11793 14025 11805 14059
rect 11839 14056 11851 14059
rect 12434 14056 12440 14068
rect 11839 14028 12440 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12618 14056 12624 14068
rect 12579 14028 12624 14056
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 12894 14056 12900 14068
rect 12759 14028 12900 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 4709 13991 4767 13997
rect 4709 13988 4721 13991
rect 3099 13960 3556 13988
rect 3620 13960 4721 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 3620 13929 3648 13960
rect 4709 13957 4721 13960
rect 4755 13957 4767 13991
rect 4709 13951 4767 13957
rect 7466 13948 7472 14000
rect 7524 13988 7530 14000
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 7524 13960 7849 13988
rect 7524 13948 7530 13960
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 9674 13988 9680 14000
rect 7837 13951 7895 13957
rect 9232 13960 9680 13988
rect 1596 13892 2084 13920
rect 3605 13923 3663 13929
rect 1596 13861 1624 13892
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 4062 13920 4068 13932
rect 3835 13892 4068 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4304 13892 5273 13920
rect 4304 13880 4310 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7650 13920 7656 13932
rect 7055 13892 7656 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 9232 13929 9260 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 11992 13960 13584 13988
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9364 13892 9781 13920
rect 9364 13880 9370 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10226 13920 10232 13932
rect 9999 13892 10232 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10284 13892 11100 13920
rect 10284 13880 10290 13892
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1581 13815 1639 13821
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2096 13824 2237 13852
rect 2096 13812 2102 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2406 13812 2412 13864
rect 2464 13852 2470 13864
rect 2501 13855 2559 13861
rect 2501 13852 2513 13855
rect 2464 13824 2513 13852
rect 2464 13812 2470 13824
rect 2501 13821 2513 13824
rect 2547 13821 2559 13855
rect 2501 13815 2559 13821
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2792 13784 2820 13815
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3510 13852 3516 13864
rect 2924 13824 2969 13852
rect 3471 13824 3516 13852
rect 2924 13812 2930 13824
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3694 13812 3700 13864
rect 3752 13852 3758 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3752 13824 3985 13852
rect 3752 13812 3758 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5994 13852 6000 13864
rect 5215 13824 6000 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 7098 13852 7104 13864
rect 7059 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13852 7803 13855
rect 8386 13852 8392 13864
rect 7791 13824 8392 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 2792 13756 5212 13784
rect 5184 13728 5212 13756
rect 6362 13744 6368 13796
rect 6420 13784 6426 13796
rect 7760 13784 7788 13815
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 10318 13852 10324 13864
rect 8496 13824 10324 13852
rect 6420 13756 7788 13784
rect 6420 13744 6426 13756
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 5074 13716 5080 13728
rect 5035 13688 5080 13716
rect 5074 13676 5080 13688
rect 5132 13676 5138 13728
rect 5166 13676 5172 13728
rect 5224 13676 5230 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7561 13719 7619 13725
rect 7248 13688 7293 13716
rect 7248 13676 7254 13688
rect 7561 13685 7573 13719
rect 7607 13716 7619 13719
rect 8496 13716 8524 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 8972 13787 9030 13793
rect 8972 13784 8984 13787
rect 8628 13756 8984 13784
rect 8628 13744 8634 13756
rect 8972 13753 8984 13756
rect 9018 13784 9030 13787
rect 9214 13784 9220 13796
rect 9018 13756 9220 13784
rect 9018 13753 9030 13756
rect 8972 13747 9030 13753
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13753 9735 13787
rect 11072 13784 11100 13892
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11992 13920 12020 13960
rect 11204 13892 12020 13920
rect 12069 13923 12127 13929
rect 11204 13880 11210 13892
rect 12069 13889 12081 13923
rect 12115 13920 12127 13923
rect 12802 13920 12808 13932
rect 12115 13892 12808 13920
rect 12115 13889 12127 13892
rect 12069 13883 12127 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13170 13920 13176 13932
rect 13131 13892 13176 13920
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 13354 13920 13360 13932
rect 13315 13892 13360 13920
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13852 11575 13855
rect 11698 13852 11704 13864
rect 11563 13824 11704 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 11698 13812 11704 13824
rect 11756 13852 11762 13864
rect 13188 13852 13216 13880
rect 13556 13861 13584 13960
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 15105 13923 15163 13929
rect 15105 13920 15117 13923
rect 14792 13892 15117 13920
rect 14792 13880 14798 13892
rect 15105 13889 15117 13892
rect 15151 13889 15163 13923
rect 15105 13883 15163 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15654 13920 15660 13932
rect 15335 13892 15660 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 11756 13824 13216 13852
rect 13541 13855 13599 13861
rect 11756 13812 11762 13824
rect 13541 13821 13553 13855
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 14090 13812 14096 13864
rect 14148 13852 14154 13864
rect 21358 13852 21364 13864
rect 14148 13824 21364 13852
rect 14148 13812 14154 13824
rect 15028 13793 15056 13824
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 15013 13787 15071 13793
rect 11072 13756 13584 13784
rect 9677 13747 9735 13753
rect 9306 13716 9312 13728
rect 7607 13688 8524 13716
rect 9267 13688 9312 13716
rect 7607 13685 7619 13688
rect 7561 13679 7619 13685
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9692 13716 9720 13747
rect 13556 13728 13584 13756
rect 15013 13753 15025 13787
rect 15059 13753 15071 13787
rect 15013 13747 15071 13753
rect 12158 13716 12164 13728
rect 9640 13688 9720 13716
rect 12119 13688 12164 13716
rect 9640 13676 9646 13688
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12253 13719 12311 13725
rect 12253 13685 12265 13719
rect 12299 13716 12311 13719
rect 12526 13716 12532 13728
rect 12299 13688 12532 13716
rect 12299 13685 12311 13688
rect 12253 13679 12311 13685
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 13081 13719 13139 13725
rect 13081 13716 13093 13719
rect 12676 13688 13093 13716
rect 12676 13676 12682 13688
rect 13081 13685 13093 13688
rect 13127 13716 13139 13719
rect 13262 13716 13268 13728
rect 13127 13688 13268 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 13538 13676 13544 13728
rect 13596 13676 13602 13728
rect 13722 13716 13728 13728
rect 13683 13688 13728 13716
rect 13722 13676 13728 13688
rect 13780 13676 13786 13728
rect 14642 13716 14648 13728
rect 14603 13688 14648 13716
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 1486 13512 1492 13524
rect 1447 13484 1492 13512
rect 1486 13472 1492 13484
rect 1544 13472 1550 13524
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2455 13484 2881 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4304 13484 4537 13512
rect 4304 13472 4310 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 5994 13512 6000 13524
rect 5955 13484 6000 13512
rect 4525 13475 4583 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6825 13515 6883 13521
rect 6825 13481 6837 13515
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 7883 13484 8217 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8662 13512 8668 13524
rect 8575 13484 8668 13512
rect 8205 13475 8263 13481
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 1762 13444 1768 13456
rect 1627 13416 1768 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 1762 13404 1768 13416
rect 1820 13404 1826 13456
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 6454 13444 6460 13456
rect 5592 13416 6460 13444
rect 5592 13404 5598 13416
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 3234 13376 3240 13388
rect 3195 13348 3240 13376
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 5626 13336 5632 13388
rect 5684 13385 5690 13388
rect 5920 13385 5948 13416
rect 6454 13404 6460 13416
rect 6512 13444 6518 13456
rect 6840 13444 6868 13475
rect 8662 13472 8668 13484
rect 8720 13512 8726 13524
rect 9030 13512 9036 13524
rect 8720 13484 9036 13512
rect 8720 13472 8726 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9585 13515 9643 13521
rect 9585 13481 9597 13515
rect 9631 13512 9643 13515
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 9631 13484 12909 13512
rect 9631 13481 9643 13484
rect 9585 13475 9643 13481
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 13228 13484 13277 13512
rect 13228 13472 13234 13484
rect 13265 13481 13277 13484
rect 13311 13512 13323 13515
rect 13630 13512 13636 13524
rect 13311 13484 13636 13512
rect 13311 13481 13323 13484
rect 13265 13475 13323 13481
rect 13630 13472 13636 13484
rect 13688 13512 13694 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13688 13484 13737 13512
rect 13688 13472 13694 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14700 13484 14841 13512
rect 14700 13472 14706 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 15562 13512 15568 13524
rect 15523 13484 15568 13512
rect 14829 13475 14887 13481
rect 15562 13472 15568 13484
rect 15620 13512 15626 13524
rect 16298 13512 16304 13524
rect 15620 13484 16304 13512
rect 15620 13472 15626 13484
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 6914 13444 6920 13456
rect 6512 13416 6920 13444
rect 6512 13404 6518 13416
rect 6914 13404 6920 13416
rect 6972 13444 6978 13456
rect 7745 13447 7803 13453
rect 6972 13416 7696 13444
rect 6972 13404 6978 13416
rect 5684 13376 5696 13385
rect 5905 13379 5963 13385
rect 5684 13348 5729 13376
rect 5684 13339 5696 13348
rect 5905 13345 5917 13379
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 6822 13376 6828 13388
rect 6411 13348 6828 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 5684 13336 5690 13339
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7006 13376 7012 13388
rect 6967 13348 7012 13376
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7668 13376 7696 13416
rect 7745 13413 7757 13447
rect 7791 13444 7803 13447
rect 9306 13444 9312 13456
rect 7791 13416 9312 13444
rect 7791 13413 7803 13416
rect 7745 13407 7803 13413
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 9490 13444 9496 13456
rect 9451 13416 9496 13444
rect 9490 13404 9496 13416
rect 9548 13444 9554 13456
rect 10226 13444 10232 13456
rect 9548 13416 10232 13444
rect 9548 13404 9554 13416
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 11790 13444 11796 13456
rect 11440 13416 11796 13444
rect 7834 13376 7840 13388
rect 7668 13348 7840 13376
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 9214 13376 9220 13388
rect 8619 13348 9220 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 9214 13336 9220 13348
rect 9272 13376 9278 13388
rect 9398 13376 9404 13388
rect 9272 13348 9404 13376
rect 9272 13336 9278 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9950 13376 9956 13388
rect 9911 13348 9956 13376
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 11440 13385 11468 13416
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 15470 13404 15476 13456
rect 15528 13444 15534 13456
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 15528 13416 15669 13444
rect 15528 13404 15534 13416
rect 15657 13413 15669 13416
rect 15703 13444 15715 13447
rect 16206 13444 16212 13456
rect 15703 13416 16212 13444
rect 15703 13413 15715 13416
rect 15657 13407 15715 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 11692 13379 11750 13385
rect 11692 13345 11704 13379
rect 11738 13376 11750 13379
rect 12066 13376 12072 13388
rect 11738 13348 12072 13376
rect 11738 13345 11750 13348
rect 11692 13339 11750 13345
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 14090 13376 14096 13388
rect 13403 13348 14096 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15838 13376 15844 13388
rect 14967 13348 15844 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 3326 13308 3332 13320
rect 3287 13280 3332 13308
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 2682 13200 2688 13252
rect 2740 13240 2746 13252
rect 3436 13240 3464 13271
rect 2740 13212 3464 13240
rect 2740 13200 2746 13212
rect 5994 13200 6000 13252
rect 6052 13240 6058 13252
rect 6362 13240 6368 13252
rect 6052 13212 6368 13240
rect 6052 13200 6058 13212
rect 6362 13200 6368 13212
rect 6420 13240 6426 13252
rect 6472 13240 6500 13271
rect 6420 13212 6500 13240
rect 6420 13200 6426 13212
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 1765 13175 1823 13181
rect 1765 13172 1777 13175
rect 1452 13144 1777 13172
rect 1452 13132 1458 13144
rect 1765 13141 1777 13144
rect 1811 13141 1823 13175
rect 1765 13135 1823 13141
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 1949 13175 2007 13181
rect 1949 13172 1961 13175
rect 1912 13144 1961 13172
rect 1912 13132 1918 13144
rect 1949 13141 1961 13144
rect 1995 13141 2007 13175
rect 1949 13135 2007 13141
rect 5626 13132 5632 13184
rect 5684 13172 5690 13184
rect 6564 13172 6592 13271
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7524 13280 7941 13308
rect 7524 13268 7530 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 7193 13243 7251 13249
rect 7193 13240 7205 13243
rect 6880 13212 7205 13240
rect 6880 13200 6886 13212
rect 7193 13209 7205 13212
rect 7239 13240 7251 13243
rect 7944 13240 7972 13271
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8536 13280 8769 13308
rect 8536 13268 8542 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8757 13271 8815 13277
rect 8864 13280 9689 13308
rect 8864 13240 8892 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 9677 13271 9735 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14642 13308 14648 13320
rect 14603 13280 14648 13308
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 10134 13240 10140 13252
rect 7239 13212 7880 13240
rect 7944 13212 8892 13240
rect 8956 13212 9352 13240
rect 10095 13212 10140 13240
rect 7239 13209 7251 13212
rect 7193 13203 7251 13209
rect 7374 13172 7380 13184
rect 5684 13144 6592 13172
rect 7335 13144 7380 13172
rect 5684 13132 5690 13144
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7852 13172 7880 13212
rect 8956 13172 8984 13212
rect 9324 13184 9352 13212
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 12802 13240 12808 13252
rect 10284 13212 10329 13240
rect 12763 13212 12808 13240
rect 10284 13200 10290 13212
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 17954 13240 17960 13252
rect 15120 13212 17960 13240
rect 9122 13172 9128 13184
rect 7852 13144 8984 13172
rect 9083 13144 9128 13172
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 15120 13172 15148 13212
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 15286 13172 15292 13184
rect 9364 13144 15148 13172
rect 15247 13144 15292 13172
rect 9364 13132 9370 13144
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1397 12971 1455 12977
rect 1397 12937 1409 12971
rect 1443 12968 1455 12971
rect 2498 12968 2504 12980
rect 1443 12940 2504 12968
rect 1443 12937 1455 12940
rect 1397 12931 1455 12937
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 4798 12968 4804 12980
rect 4479 12940 4804 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3418 12832 3424 12844
rect 2823 12804 3424 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 2924 12736 3157 12764
rect 2924 12724 2930 12736
rect 3145 12733 3157 12736
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 3973 12767 4031 12773
rect 3973 12764 3985 12767
rect 3936 12736 3985 12764
rect 3936 12724 3942 12736
rect 3973 12733 3985 12736
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 2532 12699 2590 12705
rect 2532 12665 2544 12699
rect 2578 12696 2590 12699
rect 2682 12696 2688 12708
rect 2578 12668 2688 12696
rect 2578 12665 2590 12668
rect 2532 12659 2590 12665
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 3050 12628 3056 12640
rect 3011 12600 3056 12628
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4448 12628 4476 12931
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7708 12940 7849 12968
rect 7708 12928 7714 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 7837 12931 7895 12937
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10502 12968 10508 12980
rect 10275 12940 10508 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 6454 12832 6460 12844
rect 6415 12804 6460 12832
rect 6454 12792 6460 12804
rect 6512 12792 6518 12844
rect 7852 12832 7880 12931
rect 10502 12928 10508 12940
rect 10560 12968 10566 12980
rect 11974 12968 11980 12980
rect 10560 12940 11980 12968
rect 10560 12928 10566 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 15838 12968 15844 12980
rect 13596 12940 15332 12968
rect 15799 12940 15844 12968
rect 13596 12928 13602 12940
rect 12268 12900 12296 12928
rect 8956 12872 12296 12900
rect 15304 12900 15332 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16945 12903 17003 12909
rect 16945 12900 16957 12903
rect 15304 12872 16957 12900
rect 7852 12804 8064 12832
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 8036 12764 8064 12804
rect 8185 12767 8243 12773
rect 8185 12764 8197 12767
rect 8036 12736 8197 12764
rect 7929 12727 7987 12733
rect 8185 12733 8197 12736
rect 8231 12733 8243 12767
rect 8185 12727 8243 12733
rect 6730 12705 6736 12708
rect 6724 12659 6736 12705
rect 6788 12696 6794 12708
rect 6788 12668 6824 12696
rect 6730 12656 6736 12659
rect 6788 12656 6794 12668
rect 8956 12628 8984 12872
rect 16945 12869 16957 12872
rect 16991 12869 17003 12903
rect 16945 12863 17003 12869
rect 9490 12832 9496 12844
rect 9451 12804 9496 12832
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9723 12804 10241 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10686 12832 10692 12844
rect 10551 12804 10692 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11848 12804 12265 12832
rect 11848 12792 11854 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 15654 12792 15660 12844
rect 15712 12832 15718 12844
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 15712 12804 16405 12832
rect 15712 12792 15718 12804
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 9858 12764 9864 12776
rect 9815 12736 9864 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 9858 12724 9864 12736
rect 9916 12764 9922 12776
rect 10042 12764 10048 12776
rect 9916 12736 10048 12764
rect 9916 12724 9922 12736
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 12520 12767 12578 12773
rect 12520 12733 12532 12767
rect 12566 12764 12578 12767
rect 12802 12764 12808 12776
rect 12566 12736 12808 12764
rect 12566 12733 12578 12736
rect 12520 12727 12578 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 13780 12736 14381 12764
rect 13780 12724 13786 12736
rect 14369 12733 14381 12736
rect 14415 12764 14427 12767
rect 16482 12764 16488 12776
rect 14415 12736 16488 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 16482 12724 16488 12736
rect 16540 12764 16546 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 16540 12736 18337 12764
rect 16540 12724 16546 12736
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 9398 12656 9404 12708
rect 9456 12696 9462 12708
rect 14090 12696 14096 12708
rect 9456 12668 14096 12696
rect 9456 12656 9462 12668
rect 14090 12656 14096 12668
rect 14148 12656 14154 12708
rect 14642 12705 14648 12708
rect 14636 12696 14648 12705
rect 14603 12668 14648 12696
rect 14636 12659 14648 12668
rect 14642 12656 14648 12659
rect 14700 12656 14706 12708
rect 16390 12696 16396 12708
rect 15764 12668 16396 12696
rect 3927 12600 8984 12628
rect 9309 12631 9367 12637
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9490 12628 9496 12640
rect 9355 12600 9496 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10183 12600 10609 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 10597 12591 10655 12597
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12628 10747 12631
rect 10778 12628 10784 12640
rect 10735 12600 10784 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 12710 12628 12716 12640
rect 11103 12600 12716 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13630 12628 13636 12640
rect 13412 12600 13636 12628
rect 13412 12588 13418 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 15764 12637 15792 12668
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 18080 12699 18138 12705
rect 18080 12665 18092 12699
rect 18126 12696 18138 12699
rect 21358 12696 21364 12708
rect 18126 12668 21364 12696
rect 18126 12665 18138 12668
rect 18080 12659 18138 12665
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 15749 12631 15807 12637
rect 15749 12597 15761 12631
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 16206 12628 16212 12640
rect 15988 12600 16212 12628
rect 15988 12588 15994 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 16356 12600 16401 12628
rect 16356 12588 16362 12600
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12393 1639 12427
rect 1581 12387 1639 12393
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12424 1915 12427
rect 1946 12424 1952 12436
rect 1903 12396 1952 12424
rect 1903 12393 1915 12396
rect 1857 12387 1915 12393
rect 1596 12356 1624 12387
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12424 2194 12436
rect 2682 12424 2688 12436
rect 2188 12396 2688 12424
rect 2188 12384 2194 12396
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5626 12424 5632 12436
rect 5583 12396 5632 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7156 12396 7205 12424
rect 7156 12384 7162 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7432 12396 7665 12424
rect 7432 12384 7438 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 8113 12427 8171 12433
rect 8113 12393 8125 12427
rect 8159 12424 8171 12427
rect 8662 12424 8668 12436
rect 8159 12396 8668 12424
rect 8159 12393 8171 12396
rect 8113 12387 8171 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 11790 12384 11796 12436
rect 11848 12384 11854 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 12216 12396 12265 12424
rect 12216 12384 12222 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12253 12387 12311 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 14642 12424 14648 12436
rect 14415 12396 14648 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 15344 12396 16313 12424
rect 15344 12384 15350 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 3970 12356 3976 12368
rect 1596 12328 3976 12356
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 4402 12359 4460 12365
rect 4402 12356 4414 12359
rect 4304 12328 4414 12356
rect 4304 12316 4310 12328
rect 4402 12325 4414 12328
rect 4448 12325 4460 12359
rect 6914 12356 6920 12368
rect 4402 12319 4460 12325
rect 5644 12328 6920 12356
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 1854 12288 1860 12300
rect 1719 12260 1860 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 1854 12248 1860 12260
rect 1912 12248 1918 12300
rect 2682 12248 2688 12300
rect 2740 12288 2746 12300
rect 5644 12297 5672 12328
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 7561 12359 7619 12365
rect 7561 12325 7573 12359
rect 7607 12356 7619 12359
rect 9122 12356 9128 12368
rect 7607 12328 9128 12356
rect 7607 12325 7619 12328
rect 7561 12319 7619 12325
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 9490 12316 9496 12368
rect 9548 12365 9554 12368
rect 9548 12359 9612 12365
rect 9548 12325 9566 12359
rect 9600 12325 9612 12359
rect 11808 12356 11836 12384
rect 9548 12319 9612 12325
rect 10796 12328 11836 12356
rect 9548 12316 9554 12319
rect 3154 12291 3212 12297
rect 3154 12288 3166 12291
rect 2740 12260 3166 12288
rect 2740 12248 2746 12260
rect 3154 12257 3166 12260
rect 3200 12257 3212 12291
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 3154 12251 3212 12257
rect 4172 12260 5641 12288
rect 3418 12220 3424 12232
rect 3331 12192 3424 12220
rect 3418 12180 3424 12192
rect 3476 12220 3482 12232
rect 4172 12229 4200 12260
rect 5629 12257 5641 12260
rect 5675 12257 5687 12291
rect 5896 12291 5954 12297
rect 5896 12288 5908 12291
rect 5629 12251 5687 12257
rect 5736 12260 5908 12288
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 3476 12192 4169 12220
rect 3476 12180 3482 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 5350 12180 5356 12232
rect 5408 12220 5414 12232
rect 5736 12220 5764 12260
rect 5896 12257 5908 12260
rect 5942 12288 5954 12291
rect 7466 12288 7472 12300
rect 5942 12260 7472 12288
rect 5942 12257 5954 12260
rect 5896 12251 5954 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 10796 12297 10824 12328
rect 13262 12316 13268 12368
rect 13320 12356 13326 12368
rect 13541 12359 13599 12365
rect 13541 12356 13553 12359
rect 13320 12328 13553 12356
rect 13320 12316 13326 12328
rect 13541 12325 13553 12328
rect 13587 12325 13599 12359
rect 16482 12356 16488 12368
rect 13541 12319 13599 12325
rect 15764 12328 16488 12356
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 8260 12260 9321 12288
rect 8260 12248 8266 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 11037 12291 11095 12297
rect 11037 12288 11049 12291
rect 10781 12251 10839 12257
rect 10888 12260 11049 12288
rect 5408 12192 5764 12220
rect 5408 12180 5414 12192
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 6880 12192 7757 12220
rect 6880 12180 6886 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 10888 12220 10916 12260
rect 11037 12257 11049 12260
rect 11083 12257 11095 12291
rect 11037 12251 11095 12257
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 11848 12260 12633 12288
rect 11848 12248 11854 12260
rect 12621 12257 12633 12260
rect 12667 12257 12679 12291
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12621 12251 12679 12257
rect 12912 12260 13461 12288
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 10744 12192 10916 12220
rect 12406 12192 12817 12220
rect 10744 12180 10750 12192
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 9306 12152 9312 12164
rect 8720 12124 9312 12152
rect 8720 12112 8726 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 12066 12112 12072 12164
rect 12124 12152 12130 12164
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 12124 12124 12173 12152
rect 12124 12112 12130 12124
rect 12161 12121 12173 12124
rect 12207 12152 12219 12155
rect 12406 12152 12434 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12207 12124 12434 12152
rect 12207 12121 12219 12124
rect 12161 12115 12219 12121
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 3108 12056 3617 12084
rect 3108 12044 3114 12056
rect 3605 12053 3617 12056
rect 3651 12084 3663 12087
rect 3878 12084 3884 12096
rect 3651 12056 3884 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 6880 12056 7021 12084
rect 6880 12044 6886 12056
rect 7009 12053 7021 12056
rect 7055 12053 7067 12087
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 7009 12047 7067 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 12912 12084 12940 12260
rect 13449 12257 13461 12260
rect 13495 12288 13507 12291
rect 13814 12288 13820 12300
rect 13495 12260 13820 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 15470 12248 15476 12300
rect 15528 12297 15534 12300
rect 15528 12288 15540 12297
rect 15654 12288 15660 12300
rect 15528 12260 15660 12288
rect 15528 12251 15540 12260
rect 15528 12248 15534 12251
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15764 12297 15792 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 16206 12288 16212 12300
rect 16167 12260 16212 12288
rect 15749 12251 15807 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 13630 12220 13636 12232
rect 13591 12192 13636 12220
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 16390 12220 16396 12232
rect 16351 12192 16396 12220
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 11112 12056 12940 12084
rect 11112 12044 11118 12056
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 15841 12087 15899 12093
rect 15841 12084 15853 12087
rect 14056 12056 15853 12084
rect 14056 12044 14062 12056
rect 15841 12053 15853 12056
rect 15887 12053 15899 12087
rect 15841 12047 15899 12053
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 2314 11880 2320 11892
rect 2275 11852 2320 11880
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 3292 11852 3617 11880
rect 3292 11840 3298 11852
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 7190 11880 7196 11892
rect 5767 11852 7196 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 11241 11883 11299 11889
rect 7432 11852 8294 11880
rect 7432 11840 7438 11852
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 7006 11812 7012 11824
rect 4028 11784 7012 11812
rect 4028 11772 4034 11784
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 8266 11812 8294 11852
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11790 11880 11796 11892
rect 11287 11852 11796 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12342 11880 12348 11892
rect 12216 11852 12348 11880
rect 12216 11840 12222 11852
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12526 11880 12532 11892
rect 12487 11852 12532 11880
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 14921 11883 14979 11889
rect 14921 11849 14933 11883
rect 14967 11880 14979 11883
rect 16206 11880 16212 11892
rect 14967 11852 16212 11880
rect 14967 11849 14979 11852
rect 14921 11843 14979 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 13170 11812 13176 11824
rect 8266 11784 13176 11812
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2130 11744 2136 11756
rect 1811 11716 2136 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2682 11704 2688 11756
rect 2740 11744 2746 11756
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2740 11716 3065 11744
rect 2740 11704 2746 11716
rect 3053 11713 3065 11716
rect 3099 11744 3111 11747
rect 4062 11744 4068 11756
rect 3099 11716 4068 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 4062 11704 4068 11716
rect 4120 11744 4126 11756
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 4120 11716 4169 11744
rect 4120 11704 4126 11716
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 6822 11744 6828 11756
rect 5215 11716 6828 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6972 11716 7205 11744
rect 6972 11704 6978 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 9122 11744 9128 11756
rect 9083 11716 9128 11744
rect 7193 11707 7251 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9272 11716 9321 11744
rect 9272 11704 9278 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 10686 11744 10692 11756
rect 10599 11716 10692 11744
rect 9309 11707 9367 11713
rect 10686 11704 10692 11716
rect 10744 11744 10750 11756
rect 10870 11744 10876 11756
rect 10744 11716 10876 11744
rect 10744 11704 10750 11716
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11790 11744 11796 11756
rect 11112 11716 11796 11744
rect 11112 11704 11118 11716
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11974 11744 11980 11756
rect 11935 11716 11980 11744
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12124 11716 13093 11744
rect 12124 11704 12130 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14642 11744 14648 11756
rect 14415 11716 14648 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 16482 11744 16488 11756
rect 16443 11716 16488 11744
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11676 2927 11679
rect 3878 11676 3884 11688
rect 2915 11648 3884 11676
rect 2915 11645 2927 11648
rect 2869 11639 2927 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 5258 11676 5264 11688
rect 3988 11648 5264 11676
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 2777 11611 2835 11617
rect 1903 11580 2452 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 1949 11543 2007 11549
rect 1949 11509 1961 11543
rect 1995 11540 2007 11543
rect 2314 11540 2320 11552
rect 1995 11512 2320 11540
rect 1995 11509 2007 11512
rect 1949 11503 2007 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2424 11549 2452 11580
rect 2777 11577 2789 11611
rect 2823 11608 2835 11611
rect 3602 11608 3608 11620
rect 2823 11580 3608 11608
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 3988 11552 4016 11648
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6270 11676 6276 11688
rect 6144 11648 6276 11676
rect 6144 11636 6150 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 8938 11676 8944 11688
rect 7392 11648 8944 11676
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 7392 11608 7420 11648
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9401 11679 9459 11685
rect 9401 11645 9413 11679
rect 9447 11676 9459 11679
rect 9582 11676 9588 11688
rect 9447 11648 9588 11676
rect 9447 11645 9459 11648
rect 9401 11639 9459 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10284 11648 10793 11676
rect 10284 11636 10290 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 14274 11676 14280 11688
rect 10781 11639 10839 11645
rect 12544 11648 14280 11676
rect 4672 11580 7420 11608
rect 7460 11611 7518 11617
rect 4672 11568 4678 11580
rect 7460 11577 7472 11611
rect 7506 11608 7518 11611
rect 7558 11608 7564 11620
rect 7506 11580 7564 11608
rect 7506 11577 7518 11580
rect 7460 11571 7518 11577
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10321 11611 10379 11617
rect 10321 11608 10333 11611
rect 9732 11580 10333 11608
rect 9732 11568 9738 11580
rect 10321 11577 10333 11580
rect 10367 11577 10379 11611
rect 10321 11571 10379 11577
rect 2409 11543 2467 11549
rect 2409 11509 2421 11543
rect 2455 11509 2467 11543
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 2409 11503 2467 11509
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 3970 11540 3976 11552
rect 3931 11512 3976 11540
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4522 11540 4528 11552
rect 4111 11512 4528 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 5258 11540 5264 11552
rect 5219 11512 5264 11540
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 5442 11540 5448 11552
rect 5399 11512 5448 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8444 11512 8585 11540
rect 8444 11500 8450 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9640 11512 9781 11540
rect 9640 11500 9646 11512
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 10336 11540 10364 11571
rect 10962 11568 10968 11620
rect 11020 11608 11026 11620
rect 12069 11611 12127 11617
rect 12069 11608 12081 11611
rect 11020 11580 12081 11608
rect 11020 11568 11026 11580
rect 12069 11577 12081 11580
rect 12115 11577 12127 11611
rect 12544 11608 12572 11648
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 16229 11679 16287 11685
rect 16229 11645 16241 11679
rect 16275 11676 16287 11679
rect 16390 11676 16396 11688
rect 16275 11648 16396 11676
rect 16275 11645 16287 11648
rect 16229 11639 16287 11645
rect 16390 11636 16396 11648
rect 16448 11636 16454 11688
rect 12069 11571 12127 11577
rect 12176 11580 12572 11608
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10336 11512 10885 11540
rect 9769 11503 9827 11509
rect 10873 11509 10885 11512
rect 10919 11540 10931 11543
rect 12176 11540 12204 11580
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 12676 11580 13001 11608
rect 12676 11568 12682 11580
rect 12989 11577 13001 11580
rect 13035 11577 13047 11611
rect 12989 11571 13047 11577
rect 10919 11512 12204 11540
rect 12437 11543 12495 11549
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12526 11540 12532 11552
rect 12483 11512 12532 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 14458 11540 14464 11552
rect 14419 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14550 11500 14556 11552
rect 14608 11540 14614 11552
rect 14608 11512 14653 11540
rect 14608 11500 14614 11512
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14792 11512 15117 11540
rect 14792 11500 14798 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1857 11339 1915 11345
rect 1857 11305 1869 11339
rect 1903 11305 1915 11339
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 1857 11299 1915 11305
rect 1872 11268 1900 11299
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 3234 11336 3240 11348
rect 2731 11308 3240 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 3375 11308 3985 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 3973 11305 3985 11308
rect 4019 11336 4031 11339
rect 4890 11336 4896 11348
rect 4019 11308 4896 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8527 11308 9137 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9582 11336 9588 11348
rect 9543 11308 9588 11336
rect 9125 11299 9183 11305
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 14090 11336 14096 11348
rect 14051 11308 14096 11336
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14461 11339 14519 11345
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 14550 11336 14556 11348
rect 14507 11308 14556 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 9953 11271 10011 11277
rect 9953 11268 9965 11271
rect 1872 11240 9965 11268
rect 9953 11237 9965 11240
rect 9999 11237 10011 11271
rect 9953 11231 10011 11237
rect 11793 11271 11851 11277
rect 11793 11237 11805 11271
rect 11839 11268 11851 11271
rect 14108 11268 14136 11296
rect 14366 11268 14372 11280
rect 11839 11240 14044 11268
rect 14108 11240 14372 11268
rect 11839 11237 11851 11240
rect 11793 11231 11851 11237
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1486 11200 1492 11212
rect 1443 11172 1492 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 4614 11200 4620 11212
rect 2240 11172 4620 11200
rect 1504 11132 1532 11160
rect 2133 11135 2191 11141
rect 2133 11132 2145 11135
rect 1504 11104 2145 11132
rect 2133 11101 2145 11104
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 2240 11064 2268 11172
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5902 11200 5908 11212
rect 5123 11172 5908 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6822 11209 6828 11212
rect 6816 11200 6828 11209
rect 6783 11172 6828 11200
rect 6816 11163 6828 11172
rect 6822 11160 6828 11163
rect 6880 11160 6886 11212
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11200 9551 11203
rect 10318 11200 10324 11212
rect 9539 11172 10324 11200
rect 9539 11169 9551 11172
rect 9493 11163 9551 11169
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11882 11200 11888 11212
rect 11296 11172 11888 11200
rect 11296 11160 11302 11172
rect 11882 11160 11888 11172
rect 11940 11200 11946 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11940 11172 12173 11200
rect 11940 11160 11946 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 12342 11200 12348 11212
rect 12299 11172 12348 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 2777 11135 2835 11141
rect 2777 11132 2789 11135
rect 1627 11036 2268 11064
rect 2608 11104 2789 11132
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 1949 10999 2007 11005
rect 1949 10996 1961 10999
rect 1544 10968 1961 10996
rect 1544 10956 1550 10968
rect 1949 10965 1961 10968
rect 1995 10965 2007 10999
rect 2608 10996 2636 11104
rect 2777 11101 2789 11104
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 2869 11095 2927 11101
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 2884 11064 2912 11095
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 3602 11132 3608 11144
rect 3563 11104 3608 11132
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 2740 11036 2912 11064
rect 3513 11067 3571 11073
rect 2740 11024 2746 11036
rect 3513 11033 3525 11067
rect 3559 11064 3571 11067
rect 3878 11064 3884 11076
rect 3559 11036 3884 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4908 11064 4936 11095
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 5040 11104 5085 11132
rect 5040 11092 5046 11104
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 5868 11104 6561 11132
rect 5868 11092 5874 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 8386 11132 8392 11144
rect 8347 11104 8392 11132
rect 6549 11095 6607 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 8496 11104 9689 11132
rect 5350 11064 5356 11076
rect 4908 11036 5356 11064
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7616 11036 7941 11064
rect 7616 11024 7622 11036
rect 7929 11033 7941 11036
rect 7975 11064 7987 11067
rect 8496 11064 8524 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9950 11092 9956 11144
rect 10008 11132 10014 11144
rect 10045 11135 10103 11141
rect 10045 11132 10057 11135
rect 10008 11104 10057 11132
rect 10008 11092 10014 11104
rect 10045 11101 10057 11104
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 10928 11104 12081 11132
rect 10928 11092 10934 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 7975 11036 8524 11064
rect 8941 11067 8999 11073
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 8941 11033 8953 11067
rect 8987 11064 8999 11067
rect 10594 11064 10600 11076
rect 8987 11036 10600 11064
rect 8987 11033 8999 11036
rect 8941 11027 8999 11033
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 12084 11064 12112 11095
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 12768 11104 13185 11132
rect 12768 11092 12774 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13280 11064 13308 11095
rect 12084 11036 13308 11064
rect 14016 11064 14044 11240
rect 14366 11228 14372 11240
rect 14424 11268 14430 11280
rect 14921 11271 14979 11277
rect 14921 11268 14933 11271
rect 14424 11240 14933 11268
rect 14424 11228 14430 11240
rect 14921 11237 14933 11240
rect 14967 11237 14979 11271
rect 14921 11231 14979 11237
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14875 11172 15301 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15470 11132 15476 11144
rect 15068 11104 15476 11132
rect 15068 11092 15074 11104
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 17126 11064 17132 11076
rect 14016 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 3326 10996 3332 11008
rect 2608 10968 3332 10996
rect 1949 10959 2007 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 9953 10999 10011 11005
rect 9953 10965 9965 10999
rect 9999 10996 10011 10999
rect 11790 10996 11796 11008
rect 9999 10968 11796 10996
rect 9999 10965 10011 10968
rect 9953 10959 10011 10965
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12342 10996 12348 11008
rect 12124 10968 12348 10996
rect 12124 10956 12130 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12618 10996 12624 11008
rect 12579 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12713 10999 12771 11005
rect 12713 10965 12725 10999
rect 12759 10996 12771 10999
rect 12894 10996 12900 11008
rect 12759 10968 12900 10996
rect 12759 10965 12771 10968
rect 12713 10959 12771 10965
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 4982 10792 4988 10804
rect 1627 10764 4988 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5258 10792 5264 10804
rect 5123 10764 5264 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 8113 10795 8171 10801
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 8570 10792 8576 10804
rect 8159 10764 8576 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10376 10764 10517 10792
rect 10376 10752 10382 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11020 10764 14412 10792
rect 11020 10752 11026 10764
rect 2958 10684 2964 10736
rect 3016 10724 3022 10736
rect 4065 10727 4123 10733
rect 4065 10724 4077 10727
rect 3016 10696 4077 10724
rect 3016 10684 3022 10696
rect 4065 10693 4077 10696
rect 4111 10724 4123 10727
rect 14384 10724 14412 10764
rect 14458 10752 14464 10804
rect 14516 10792 14522 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 14516 10764 14933 10792
rect 14516 10752 14522 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 16574 10724 16580 10736
rect 4111 10696 4752 10724
rect 14384 10696 16580 10724
rect 4111 10693 4123 10696
rect 4065 10687 4123 10693
rect 4356 10600 4384 10696
rect 4724 10665 4752 10696
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4709 10619 4767 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5408 10628 5641 10656
rect 5408 10616 5414 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5902 10656 5908 10668
rect 5863 10628 5908 10656
rect 5629 10619 5687 10625
rect 5902 10616 5908 10628
rect 5960 10616 5966 10668
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6604 10628 6745 10656
rect 6604 10616 6610 10628
rect 6733 10625 6745 10628
rect 6779 10656 6791 10659
rect 6822 10656 6828 10668
rect 6779 10628 6828 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 6822 10616 6828 10628
rect 6880 10656 6886 10668
rect 7558 10656 7564 10668
rect 6880 10628 7052 10656
rect 7519 10628 7564 10656
rect 6880 10616 6886 10628
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 3970 10588 3976 10600
rect 1811 10560 3976 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4338 10548 4344 10600
rect 4396 10548 4402 10600
rect 5442 10548 5448 10600
rect 5500 10588 5506 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5500 10560 5549 10588
rect 5500 10548 5506 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 6914 10588 6920 10600
rect 6875 10560 6920 10588
rect 5537 10551 5595 10557
rect 6914 10548 6920 10560
rect 6972 10548 6978 10600
rect 7024 10588 7052 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 11238 10656 11244 10668
rect 11195 10628 11244 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 8386 10588 8392 10600
rect 7024 10560 7880 10588
rect 8347 10560 8392 10588
rect 2032 10523 2090 10529
rect 2032 10489 2044 10523
rect 2078 10520 2090 10523
rect 2498 10520 2504 10532
rect 2078 10492 2504 10520
rect 2078 10489 2090 10492
rect 2032 10483 2090 10489
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 6825 10523 6883 10529
rect 6825 10489 6837 10523
rect 6871 10520 6883 10523
rect 7006 10520 7012 10532
rect 6871 10492 7012 10520
rect 6871 10489 6883 10492
rect 6825 10483 6883 10489
rect 7006 10480 7012 10492
rect 7064 10480 7070 10532
rect 7745 10523 7803 10529
rect 7745 10520 7757 10523
rect 7300 10492 7757 10520
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 4212 10424 4261 10452
rect 4212 10412 4218 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4614 10452 4620 10464
rect 4575 10424 4620 10452
rect 4249 10415 4307 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 7300 10461 7328 10492
rect 7745 10489 7757 10492
rect 7791 10489 7803 10523
rect 7852 10520 7880 10560
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 8645 10591 8703 10597
rect 8645 10588 8657 10591
rect 8536 10560 8657 10588
rect 8536 10548 8542 10560
rect 8645 10557 8657 10560
rect 8691 10557 8703 10591
rect 8645 10551 8703 10557
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 11164 10588 11192 10619
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 14369 10659 14427 10665
rect 12483 10628 12848 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 9180 10560 11192 10588
rect 12529 10591 12587 10597
rect 9180 10548 9186 10560
rect 12529 10557 12541 10591
rect 12575 10588 12587 10591
rect 12713 10591 12771 10597
rect 12713 10588 12725 10591
rect 12575 10560 12725 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 12713 10557 12725 10560
rect 12759 10557 12771 10591
rect 12820 10588 12848 10628
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 15010 10656 15016 10668
rect 14415 10628 15016 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 12820 10560 13124 10588
rect 12713 10551 12771 10557
rect 9140 10520 9168 10548
rect 13096 10532 13124 10560
rect 7852 10492 9168 10520
rect 10873 10523 10931 10529
rect 7745 10483 7803 10489
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 12618 10520 12624 10532
rect 10919 10492 12624 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 12618 10480 12624 10492
rect 12676 10520 12682 10532
rect 12802 10520 12808 10532
rect 12676 10492 12808 10520
rect 12676 10480 12682 10492
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 12894 10480 12900 10532
rect 12952 10529 12958 10532
rect 12952 10523 13016 10529
rect 12952 10489 12970 10523
rect 13004 10489 13016 10523
rect 12952 10483 13016 10489
rect 12952 10480 12958 10483
rect 13078 10480 13084 10532
rect 13136 10480 13142 10532
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5316 10424 5457 10452
rect 5316 10412 5322 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 5445 10415 5503 10421
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10421 7343 10455
rect 7650 10452 7656 10464
rect 7611 10424 7656 10452
rect 7285 10415 7343 10421
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 9766 10452 9772 10464
rect 9727 10424 9772 10452
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10318 10452 10324 10464
rect 10279 10424 10324 10452
rect 10318 10412 10324 10424
rect 10376 10452 10382 10464
rect 10962 10452 10968 10464
rect 10376 10424 10968 10452
rect 10376 10412 10382 10424
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 11882 10452 11888 10464
rect 11839 10424 11888 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12492 10424 12541 10452
rect 12492 10412 12498 10424
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 14090 10452 14096 10464
rect 14051 10424 14096 10452
rect 12529 10415 12587 10421
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 14734 10452 14740 10464
rect 14599 10424 14740 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10217 1639 10251
rect 1581 10211 1639 10217
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2038 10248 2044 10260
rect 1903 10220 2044 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 1596 10180 1624 10211
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2222 10248 2228 10260
rect 2179 10220 2228 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2682 10248 2688 10260
rect 2363 10220 2688 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 3881 10251 3939 10257
rect 3881 10217 3893 10251
rect 3927 10248 3939 10251
rect 4246 10248 4252 10260
rect 3927 10220 4252 10248
rect 3927 10217 3939 10220
rect 3881 10211 3939 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 4672 10220 5365 10248
rect 4672 10208 4678 10220
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5353 10211 5411 10217
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 7650 10248 7656 10260
rect 7147 10220 7656 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9447 10220 9965 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 9953 10211 10011 10217
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 10100 10220 10425 10248
rect 10100 10208 10106 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 14461 10251 14519 10257
rect 14461 10248 14473 10251
rect 11296 10220 14473 10248
rect 11296 10208 11302 10220
rect 14461 10217 14473 10220
rect 14507 10217 14519 10251
rect 14461 10211 14519 10217
rect 3694 10180 3700 10192
rect 1596 10152 3700 10180
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 4890 10140 4896 10192
rect 4948 10180 4954 10192
rect 4994 10183 5052 10189
rect 4994 10180 5006 10183
rect 4948 10152 5006 10180
rect 4948 10140 4954 10152
rect 4994 10149 5006 10152
rect 5040 10180 5052 10183
rect 6822 10180 6828 10192
rect 5040 10152 6828 10180
rect 5040 10149 5052 10152
rect 4994 10143 5052 10149
rect 6822 10140 6828 10152
rect 6880 10180 6886 10192
rect 6880 10152 7880 10180
rect 6880 10140 6886 10152
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1486 10112 1492 10124
rect 1443 10084 1492 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 3441 10115 3499 10121
rect 3441 10081 3453 10115
rect 3487 10112 3499 10115
rect 3602 10112 3608 10124
rect 3487 10084 3608 10112
rect 3487 10081 3499 10084
rect 3441 10075 3499 10081
rect 1964 9908 1992 10075
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 3988 10084 5273 10112
rect 3988 10056 4016 10084
rect 5261 10081 5273 10084
rect 5307 10112 5319 10115
rect 5810 10112 5816 10124
rect 5307 10084 5816 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6512 10084 6745 10112
rect 6512 10072 6518 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 6733 10075 6791 10081
rect 7576 10084 7665 10112
rect 3697 10047 3755 10053
rect 3697 10013 3709 10047
rect 3743 10044 3755 10047
rect 3970 10044 3976 10056
rect 3743 10016 3976 10044
rect 3743 10013 3755 10016
rect 3697 10007 3755 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 6656 9976 6684 10007
rect 6730 9976 6736 9988
rect 6656 9948 6736 9976
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 7576 9976 7604 10084
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 7852 10053 7880 10152
rect 10226 10140 10232 10192
rect 10284 10180 10290 10192
rect 10321 10183 10379 10189
rect 10321 10180 10333 10183
rect 10284 10152 10333 10180
rect 10284 10140 10290 10152
rect 10321 10149 10333 10152
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 11440 10152 11836 10180
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 11440 10121 11468 10152
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10081 11483 10115
rect 11681 10115 11739 10121
rect 11681 10112 11693 10115
rect 11425 10075 11483 10081
rect 11532 10084 11693 10112
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 9180 10016 9229 10044
rect 9180 10004 9186 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10226 10044 10232 10056
rect 9824 10016 10232 10044
rect 9824 10004 9830 10016
rect 10226 10004 10232 10016
rect 10284 10044 10290 10056
rect 10505 10047 10563 10053
rect 10505 10044 10517 10047
rect 10284 10016 10517 10044
rect 10284 10004 10290 10016
rect 10505 10013 10517 10016
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11532 10044 11560 10084
rect 11681 10081 11693 10084
rect 11727 10081 11739 10115
rect 11808 10112 11836 10152
rect 12986 10140 12992 10192
rect 13044 10180 13050 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 13044 10152 13185 10180
rect 13044 10140 13050 10152
rect 13173 10149 13185 10152
rect 13219 10180 13231 10183
rect 13219 10152 13952 10180
rect 13219 10149 13231 10152
rect 13173 10143 13231 10149
rect 12434 10112 12440 10124
rect 11808 10084 12440 10112
rect 11681 10075 11739 10081
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 13188 10084 13369 10112
rect 13188 10056 13216 10084
rect 13357 10081 13369 10084
rect 13403 10112 13415 10115
rect 13446 10112 13452 10124
rect 13403 10084 13452 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13446 10072 13452 10084
rect 13504 10112 13510 10124
rect 13924 10121 13952 10152
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 15574 10183 15632 10189
rect 15574 10180 15586 10183
rect 14148 10152 15586 10180
rect 14148 10140 14154 10152
rect 15574 10149 15586 10152
rect 15620 10149 15632 10183
rect 15574 10143 15632 10149
rect 13817 10115 13875 10121
rect 13817 10112 13829 10115
rect 13504 10084 13829 10112
rect 13504 10072 13510 10084
rect 13817 10081 13829 10084
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 16114 10112 16120 10124
rect 13955 10084 16120 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 11112 10016 11560 10044
rect 11112 10004 11118 10016
rect 13170 10004 13176 10056
rect 13228 10004 13234 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14642 10044 14648 10056
rect 14139 10016 14648 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 15838 10044 15844 10056
rect 15799 10016 15844 10044
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 9306 9976 9312 9988
rect 7576 9948 9312 9976
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 9784 9948 11192 9976
rect 4890 9908 4896 9920
rect 1964 9880 4896 9908
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 5960 9880 7297 9908
rect 5960 9868 5966 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9784 9908 9812 9948
rect 9272 9880 9812 9908
rect 9861 9911 9919 9917
rect 9272 9868 9278 9880
rect 9861 9877 9873 9911
rect 9907 9908 9919 9911
rect 11054 9908 11060 9920
rect 9907 9880 11060 9908
rect 9907 9877 9919 9880
rect 9861 9871 9919 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11164 9908 11192 9948
rect 12342 9908 12348 9920
rect 11164 9880 12348 9908
rect 12342 9868 12348 9880
rect 12400 9908 12406 9920
rect 12710 9908 12716 9920
rect 12400 9880 12716 9908
rect 12400 9868 12406 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12805 9911 12863 9917
rect 12805 9877 12817 9911
rect 12851 9908 12863 9911
rect 12894 9908 12900 9920
rect 12851 9880 12900 9908
rect 12851 9877 12863 9880
rect 12805 9871 12863 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13446 9908 13452 9920
rect 13407 9880 13452 9908
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 9214 9704 9220 9716
rect 3752 9676 9220 9704
rect 3752 9664 3758 9676
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 10318 9704 10324 9716
rect 9324 9676 10324 9704
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 1903 9608 3740 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 1412 9540 2237 9568
rect 1412 9512 1440 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2314 9528 2320 9580
rect 2372 9568 2378 9580
rect 2372 9540 2636 9568
rect 2372 9528 2378 9540
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1636 9472 1685 9500
rect 1636 9460 1642 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1673 9463 1731 9469
rect 1688 9432 1716 9463
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2056 9472 2421 9500
rect 2056 9432 2084 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 1688 9404 2084 9432
rect 2608 9432 2636 9540
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 2740 9472 2785 9500
rect 2740 9460 2746 9472
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2608 9404 2789 9432
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 3712 9432 3740 9608
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3844 9608 3985 9636
rect 3844 9596 3850 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 4890 9636 4896 9648
rect 4851 9608 4896 9636
rect 3973 9599 4031 9605
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 9324 9636 9352 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 8536 9608 9352 9636
rect 8536 9596 8542 9608
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 11517 9639 11575 9645
rect 11020 9608 11468 9636
rect 11020 9596 11026 9608
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4212 9540 4537 9568
rect 4212 9528 4218 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5258 9568 5264 9580
rect 4856 9540 5264 9568
rect 4856 9528 4862 9540
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 5718 9568 5724 9580
rect 5583 9540 5724 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 8294 9568 8300 9580
rect 8128 9540 8300 9568
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 4304 9472 4353 9500
rect 4304 9460 4310 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5902 9500 5908 9512
rect 4479 9472 5908 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6178 9500 6184 9512
rect 6139 9472 6184 9500
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 8128 9500 8156 9540
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 8404 9540 9321 9568
rect 8404 9512 8432 9540
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 10686 9528 10692 9580
rect 10744 9568 10750 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10744 9540 10885 9568
rect 10744 9528 10750 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 11054 9568 11060 9580
rect 11015 9540 11060 9568
rect 10873 9531 10931 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 11440 9568 11468 9608
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 11563 9608 12434 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11440 9540 11805 9568
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 6288 9472 8156 9500
rect 8205 9503 8263 9509
rect 6288 9432 6316 9472
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8386 9500 8392 9512
rect 8251 9472 8392 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 3712 9404 6316 9432
rect 2777 9395 2835 9401
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 7938 9435 7996 9441
rect 7938 9432 7950 9435
rect 7524 9404 7950 9432
rect 7524 9392 7530 9404
rect 7938 9401 7950 9404
rect 7984 9401 7996 9435
rect 7938 9395 7996 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2866 9364 2872 9376
rect 2179 9336 2872 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3510 9364 3516 9376
rect 3016 9336 3516 9364
rect 3016 9324 3022 9336
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5534 9364 5540 9376
rect 5399 9336 5540 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5868 9336 6009 9364
rect 5868 9324 5874 9336
rect 5997 9333 6009 9336
rect 6043 9364 6055 9367
rect 8220 9364 8248 9463
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9225 9503 9283 9509
rect 9225 9469 9237 9503
rect 9271 9500 9283 9503
rect 9950 9500 9956 9512
rect 9271 9472 9956 9500
rect 9271 9469 9283 9472
rect 9225 9463 9283 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 12406 9500 12434 9608
rect 12526 9596 12532 9648
rect 12584 9636 12590 9648
rect 12584 9608 13308 9636
rect 12584 9596 12590 9608
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13280 9577 13308 9608
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 13964 9608 14565 9636
rect 13964 9596 13970 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12952 9540 13093 9568
rect 12952 9528 12958 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14090 9568 14096 9580
rect 14047 9540 14096 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 13357 9503 13415 9509
rect 12406 9472 12664 9500
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 9554 9435 9612 9441
rect 9554 9432 9566 9435
rect 9180 9404 9566 9432
rect 9180 9392 9186 9404
rect 9554 9401 9566 9404
rect 9600 9401 9612 9435
rect 9554 9395 9612 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11790 9432 11796 9444
rect 11112 9404 11796 9432
rect 11112 9392 11118 9404
rect 11790 9392 11796 9404
rect 11848 9432 11854 9444
rect 11977 9435 12035 9441
rect 11977 9432 11989 9435
rect 11848 9404 11989 9432
rect 11848 9392 11854 9404
rect 11977 9401 11989 9404
rect 12023 9401 12035 9435
rect 11977 9395 12035 9401
rect 12069 9435 12127 9441
rect 12069 9401 12081 9435
rect 12115 9432 12127 9435
rect 12529 9435 12587 9441
rect 12529 9432 12541 9435
rect 12115 9404 12541 9432
rect 12115 9401 12127 9404
rect 12069 9395 12127 9401
rect 12529 9401 12541 9404
rect 12575 9401 12587 9435
rect 12636 9432 12664 9472
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13446 9500 13452 9512
rect 13403 9472 13452 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 13596 9472 14197 9500
rect 13596 9460 13602 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 18690 9432 18696 9444
rect 12636 9404 18696 9432
rect 12529 9395 12587 9401
rect 18690 9392 18696 9404
rect 18748 9392 18754 9444
rect 9030 9364 9036 9376
rect 6043 9336 8248 9364
rect 8991 9336 9036 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 12437 9367 12495 9373
rect 12437 9364 12449 9367
rect 12216 9336 12449 9364
rect 12216 9324 12222 9336
rect 12437 9333 12449 9336
rect 12483 9333 12495 9367
rect 12437 9327 12495 9333
rect 13725 9367 13783 9373
rect 13725 9333 13737 9367
rect 13771 9364 13783 9367
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 13771 9336 14105 9364
rect 13771 9333 13783 9336
rect 13725 9327 13783 9333
rect 14093 9333 14105 9336
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1728 9132 1869 9160
rect 1728 9120 1734 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 1857 9123 1915 9129
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2363 9132 2789 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 2777 9123 2835 9129
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 3936 9132 4261 9160
rect 3936 9120 3942 9132
rect 4249 9129 4261 9132
rect 4295 9160 4307 9163
rect 5074 9160 5080 9172
rect 4295 9132 5080 9160
rect 4295 9129 4307 9132
rect 4249 9123 4307 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5718 9160 5724 9172
rect 5679 9132 5724 9160
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7742 9160 7748 9172
rect 7699 9132 7748 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8159 9132 8248 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 5736 9092 5764 9120
rect 6058 9095 6116 9101
rect 6058 9092 6070 9095
rect 1636 9064 5672 9092
rect 5736 9064 6070 9092
rect 1636 9052 1642 9064
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 9024 1458 9036
rect 1673 9027 1731 9033
rect 1673 9024 1685 9027
rect 1452 8996 1685 9024
rect 1452 8984 1458 8996
rect 1673 8993 1685 8996
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 2096 8996 2237 9024
rect 2096 8984 2102 8996
rect 2225 8993 2237 8996
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3510 9024 3516 9036
rect 3191 8996 3516 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4608 9027 4666 9033
rect 4608 8993 4620 9027
rect 4654 9024 4666 9027
rect 4890 9024 4896 9036
rect 4654 8996 4896 9024
rect 4654 8993 4666 8996
rect 4608 8987 4666 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5644 9024 5672 9064
rect 6058 9061 6070 9064
rect 6104 9061 6116 9095
rect 8220 9092 8248 9132
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8352 9132 10456 9160
rect 8352 9120 8358 9132
rect 8754 9092 8760 9104
rect 6058 9055 6116 9061
rect 6196 9064 8156 9092
rect 8220 9064 8760 9092
rect 6196 9024 6224 9064
rect 5644 8996 6224 9024
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 8128 9024 8156 9064
rect 8754 9052 8760 9064
rect 8812 9092 8818 9104
rect 10134 9092 10140 9104
rect 8812 9064 10140 9092
rect 8812 9052 8818 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10226 9052 10232 9104
rect 10284 9101 10290 9104
rect 10284 9092 10296 9101
rect 10428 9092 10456 9132
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 10560 9132 11253 9160
rect 10560 9120 10566 9132
rect 11241 9129 11253 9132
rect 11287 9129 11299 9163
rect 11241 9123 11299 9129
rect 11701 9163 11759 9169
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11747 9132 12081 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 12529 9163 12587 9169
rect 12216 9132 12261 9160
rect 12216 9120 12222 9132
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 13538 9160 13544 9172
rect 12575 9132 13544 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 14608 9132 14657 9160
rect 14608 9120 14614 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 13262 9092 13268 9104
rect 10284 9064 10329 9092
rect 10428 9064 13268 9092
rect 10284 9055 10296 9064
rect 10284 9052 10290 9055
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 17126 9092 17132 9104
rect 13464 9064 17132 9092
rect 8128 8996 10640 9024
rect 8021 8987 8079 8993
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2409 8959 2467 8965
rect 2409 8956 2421 8959
rect 2188 8928 2421 8956
rect 2188 8916 2194 8928
rect 2409 8925 2421 8928
rect 2455 8925 2467 8959
rect 2409 8919 2467 8925
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3234 8956 3240 8968
rect 2648 8928 3096 8956
rect 3195 8928 3240 8956
rect 2648 8916 2654 8928
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 3068 8888 3096 8928
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3344 8888 3372 8919
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 4028 8928 4353 8956
rect 4028 8916 4034 8928
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 4341 8919 4399 8925
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 8036 8956 8064 8987
rect 8110 8956 8116 8968
rect 8036 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 7193 8891 7251 8897
rect 1627 8860 2774 8888
rect 3068 8860 3372 8888
rect 3528 8860 4384 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 2746 8820 2774 8860
rect 3528 8820 3556 8860
rect 3694 8820 3700 8832
rect 2746 8792 3556 8820
rect 3655 8792 3700 8820
rect 3694 8780 3700 8792
rect 3752 8820 3758 8832
rect 4246 8820 4252 8832
rect 3752 8792 4252 8820
rect 3752 8780 3758 8792
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4356 8820 4384 8860
rect 7193 8857 7205 8891
rect 7239 8888 7251 8891
rect 7466 8888 7472 8900
rect 7239 8860 7472 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7466 8848 7472 8860
rect 7524 8888 7530 8900
rect 8220 8888 8248 8919
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8444 8928 8493 8956
rect 8444 8916 8450 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9398 8956 9404 8968
rect 8720 8928 9404 8956
rect 8720 8916 8726 8928
rect 9398 8916 9404 8928
rect 9456 8916 9462 8968
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 7524 8860 8248 8888
rect 8404 8860 9628 8888
rect 7524 8848 7530 8860
rect 8404 8820 8432 8860
rect 9122 8820 9128 8832
rect 4356 8792 8432 8820
rect 9083 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9600 8820 9628 8860
rect 10318 8820 10324 8832
rect 9600 8792 10324 8820
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 10520 8820 10548 8919
rect 10612 8888 10640 8996
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11020 8996 11345 9024
rect 11020 8984 11026 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 12894 9024 12900 9036
rect 11333 8987 11391 8993
rect 11992 8996 12900 9024
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11992 8965 12020 8996
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 8993 13047 9027
rect 13464 9024 13492 9064
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 13630 9024 13636 9036
rect 12989 8987 13047 8993
rect 13280 8996 13492 9024
rect 13591 8996 13636 9024
rect 11057 8959 11115 8965
rect 11057 8956 11069 8959
rect 10928 8928 11069 8956
rect 10928 8916 10934 8928
rect 11057 8925 11069 8928
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8925 12035 8959
rect 11977 8919 12035 8925
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 13004 8956 13032 8987
rect 12216 8928 13032 8956
rect 12216 8916 12222 8928
rect 12250 8888 12256 8900
rect 10612 8860 12256 8888
rect 12250 8848 12256 8860
rect 12308 8848 12314 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 13280 8888 13308 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8925 13415 8959
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13357 8919 13415 8925
rect 12768 8860 13308 8888
rect 13372 8888 13400 8919
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 14056 8928 14381 8956
rect 14056 8916 14062 8928
rect 14369 8925 14381 8928
rect 14415 8925 14427 8959
rect 14369 8919 14427 8925
rect 13906 8888 13912 8900
rect 13372 8860 13912 8888
rect 12768 8848 12774 8860
rect 13906 8848 13912 8860
rect 13964 8848 13970 8900
rect 15286 8888 15292 8900
rect 14016 8860 15292 8888
rect 12434 8820 12440 8832
rect 10520 8792 12440 8820
rect 12434 8780 12440 8792
rect 12492 8820 12498 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 12492 8792 13185 8820
rect 12492 8780 12498 8792
rect 13173 8789 13185 8792
rect 13219 8820 13231 8823
rect 13722 8820 13728 8832
rect 13219 8792 13728 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14016 8829 14044 8860
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 14001 8823 14059 8829
rect 14001 8789 14013 8823
rect 14047 8789 14059 8823
rect 14001 8783 14059 8789
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15194 8820 15200 8832
rect 14967 8792 15200 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15194 8780 15200 8792
rect 15252 8780 15258 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 3510 8616 3516 8628
rect 1627 8588 3372 8616
rect 3471 8588 3516 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 3344 8548 3372 8588
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5534 8616 5540 8628
rect 4948 8588 5304 8616
rect 5495 8588 5540 8616
rect 4948 8576 4954 8588
rect 3344 8520 5212 8548
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3160 8452 4077 8480
rect 3160 8424 3188 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4890 8480 4896 8492
rect 4488 8452 4896 8480
rect 4488 8440 4494 8452
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5074 8480 5080 8492
rect 5031 8452 5080 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 1394 8412 1400 8424
rect 1307 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8412 1458 8424
rect 2682 8412 2688 8424
rect 1452 8384 2688 8412
rect 1452 8372 1458 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 2981 8415 3039 8421
rect 2981 8381 2993 8415
rect 3027 8412 3039 8415
rect 3142 8412 3148 8424
rect 3027 8384 3148 8412
rect 3027 8381 3039 8384
rect 2981 8375 3039 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3970 8412 3976 8424
rect 3283 8384 3976 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 1673 8347 1731 8353
rect 1673 8344 1685 8347
rect 1544 8316 1685 8344
rect 1544 8304 1550 8316
rect 1673 8313 1685 8316
rect 1719 8313 1731 8347
rect 1673 8307 1731 8313
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3252 8344 3280 8375
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 2924 8316 3280 8344
rect 2924 8304 2930 8316
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 3752 8316 3893 8344
rect 3752 8304 3758 8316
rect 3881 8313 3893 8316
rect 3927 8344 3939 8347
rect 4617 8347 4675 8353
rect 3927 8316 4476 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 2590 8276 2596 8288
rect 1903 8248 2596 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 3326 8276 3332 8288
rect 3287 8248 3332 8276
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3973 8279 4031 8285
rect 3973 8245 3985 8279
rect 4019 8276 4031 8279
rect 4246 8276 4252 8288
rect 4019 8248 4252 8276
rect 4019 8245 4031 8248
rect 3973 8239 4031 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4448 8276 4476 8316
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 5077 8347 5135 8353
rect 5077 8344 5089 8347
rect 4663 8316 5089 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 5077 8313 5089 8316
rect 5123 8313 5135 8347
rect 5184 8344 5212 8520
rect 5276 8412 5304 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6730 8616 6736 8628
rect 6236 8588 6736 8616
rect 6236 8576 6242 8588
rect 6730 8576 6736 8588
rect 6788 8616 6794 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 6788 8588 7849 8616
rect 6788 8576 6794 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 7837 8579 7895 8585
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8662 8616 8668 8628
rect 8343 8588 8668 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9490 8616 9496 8628
rect 9263 8588 9496 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6012 8520 6469 8548
rect 6012 8489 6040 8520
rect 6457 8517 6469 8520
rect 6503 8517 6515 8551
rect 6457 8511 6515 8517
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 8846 8548 8852 8560
rect 7708 8520 8852 8548
rect 7708 8508 7714 8520
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 9140 8548 9168 8579
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 11146 8616 11152 8628
rect 10152 8588 11152 8616
rect 10152 8548 10180 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 9140 8520 10180 8548
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10689 8551 10747 8557
rect 10689 8548 10701 8551
rect 10652 8520 10701 8548
rect 10652 8508 10658 8520
rect 10689 8517 10701 8520
rect 10735 8517 10747 8551
rect 10689 8511 10747 8517
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 11885 8551 11943 8557
rect 10836 8520 11284 8548
rect 10836 8508 10842 8520
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 6104 8412 6132 8443
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6236 8452 7021 8480
rect 6236 8440 6242 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 9122 8480 9128 8492
rect 8619 8452 9128 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9456 8452 9689 8480
rect 9456 8440 9462 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 9858 8480 9864 8492
rect 9771 8452 9864 8480
rect 9677 8443 9735 8449
rect 9858 8440 9864 8452
rect 9916 8480 9922 8492
rect 10226 8480 10232 8492
rect 9916 8452 10232 8480
rect 9916 8440 9922 8452
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 10962 8480 10968 8492
rect 10376 8452 10968 8480
rect 10376 8440 10382 8452
rect 10962 8440 10968 8452
rect 11020 8480 11026 8492
rect 11256 8489 11284 8520
rect 11885 8517 11897 8551
rect 11931 8548 11943 8551
rect 12158 8548 12164 8560
rect 11931 8520 12164 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 14734 8548 14740 8560
rect 12308 8520 14740 8548
rect 12308 8508 12314 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 11020 8452 11161 8480
rect 11020 8440 11026 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 12710 8480 12716 8492
rect 11241 8443 11299 8449
rect 12406 8452 12716 8480
rect 7650 8412 7656 8424
rect 5276 8384 6132 8412
rect 6748 8384 7656 8412
rect 6748 8344 6776 8384
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 9030 8412 9036 8424
rect 8067 8384 9036 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 9030 8372 9036 8384
rect 9088 8412 9094 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 9088 8384 11713 8412
rect 9088 8372 9094 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 12406 8412 12434 8452
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12860 8452 12909 8480
rect 12860 8440 12866 8452
rect 12897 8449 12909 8452
rect 12943 8480 12955 8483
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 12943 8452 14197 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 14185 8449 14197 8452
rect 14231 8480 14243 8483
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14231 8452 15117 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 12986 8412 12992 8424
rect 11701 8375 11759 8381
rect 11808 8384 12434 8412
rect 12544 8384 12992 8412
rect 5184 8316 6776 8344
rect 6825 8347 6883 8353
rect 5077 8307 5135 8313
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 7006 8344 7012 8356
rect 6871 8316 7012 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 7282 8344 7288 8356
rect 7116 8316 7288 8344
rect 4890 8276 4896 8288
rect 4448 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 5316 8248 5457 8276
rect 5316 8236 5322 8248
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5445 8239 5503 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7116 8276 7144 8316
rect 7282 8304 7288 8316
rect 7340 8344 7346 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 7340 8316 7389 8344
rect 7340 8304 7346 8316
rect 7377 8313 7389 8316
rect 7423 8344 7435 8347
rect 8202 8344 8208 8356
rect 7423 8316 8208 8344
rect 7423 8313 7435 8316
rect 7377 8307 7435 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 8803 8316 10057 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 10045 8313 10057 8316
rect 10091 8313 10103 8347
rect 10045 8307 10103 8313
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 11808 8344 11836 8384
rect 12544 8344 12572 8384
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 13262 8412 13268 8424
rect 13219 8384 13268 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13998 8412 14004 8424
rect 13959 8384 14004 8412
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14608 8384 14933 8412
rect 14608 8372 14614 8384
rect 14921 8381 14933 8384
rect 14967 8412 14979 8415
rect 15654 8412 15660 8424
rect 14967 8384 15660 8412
rect 14967 8381 14979 8384
rect 14921 8375 14979 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 12710 8344 12716 8356
rect 10192 8316 11836 8344
rect 11900 8316 12572 8344
rect 12623 8316 12716 8344
rect 10192 8304 10198 8316
rect 8662 8276 8668 8288
rect 6963 8248 7144 8276
rect 8623 8248 8668 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 9582 8276 9588 8288
rect 9543 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 11054 8276 11060 8288
rect 11015 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11900 8276 11928 8316
rect 12710 8304 12716 8316
rect 12768 8344 12774 8356
rect 13081 8347 13139 8353
rect 13081 8344 13093 8347
rect 12768 8316 13093 8344
rect 12768 8304 12774 8316
rect 13081 8313 13093 8316
rect 13127 8344 13139 8347
rect 13354 8344 13360 8356
rect 13127 8316 13360 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 13872 8316 14105 8344
rect 13872 8304 13878 8316
rect 14093 8313 14105 8316
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14240 8316 15025 8344
rect 14240 8304 14246 8316
rect 15013 8313 15025 8316
rect 15059 8344 15071 8347
rect 15194 8344 15200 8356
rect 15059 8316 15200 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 15194 8304 15200 8316
rect 15252 8344 15258 8356
rect 16390 8344 16396 8356
rect 15252 8316 16396 8344
rect 15252 8304 15258 8316
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 13538 8276 13544 8288
rect 11204 8248 11928 8276
rect 13499 8248 13544 8276
rect 11204 8236 11210 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 14550 8276 14556 8288
rect 14511 8248 14556 8276
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8041 1455 8075
rect 1397 8035 1455 8041
rect 1412 8004 1440 8035
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 12710 8072 12716 8084
rect 1636 8044 12716 8072
rect 1636 8032 1642 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 13906 8072 13912 8084
rect 13867 8044 13912 8072
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 2130 8004 2136 8016
rect 1412 7976 2136 8004
rect 2130 7964 2136 7976
rect 2188 7964 2194 8016
rect 2590 8013 2596 8016
rect 2532 8007 2596 8013
rect 2532 7973 2544 8007
rect 2578 7973 2596 8007
rect 2532 7967 2596 7973
rect 2590 7964 2596 7967
rect 2648 7964 2654 8016
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 5258 8004 5264 8016
rect 4120 7976 5264 8004
rect 4120 7964 4126 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5568 8007 5626 8013
rect 5568 7973 5580 8007
rect 5614 8004 5626 8007
rect 6178 8004 6184 8016
rect 5614 7976 6184 8004
rect 5614 7973 5626 7976
rect 5568 7967 5626 7973
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 7009 8007 7067 8013
rect 7009 7973 7021 8007
rect 7055 8004 7067 8007
rect 7098 8004 7104 8016
rect 7055 7976 7104 8004
rect 7055 7973 7067 7976
rect 7009 7967 7067 7973
rect 7098 7964 7104 7976
rect 7156 7964 7162 8016
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 9677 8007 9735 8013
rect 9677 8004 9689 8007
rect 7708 7976 9689 8004
rect 7708 7964 7714 7976
rect 9677 7973 9689 7976
rect 9723 8004 9735 8007
rect 9766 8004 9772 8016
rect 9723 7976 9772 8004
rect 9723 7973 9735 7976
rect 9677 7967 9735 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10686 8013 10692 8016
rect 10680 7967 10692 8013
rect 10744 8004 10750 8016
rect 10744 7976 10780 8004
rect 10686 7964 10692 7967
rect 10744 7964 10750 7976
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11790 8004 11796 8016
rect 11112 7976 11796 8004
rect 11112 7964 11118 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 13924 8004 13952 8032
rect 14614 8007 14672 8013
rect 14614 8004 14626 8007
rect 12544 7976 13768 8004
rect 13924 7976 14626 8004
rect 12544 7948 12572 7976
rect 13740 7948 13768 7976
rect 14614 7973 14626 7976
rect 14660 7973 14672 8007
rect 15838 8004 15844 8016
rect 14614 7967 14672 7973
rect 14752 7976 15844 8004
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 2866 7936 2872 7948
rect 2823 7908 2872 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 3016 7908 3249 7936
rect 3016 7896 3022 7908
rect 3237 7905 3249 7908
rect 3283 7905 3295 7939
rect 3237 7899 3295 7905
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 5810 7936 5816 7948
rect 3375 7908 4200 7936
rect 5771 7908 5816 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 4172 7877 4200 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7282 7936 7288 7948
rect 6963 7908 7288 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7432 7908 7757 7936
rect 7432 7896 7438 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9490 7936 9496 7948
rect 8996 7908 9496 7936
rect 8996 7896 9002 7908
rect 9490 7896 9496 7908
rect 9548 7936 9554 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9548 7908 9597 7936
rect 9548 7896 9554 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 12526 7936 12532 7948
rect 12439 7908 12532 7936
rect 9585 7899 9643 7905
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12802 7945 12808 7948
rect 12796 7936 12808 7945
rect 12763 7908 12808 7936
rect 12796 7899 12808 7908
rect 12802 7896 12808 7899
rect 12860 7896 12866 7948
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 13780 7908 14381 7936
rect 13780 7896 13786 7908
rect 14369 7905 14381 7908
rect 14415 7936 14427 7939
rect 14752 7936 14780 7976
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 16097 7939 16155 7945
rect 16097 7936 16109 7939
rect 14415 7908 14780 7936
rect 15764 7908 16109 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3200 7840 3433 7868
rect 3200 7828 3206 7840
rect 3421 7837 3433 7840
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 6270 7868 6276 7880
rect 4203 7840 4844 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4430 7800 4436 7812
rect 4391 7772 4436 7800
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 2866 7732 2872 7744
rect 2827 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3476 7704 3893 7732
rect 3476 7692 3482 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 3881 7695 3939 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4816 7732 4844 7840
rect 5828 7840 6276 7868
rect 5828 7812 5856 7840
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 7190 7868 7196 7880
rect 7151 7840 7196 7868
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7760 7840 7849 7868
rect 7760 7812 7788 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8294 7868 8300 7880
rect 8067 7840 8300 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 5810 7760 5816 7812
rect 5868 7760 5874 7812
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6457 7803 6515 7809
rect 6457 7800 6469 7803
rect 5960 7772 6469 7800
rect 5960 7760 5966 7772
rect 6457 7769 6469 7772
rect 6503 7800 6515 7803
rect 6503 7772 7696 7800
rect 6503 7769 6515 7772
rect 6457 7763 6515 7769
rect 7668 7744 7696 7772
rect 7742 7760 7748 7812
rect 7800 7760 7806 7812
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 9217 7803 9275 7809
rect 9217 7800 9229 7803
rect 8720 7772 9229 7800
rect 8720 7760 8726 7772
rect 9217 7769 9229 7772
rect 9263 7769 9275 7803
rect 9217 7763 9275 7769
rect 15764 7744 15792 7908
rect 16097 7905 16109 7908
rect 16143 7905 16155 7939
rect 16097 7899 16155 7905
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 15896 7840 15941 7868
rect 15896 7828 15902 7840
rect 6086 7732 6092 7744
rect 4816 7704 6092 7732
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7377 7735 7435 7741
rect 7377 7732 7389 7735
rect 7156 7704 7389 7732
rect 7156 7692 7162 7704
rect 7377 7701 7389 7704
rect 7423 7701 7435 7735
rect 7650 7732 7656 7744
rect 7563 7704 7656 7732
rect 7377 7695 7435 7701
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 11146 7732 11152 7744
rect 7708 7704 11152 7732
rect 7708 7692 7714 7704
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 15746 7732 15752 7744
rect 15707 7704 15752 7732
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 17218 7732 17224 7744
rect 17179 7704 17224 7732
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 3292 7500 3525 7528
rect 3292 7488 3298 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 3936 7500 4353 7528
rect 3936 7488 3942 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 5810 7528 5816 7540
rect 4663 7500 5816 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 3160 7432 4108 7460
rect 3160 7404 3188 7432
rect 2774 7392 2780 7404
rect 2735 7364 2780 7392
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3142 7392 3148 7404
rect 3007 7364 3148 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 4080 7401 4108 7432
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7324 2010 7336
rect 3326 7324 3332 7336
rect 2004 7296 3332 7324
rect 2004 7284 2010 7296
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4632 7324 4660 7491
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 7374 7528 7380 7540
rect 6319 7500 7380 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8536 7500 8953 7528
rect 8536 7488 8542 7500
rect 8941 7497 8953 7500
rect 8987 7528 8999 7531
rect 10778 7528 10784 7540
rect 8987 7500 10784 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 4706 7420 4712 7472
rect 4764 7460 4770 7472
rect 5074 7460 5080 7472
rect 4764 7432 5080 7460
rect 4764 7420 4770 7432
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 7190 7460 7196 7472
rect 7116 7432 7196 7460
rect 5718 7392 5724 7404
rect 5679 7364 5724 7392
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 7116 7401 7144 7432
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 7101 7395 7159 7401
rect 6512 7364 6868 7392
rect 6512 7352 6518 7364
rect 4019 7296 4660 7324
rect 5905 7327 5963 7333
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6546 7324 6552 7336
rect 5951 7296 6552 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 6840 7333 6868 7364
rect 7101 7361 7113 7395
rect 7147 7361 7159 7395
rect 7282 7392 7288 7404
rect 7243 7364 7288 7392
rect 7101 7355 7159 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 9674 7392 9680 7404
rect 9635 7364 9680 7392
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12342 7392 12348 7404
rect 12207 7364 12348 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 13964 7364 14197 7392
rect 13964 7352 13970 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7392 14427 7395
rect 14550 7392 14556 7404
rect 14415 7364 14556 7392
rect 14415 7361 14427 7364
rect 14369 7355 14427 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15746 7392 15752 7404
rect 15151 7364 15752 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7561 7327 7619 7333
rect 7561 7324 7573 7327
rect 6972 7296 7573 7324
rect 6972 7284 6978 7296
rect 7561 7293 7573 7296
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9548 7296 9781 7324
rect 9548 7284 9554 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 15286 7324 15292 7336
rect 12308 7296 12388 7324
rect 15247 7296 15292 7324
rect 12308 7284 12314 7296
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7256 2743 7259
rect 3145 7259 3203 7265
rect 3145 7256 3157 7259
rect 2731 7228 3157 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3145 7225 3157 7228
rect 3191 7225 3203 7259
rect 3145 7219 3203 7225
rect 3510 7216 3516 7268
rect 3568 7256 3574 7268
rect 4709 7259 4767 7265
rect 4709 7256 4721 7259
rect 3568 7228 4721 7256
rect 3568 7216 3574 7228
rect 4709 7225 4721 7228
rect 4755 7225 4767 7259
rect 4709 7219 4767 7225
rect 5813 7259 5871 7265
rect 5813 7225 5825 7259
rect 5859 7256 5871 7259
rect 7828 7259 7886 7265
rect 5859 7228 6316 7256
rect 5859 7225 5871 7228
rect 5813 7219 5871 7225
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2222 7188 2228 7200
rect 2179 7160 2228 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2406 7188 2412 7200
rect 2363 7160 2412 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 4338 7188 4344 7200
rect 3292 7160 4344 7188
rect 3292 7148 3298 7160
rect 4338 7148 4344 7160
rect 4396 7188 4402 7200
rect 4893 7191 4951 7197
rect 4893 7188 4905 7191
rect 4396 7160 4905 7188
rect 4396 7148 4402 7160
rect 4893 7157 4905 7160
rect 4939 7157 4951 7191
rect 4893 7151 4951 7157
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 5215 7160 5457 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 5445 7157 5457 7160
rect 5491 7188 5503 7191
rect 5534 7188 5540 7200
rect 5491 7160 5540 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 6288 7188 6316 7228
rect 7828 7225 7840 7259
rect 7874 7256 7886 7259
rect 8294 7256 8300 7268
rect 7874 7228 8300 7256
rect 7874 7225 7886 7228
rect 7828 7219 7886 7225
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 8662 7216 8668 7268
rect 8720 7256 8726 7268
rect 11054 7256 11060 7268
rect 8720 7228 11060 7256
rect 8720 7216 8726 7228
rect 11054 7216 11060 7228
rect 11112 7256 11118 7268
rect 12360 7265 12388 7296
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 12345 7259 12403 7265
rect 11112 7228 12296 7256
rect 11112 7216 11118 7228
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 6288 7160 6469 7188
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 6917 7191 6975 7197
rect 6917 7188 6929 7191
rect 6880 7160 6929 7188
rect 6880 7148 6886 7160
rect 6917 7157 6929 7160
rect 6963 7157 6975 7191
rect 6917 7151 6975 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10229 7191 10287 7197
rect 9916 7160 9961 7188
rect 9916 7148 9922 7160
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10870 7188 10876 7200
rect 10275 7160 10876 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 12268 7197 12296 7228
rect 12345 7225 12357 7259
rect 12391 7225 12403 7259
rect 12345 7219 12403 7225
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 14461 7259 14519 7265
rect 14461 7256 14473 7259
rect 12952 7228 14473 7256
rect 12952 7216 12958 7228
rect 14461 7225 14473 7228
rect 14507 7225 14519 7259
rect 14461 7219 14519 7225
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7157 12311 7191
rect 12253 7151 12311 7157
rect 12713 7191 12771 7197
rect 12713 7157 12725 7191
rect 12759 7188 12771 7191
rect 14274 7188 14280 7200
rect 12759 7160 14280 7188
rect 12759 7157 12771 7160
rect 12713 7151 12771 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7188 14887 7191
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 14875 7160 15209 7188
rect 14875 7157 14887 7160
rect 14829 7151 14887 7157
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15436 7160 15669 7188
rect 15436 7148 15442 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 1670 6944 1676 6996
rect 1728 6944 1734 6996
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 5074 6984 5080 6996
rect 3375 6956 5080 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 5258 6984 5264 6996
rect 5219 6956 5264 6984
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7190 6944 7196 6996
rect 7248 6944 7254 6996
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 9674 6944 9680 6996
rect 9732 6944 9738 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10137 6987 10195 6993
rect 10137 6984 10149 6987
rect 9916 6956 10149 6984
rect 9916 6944 9922 6956
rect 10137 6953 10149 6956
rect 10183 6953 10195 6987
rect 10137 6947 10195 6953
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10686 6984 10692 6996
rect 10376 6956 10692 6984
rect 10376 6944 10382 6956
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 1688 6916 1716 6944
rect 3418 6916 3424 6928
rect 1688 6888 3424 6916
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 4249 6919 4307 6925
rect 4249 6885 4261 6919
rect 4295 6916 4307 6919
rect 4982 6916 4988 6928
rect 4295 6888 4988 6916
rect 4295 6885 4307 6888
rect 4249 6879 4307 6885
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 5626 6916 5632 6928
rect 5368 6888 5632 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1486 6848 1492 6860
rect 1443 6820 1492 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 2501 6851 2559 6857
rect 1719 6820 2452 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1688 6780 1716 6811
rect 1360 6752 1716 6780
rect 1360 6740 1366 6752
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 2424 6712 2452 6820
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2866 6848 2872 6860
rect 2547 6820 2872 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4341 6851 4399 6857
rect 3384 6820 4292 6848
rect 3384 6808 3390 6820
rect 2590 6780 2596 6792
rect 2551 6752 2596 6780
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3283 6752 3924 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3896 6721 3924 6752
rect 3881 6715 3939 6721
rect 1903 6684 2360 6712
rect 2424 6684 3832 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2332 6644 2360 6684
rect 3326 6644 3332 6656
rect 2332 6616 3332 6644
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3694 6644 3700 6656
rect 3655 6616 3700 6644
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3804 6644 3832 6684
rect 3881 6681 3893 6715
rect 3927 6681 3939 6715
rect 4264 6712 4292 6820
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4798 6848 4804 6860
rect 4387 6820 4804 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4893 6851 4951 6857
rect 4893 6817 4905 6851
rect 4939 6848 4951 6851
rect 5368 6848 5396 6888
rect 5626 6876 5632 6888
rect 5684 6916 5690 6928
rect 6362 6916 6368 6928
rect 5684 6888 6368 6916
rect 5684 6876 5690 6888
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 6580 6919 6638 6925
rect 6580 6885 6592 6919
rect 6626 6916 6638 6919
rect 7208 6916 7236 6944
rect 9692 6916 9720 6944
rect 10888 6916 10916 6947
rect 10962 6944 10968 6996
rect 11020 6984 11026 6996
rect 14734 6984 14740 6996
rect 11020 6956 14504 6984
rect 14695 6956 14740 6984
rect 11020 6944 11026 6956
rect 11054 6916 11060 6928
rect 6626 6888 7236 6916
rect 9508 6888 11060 6916
rect 6626 6885 6638 6888
rect 6580 6879 6638 6885
rect 5718 6848 5724 6860
rect 4939 6820 5396 6848
rect 5460 6820 5724 6848
rect 4939 6817 4951 6820
rect 4893 6811 4951 6817
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4982 6780 4988 6792
rect 4571 6752 4988 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5460 6721 5488 6820
rect 5718 6808 5724 6820
rect 5776 6848 5782 6860
rect 7184 6851 7242 6857
rect 7184 6848 7196 6851
rect 5776 6820 7196 6848
rect 5776 6808 5782 6820
rect 7184 6817 7196 6820
rect 7230 6848 7242 6851
rect 7466 6848 7472 6860
rect 7230 6820 7472 6848
rect 7230 6817 7242 6820
rect 7184 6811 7242 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 9508 6848 9536 6888
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 11790 6876 11796 6928
rect 11848 6916 11854 6928
rect 11986 6919 12044 6925
rect 11986 6916 11998 6919
rect 11848 6888 11998 6916
rect 11848 6876 11854 6888
rect 11986 6885 11998 6888
rect 12032 6885 12044 6919
rect 14476 6916 14504 6956
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 11986 6879 12044 6885
rect 12084 6888 14320 6916
rect 14476 6888 14780 6916
rect 9416 6820 9536 6848
rect 9677 6851 9735 6857
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 6914 6780 6920 6792
rect 6871 6752 6920 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 9416 6789 9444 6820
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9766 6848 9772 6860
rect 9723 6820 9772 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 12084 6848 12112 6888
rect 9876 6820 12112 6848
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6749 9459 6783
rect 9582 6780 9588 6792
rect 9543 6752 9588 6780
rect 9401 6743 9459 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 5445 6715 5503 6721
rect 4264 6684 5396 6712
rect 3881 6675 3939 6681
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 3804 6616 4721 6644
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4856 6616 5089 6644
rect 4856 6604 4862 6616
rect 5077 6613 5089 6616
rect 5123 6613 5135 6647
rect 5368 6644 5396 6684
rect 5445 6681 5457 6715
rect 5491 6681 5503 6715
rect 5445 6675 5503 6681
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8662 6712 8668 6724
rect 7984 6684 8668 6712
rect 7984 6672 7990 6684
rect 8662 6672 8668 6684
rect 8720 6712 8726 6724
rect 9766 6712 9772 6724
rect 8720 6684 9772 6712
rect 8720 6672 8726 6684
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 9876 6644 9904 6820
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 12216 6820 12357 6848
rect 12216 6808 12222 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 14292 6848 14320 6888
rect 14458 6848 14464 6860
rect 14292 6820 14464 6848
rect 12345 6811 12403 6817
rect 14458 6808 14464 6820
rect 14516 6848 14522 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14516 6820 14657 6848
rect 14516 6808 14522 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14752 6848 14780 6888
rect 19058 6848 19064 6860
rect 14752 6820 19064 6848
rect 14645 6811 14703 6817
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10962 6780 10968 6792
rect 10008 6752 10968 6780
rect 10008 6740 10014 6752
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6780 12311 6783
rect 12526 6780 12532 6792
rect 12299 6752 12532 6780
rect 12299 6749 12311 6752
rect 12253 6743 12311 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 14550 6780 14556 6792
rect 14511 6752 14556 6780
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 10744 6684 11376 6712
rect 10744 6672 10750 6684
rect 5368 6616 9904 6644
rect 10045 6647 10103 6653
rect 5077 6607 5135 6613
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10778 6644 10784 6656
rect 10091 6616 10784 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11348 6644 11376 6684
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 16298 6712 16304 6724
rect 12492 6684 16304 6712
rect 12492 6672 12498 6684
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 12526 6644 12532 6656
rect 11348 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 15105 6647 15163 6653
rect 15105 6613 15117 6647
rect 15151 6644 15163 6647
rect 15470 6644 15476 6656
rect 15151 6616 15476 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 3237 6443 3295 6449
rect 1627 6412 3188 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 3160 6372 3188 6412
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 3326 6440 3332 6452
rect 3283 6412 3332 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 3326 6400 3332 6412
rect 3384 6440 3390 6452
rect 3602 6440 3608 6452
rect 3384 6412 3608 6440
rect 3384 6400 3390 6412
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 6822 6440 6828 6452
rect 4080 6412 6828 6440
rect 4080 6372 4108 6412
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7800 6412 7849 6440
rect 7800 6400 7806 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 7837 6403 7895 6409
rect 7944 6412 12480 6440
rect 3160 6344 4108 6372
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 5445 6375 5503 6381
rect 5445 6372 5457 6375
rect 4212 6344 5457 6372
rect 4212 6332 4218 6344
rect 5445 6341 5457 6344
rect 5491 6341 5503 6375
rect 7944 6372 7972 6412
rect 5445 6335 5503 6341
rect 5552 6344 7972 6372
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 1670 6236 1676 6248
rect 1443 6208 1676 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 1670 6196 1676 6208
rect 1728 6196 1734 6248
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 2102 6171 2160 6177
rect 2102 6168 2114 6171
rect 1820 6140 2114 6168
rect 1820 6128 1826 6140
rect 2102 6137 2114 6140
rect 2148 6168 2160 6171
rect 3142 6168 3148 6180
rect 2148 6140 3148 6168
rect 2148 6137 2160 6140
rect 2102 6131 2160 6137
rect 3142 6128 3148 6140
rect 3200 6168 3206 6180
rect 3988 6168 4016 6267
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4764 6276 4813 6304
rect 4764 6264 4770 6276
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 4982 6304 4988 6316
rect 4895 6276 4988 6304
rect 4801 6267 4859 6273
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 5132 6276 5181 6304
rect 5132 6264 5138 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 5000 6236 5028 6264
rect 5552 6236 5580 6344
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 12250 6372 12256 6384
rect 10560 6344 10605 6372
rect 10704 6344 12256 6372
rect 10560 6332 10566 6344
rect 6086 6304 6092 6316
rect 6047 6276 6092 6304
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 7190 6304 7196 6316
rect 6595 6276 7052 6304
rect 7151 6276 7196 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 5718 6236 5724 6248
rect 4580 6208 5580 6236
rect 5679 6208 5724 6236
rect 4580 6196 4586 6208
rect 5718 6196 5724 6208
rect 5776 6236 5782 6248
rect 5994 6236 6000 6248
rect 5776 6208 6000 6236
rect 5776 6196 5782 6208
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6730 6236 6736 6248
rect 6691 6208 6736 6236
rect 6730 6196 6736 6208
rect 6788 6196 6794 6248
rect 7024 6236 7052 6276
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 7524 6276 8401 6304
rect 7524 6264 7530 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 10704 6304 10732 6344
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 8389 6267 8447 6273
rect 10336 6276 10732 6304
rect 7742 6236 7748 6248
rect 7024 6208 7748 6236
rect 7742 6196 7748 6208
rect 7800 6236 7806 6248
rect 10336 6236 10364 6276
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 10836 6276 10977 6304
rect 10836 6264 10842 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 12452 6304 12480 6412
rect 14016 6412 18337 6440
rect 12529 6375 12587 6381
rect 12529 6341 12541 6375
rect 12575 6372 12587 6375
rect 12894 6372 12900 6384
rect 12575 6344 12900 6372
rect 12575 6341 12587 6344
rect 12529 6335 12587 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 14016 6304 14044 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 12452 6276 14044 6304
rect 11977 6267 12035 6273
rect 7800 6208 10364 6236
rect 10413 6239 10471 6245
rect 7800 6196 7806 6208
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10686 6236 10692 6248
rect 10459 6208 10692 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10870 6236 10876 6248
rect 10831 6208 10876 6236
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11072 6236 11100 6267
rect 10980 6208 11100 6236
rect 11992 6236 12020 6267
rect 11992 6208 12434 6236
rect 3200 6140 4016 6168
rect 4709 6171 4767 6177
rect 3200 6128 3206 6140
rect 4709 6137 4721 6171
rect 4755 6168 4767 6171
rect 5258 6168 5264 6180
rect 4755 6140 5264 6168
rect 4755 6137 4767 6140
rect 4709 6131 4767 6137
rect 5258 6128 5264 6140
rect 5316 6168 5322 6180
rect 6822 6168 6828 6180
rect 5316 6140 6828 6168
rect 5316 6128 5322 6140
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 7282 6168 7288 6180
rect 7243 6140 7288 6168
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 10226 6177 10232 6180
rect 8297 6171 8355 6177
rect 8297 6168 8309 6171
rect 7760 6140 8309 6168
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1673 6103 1731 6109
rect 1673 6100 1685 6103
rect 1452 6072 1685 6100
rect 1452 6060 1458 6072
rect 1673 6069 1685 6072
rect 1719 6069 1731 6103
rect 1673 6063 1731 6069
rect 3421 6103 3479 6109
rect 3421 6069 3433 6103
rect 3467 6100 3479 6103
rect 3602 6100 3608 6112
rect 3467 6072 3608 6100
rect 3467 6069 3479 6072
rect 3421 6063 3479 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 3927 6072 4353 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 4341 6069 4353 6072
rect 4387 6069 4399 6103
rect 4341 6063 4399 6069
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5813 6103 5871 6109
rect 5813 6100 5825 6103
rect 4948 6072 5825 6100
rect 4948 6060 4954 6072
rect 5813 6069 5825 6072
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6178 6100 6184 6112
rect 6052 6072 6184 6100
rect 6052 6060 6058 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6914 6100 6920 6112
rect 6788 6072 6920 6100
rect 6788 6060 6794 6072
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7374 6100 7380 6112
rect 7335 6072 7380 6100
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7760 6109 7788 6140
rect 8297 6137 8309 6140
rect 8343 6137 8355 6171
rect 10168 6171 10232 6177
rect 10168 6168 10180 6171
rect 10139 6140 10180 6168
rect 8297 6131 8355 6137
rect 10168 6137 10180 6140
rect 10214 6137 10232 6171
rect 10168 6131 10232 6137
rect 10226 6128 10232 6131
rect 10284 6168 10290 6180
rect 10980 6168 11008 6208
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 10284 6140 11008 6168
rect 11072 6140 12173 6168
rect 10284 6128 10290 6140
rect 7745 6103 7803 6109
rect 7745 6069 7757 6103
rect 7791 6069 7803 6103
rect 8202 6100 8208 6112
rect 8163 6072 8208 6100
rect 7745 6063 7803 6069
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8812 6072 9045 6100
rect 8812 6060 8818 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 11072 6100 11100 6140
rect 12161 6137 12173 6140
rect 12207 6137 12219 6171
rect 12161 6131 12219 6137
rect 9272 6072 11100 6100
rect 12069 6103 12127 6109
rect 9272 6060 9278 6072
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12250 6100 12256 6112
rect 12115 6072 12256 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12406 6100 12434 6208
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 15252 6208 16957 6236
rect 15252 6196 15258 6208
rect 16945 6205 16957 6208
rect 16991 6205 17003 6239
rect 16945 6199 17003 6205
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 14930 6171 14988 6177
rect 14930 6168 14942 6171
rect 14516 6140 14942 6168
rect 14516 6128 14522 6140
rect 14930 6137 14942 6140
rect 14976 6137 14988 6171
rect 14930 6131 14988 6137
rect 17212 6171 17270 6177
rect 17212 6137 17224 6171
rect 17258 6168 17270 6171
rect 17402 6168 17408 6180
rect 17258 6140 17408 6168
rect 17258 6137 17270 6140
rect 17212 6131 17270 6137
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 12802 6100 12808 6112
rect 12406 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6100 12866 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 12860 6072 13829 6100
rect 12860 6060 12866 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14642 6100 14648 6112
rect 14332 6072 14648 6100
rect 14332 6060 14338 6072
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15286 6100 15292 6112
rect 15247 6072 15292 6100
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 16761 6103 16819 6109
rect 16761 6069 16773 6103
rect 16807 6100 16819 6103
rect 17862 6100 17868 6112
rect 16807 6072 17868 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1762 5896 1768 5908
rect 1723 5868 1768 5896
rect 1762 5856 1768 5868
rect 1820 5856 1826 5908
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3200 5868 3740 5896
rect 3200 5856 3206 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 2464 5800 3617 5828
rect 2464 5788 2470 5800
rect 3605 5797 3617 5800
rect 3651 5797 3663 5831
rect 3605 5791 3663 5797
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 2889 5763 2947 5769
rect 2889 5729 2901 5763
rect 2935 5760 2947 5763
rect 2935 5732 3372 5760
rect 2935 5729 2947 5732
rect 2889 5723 2947 5729
rect 3142 5692 3148 5704
rect 3103 5664 3148 5692
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3344 5692 3372 5732
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 3712 5760 3740 5868
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3844 5868 3893 5896
rect 3844 5856 3850 5868
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 4246 5896 4252 5908
rect 4159 5868 4252 5896
rect 3881 5859 3939 5865
rect 4246 5856 4252 5868
rect 4304 5896 4310 5908
rect 5442 5896 5448 5908
rect 4304 5868 5448 5896
rect 4304 5856 4310 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 6052 5868 6101 5896
rect 6052 5856 6058 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 7190 5896 7196 5908
rect 6503 5868 7196 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7340 5868 7941 5896
rect 7340 5856 7346 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 7929 5859 7987 5865
rect 8128 5868 8401 5896
rect 8128 5840 8156 5868
rect 8389 5865 8401 5868
rect 8435 5896 8447 5899
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8435 5868 8953 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 8941 5865 8953 5868
rect 8987 5896 8999 5899
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8987 5868 9137 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9309 5899 9367 5905
rect 9309 5865 9321 5899
rect 9355 5896 9367 5899
rect 10226 5896 10232 5908
rect 9355 5868 10232 5896
rect 9355 5865 9367 5868
rect 9309 5859 9367 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 10781 5899 10839 5905
rect 10781 5865 10793 5899
rect 10827 5896 10839 5899
rect 10870 5896 10876 5908
rect 10827 5868 10876 5896
rect 10827 5865 10839 5868
rect 10781 5859 10839 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11149 5899 11207 5905
rect 11149 5896 11161 5899
rect 11020 5868 11161 5896
rect 11020 5856 11026 5868
rect 11149 5865 11161 5868
rect 11195 5865 11207 5899
rect 11149 5859 11207 5865
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11885 5899 11943 5905
rect 11287 5868 11652 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 4338 5828 4344 5840
rect 4299 5800 4344 5828
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 6273 5831 6331 5837
rect 6273 5828 6285 5831
rect 5592 5800 6285 5828
rect 5592 5788 5598 5800
rect 6273 5797 6285 5800
rect 6319 5828 6331 5831
rect 6638 5828 6644 5840
rect 6319 5800 6644 5828
rect 6319 5797 6331 5800
rect 6273 5791 6331 5797
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 7592 5831 7650 5837
rect 7592 5828 7604 5831
rect 7524 5800 7604 5828
rect 7524 5788 7530 5800
rect 7592 5797 7604 5800
rect 7638 5828 7650 5831
rect 7638 5800 8064 5828
rect 7638 5797 7650 5800
rect 7592 5791 7650 5797
rect 4982 5769 4988 5772
rect 4976 5760 4988 5769
rect 3476 5732 3521 5760
rect 3712 5732 4752 5760
rect 4943 5732 4988 5760
rect 3476 5720 3482 5732
rect 4522 5692 4528 5704
rect 3344 5664 4528 5692
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4724 5701 4752 5732
rect 4976 5723 4988 5732
rect 4982 5720 4988 5723
rect 5040 5720 5046 5772
rect 5718 5720 5724 5772
rect 5776 5760 5782 5772
rect 7926 5760 7932 5772
rect 5776 5732 7932 5760
rect 5776 5720 5782 5732
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8036 5760 8064 5800
rect 8110 5788 8116 5840
rect 8168 5788 8174 5840
rect 8297 5831 8355 5837
rect 8297 5797 8309 5831
rect 8343 5828 8355 5831
rect 8849 5831 8907 5837
rect 8849 5828 8861 5831
rect 8343 5800 8861 5828
rect 8343 5797 8355 5800
rect 8297 5791 8355 5797
rect 8849 5797 8861 5800
rect 8895 5828 8907 5831
rect 9950 5828 9956 5840
rect 8895 5800 9956 5828
rect 8895 5797 8907 5800
rect 8849 5791 8907 5797
rect 9950 5788 9956 5800
rect 10008 5788 10014 5840
rect 10444 5831 10502 5837
rect 10444 5797 10456 5831
rect 10490 5828 10502 5831
rect 11054 5828 11060 5840
rect 10490 5800 11060 5828
rect 10490 5797 10502 5800
rect 10444 5791 10502 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 8941 5763 8999 5769
rect 8036 5732 8340 5760
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 7834 5692 7840 5704
rect 7795 5664 7840 5692
rect 4709 5655 4767 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 4246 5624 4252 5636
rect 1627 5596 2176 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 2148 5556 2176 5596
rect 3160 5596 4252 5624
rect 3160 5556 3188 5596
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 2148 5528 3188 5556
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3786 5556 3792 5568
rect 3375 5528 3792 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4724 5556 4752 5655
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8312 5692 8340 5732
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 11624 5760 11652 5868
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 12066 5896 12072 5908
rect 11931 5868 12072 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14366 5896 14372 5908
rect 14231 5868 14372 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14366 5856 14372 5868
rect 14424 5896 14430 5908
rect 15105 5899 15163 5905
rect 14424 5868 14679 5896
rect 14424 5856 14430 5868
rect 11701 5831 11759 5837
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 11974 5828 11980 5840
rect 11747 5800 11980 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 13078 5828 13084 5840
rect 12636 5800 13084 5828
rect 12066 5760 12072 5772
rect 8987 5732 11560 5760
rect 11624 5732 12072 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8312 5664 8493 5692
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 10686 5692 10692 5704
rect 10647 5664 10692 5692
rect 8481 5655 8539 5661
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 11112 5664 11345 5692
rect 11112 5652 11118 5664
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 5902 5584 5908 5636
rect 5960 5624 5966 5636
rect 5960 5596 6776 5624
rect 5960 5584 5966 5596
rect 5920 5556 5948 5584
rect 6748 5568 6776 5596
rect 4724 5528 5948 5556
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 6638 5556 6644 5568
rect 6144 5528 6644 5556
rect 6144 5516 6150 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 7834 5556 7840 5568
rect 6788 5528 7840 5556
rect 6788 5516 6794 5528
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 10778 5556 10784 5568
rect 7984 5528 10784 5556
rect 7984 5516 7990 5528
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 11532 5556 11560 5732
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 12636 5769 12664 5800
rect 13078 5788 13084 5800
rect 13136 5788 13142 5840
rect 14651 5769 14679 5868
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15565 5899 15623 5905
rect 15565 5896 15577 5899
rect 15151 5868 15577 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15565 5865 15577 5868
rect 15611 5865 15623 5899
rect 17862 5896 17868 5908
rect 17823 5868 17868 5896
rect 15565 5859 15623 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 21358 5896 21364 5908
rect 21319 5868 21364 5896
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 14737 5831 14795 5837
rect 14737 5797 14749 5831
rect 14783 5828 14795 5831
rect 15286 5828 15292 5840
rect 14783 5800 15292 5828
rect 14783 5797 14795 5800
rect 14737 5791 14795 5797
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 17957 5831 18015 5837
rect 17957 5828 17969 5831
rect 15580 5800 17969 5828
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12584 5732 12633 5760
rect 12584 5720 12590 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12888 5763 12946 5769
rect 12888 5729 12900 5763
rect 12934 5760 12946 5763
rect 14645 5763 14703 5769
rect 12934 5732 14596 5760
rect 12934 5729 12946 5732
rect 12888 5723 12946 5729
rect 14568 5704 14596 5732
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 14826 5720 14832 5772
rect 14884 5760 14890 5772
rect 15580 5760 15608 5800
rect 17957 5797 17969 5800
rect 18003 5797 18015 5831
rect 17957 5791 18015 5797
rect 14884 5732 15608 5760
rect 16292 5763 16350 5769
rect 14884 5720 14890 5732
rect 16292 5729 16304 5763
rect 16338 5760 16350 5763
rect 21269 5763 21327 5769
rect 16338 5732 17632 5760
rect 16338 5729 16350 5732
rect 16292 5723 16350 5729
rect 14550 5692 14556 5704
rect 14511 5664 14556 5692
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14792 5664 15301 5692
rect 14792 5652 14798 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 14001 5627 14059 5633
rect 14001 5593 14013 5627
rect 14047 5624 14059 5627
rect 14752 5624 14780 5652
rect 14047 5596 14780 5624
rect 14047 5593 14059 5596
rect 14001 5587 14059 5593
rect 15194 5584 15200 5636
rect 15252 5624 15258 5636
rect 16040 5624 16068 5655
rect 17604 5636 17632 5732
rect 21269 5729 21281 5763
rect 21315 5760 21327 5763
rect 21542 5760 21548 5772
rect 21315 5732 21548 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 17402 5624 17408 5636
rect 15252 5596 16068 5624
rect 17363 5596 17408 5624
rect 15252 5584 15258 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 18064 5624 18092 5655
rect 17644 5596 18092 5624
rect 17644 5584 17650 5596
rect 14366 5556 14372 5568
rect 11532 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15933 5559 15991 5565
rect 15933 5556 15945 5559
rect 15620 5528 15945 5556
rect 15620 5516 15626 5528
rect 15933 5525 15945 5528
rect 15979 5525 15991 5559
rect 17494 5556 17500 5568
rect 17455 5528 17500 5556
rect 15933 5519 15991 5525
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 4154 5352 4160 5364
rect 1596 5324 4160 5352
rect 1486 5148 1492 5160
rect 1399 5120 1492 5148
rect 1486 5108 1492 5120
rect 1544 5148 1550 5160
rect 1596 5148 1624 5324
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 5350 5352 5356 5364
rect 4663 5324 5356 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5500 5324 6469 5352
rect 5500 5312 5506 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7377 5355 7435 5361
rect 7377 5321 7389 5355
rect 7423 5352 7435 5355
rect 8202 5352 8208 5364
rect 7423 5324 8208 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 9907 5324 19196 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 1854 5284 1860 5296
rect 1719 5256 1860 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 1854 5244 1860 5256
rect 1912 5244 1918 5296
rect 4065 5287 4123 5293
rect 4065 5253 4077 5287
rect 4111 5284 4123 5287
rect 7466 5284 7472 5296
rect 4111 5256 7328 5284
rect 7427 5256 7472 5284
rect 4111 5253 4123 5256
rect 4065 5247 4123 5253
rect 3142 5176 3148 5228
rect 3200 5176 3206 5228
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3384 5188 3433 5216
rect 3384 5176 3390 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3421 5179 3479 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4522 5176 4528 5228
rect 4580 5216 4586 5228
rect 4982 5216 4988 5228
rect 4580 5188 4988 5216
rect 4580 5176 4586 5188
rect 4982 5176 4988 5188
rect 5040 5216 5046 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 5040 5188 5181 5216
rect 5040 5176 5046 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 6178 5216 6184 5228
rect 5583 5188 6184 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7190 5216 7196 5228
rect 6871 5188 7196 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 1544 5120 1624 5148
rect 1544 5108 1550 5120
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2130 5157 2136 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1820 5120 1869 5148
rect 1820 5108 1826 5120
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 2124 5111 2136 5157
rect 2188 5148 2194 5160
rect 2188 5120 2224 5148
rect 1872 5080 1900 5111
rect 2130 5108 2136 5111
rect 2188 5108 2194 5120
rect 3160 5080 3188 5176
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 5994 5148 6000 5160
rect 5000 5120 6000 5148
rect 1872 5052 3188 5080
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 5000 5089 5028 5120
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6638 5148 6644 5160
rect 6135 5120 6644 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 4341 5083 4399 5089
rect 4341 5080 4353 5083
rect 4028 5052 4353 5080
rect 4028 5040 4034 5052
rect 4341 5049 4353 5052
rect 4387 5049 4399 5083
rect 4341 5043 4399 5049
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5049 5043 5083
rect 4985 5043 5043 5049
rect 5077 5083 5135 5089
rect 5077 5049 5089 5083
rect 5123 5080 5135 5083
rect 5810 5080 5816 5092
rect 5123 5052 5816 5080
rect 5123 5049 5135 5052
rect 5077 5043 5135 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6362 5080 6368 5092
rect 5951 5052 6368 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 6917 5083 6975 5089
rect 6917 5049 6929 5083
rect 6963 5080 6975 5083
rect 7190 5080 7196 5092
rect 6963 5052 7196 5080
rect 6963 5049 6975 5052
rect 6917 5043 6975 5049
rect 7190 5040 7196 5052
rect 7248 5040 7254 5092
rect 7300 5080 7328 5256
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 12526 5284 12532 5296
rect 9456 5256 12532 5284
rect 9456 5244 9462 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16761 5287 16819 5293
rect 16761 5284 16773 5287
rect 16540 5256 16773 5284
rect 16540 5244 16546 5256
rect 16761 5253 16773 5256
rect 16807 5284 16819 5287
rect 17586 5284 17592 5296
rect 16807 5256 17592 5284
rect 16807 5253 16819 5256
rect 16761 5247 16819 5253
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10284 5188 10517 5216
rect 10284 5176 10290 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11112 5188 11345 5216
rect 11112 5176 11118 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 11333 5179 11391 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 11848 5188 12265 5216
rect 11848 5176 11854 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 12710 5216 12716 5228
rect 12299 5188 12716 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14734 5216 14740 5228
rect 14695 5188 14740 5216
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 15252 5188 15393 5216
rect 15252 5176 15258 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 17218 5216 17224 5228
rect 15381 5179 15439 5185
rect 16408 5188 17224 5216
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8846 5148 8852 5160
rect 7892 5120 8852 5148
rect 7892 5108 7898 5120
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 10870 5148 10876 5160
rect 10367 5120 10876 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 12158 5148 12164 5160
rect 12119 5120 12164 5148
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 13348 5151 13406 5157
rect 13348 5117 13360 5151
rect 13394 5148 13406 5151
rect 14752 5148 14780 5176
rect 13394 5120 14780 5148
rect 13394 5117 13406 5120
rect 13348 5111 13406 5117
rect 8604 5083 8662 5089
rect 7300 5052 8248 5080
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3326 5012 3332 5024
rect 3283 4984 3332 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4120 4984 4169 5012
rect 4120 4972 4126 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 5718 5012 5724 5024
rect 5679 4984 5724 5012
rect 4157 4975 4215 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 6181 5015 6239 5021
rect 6181 5012 6193 5015
rect 6144 4984 6193 5012
rect 6144 4972 6150 4984
rect 6181 4981 6193 4984
rect 6227 4981 6239 5015
rect 6181 4975 6239 4981
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 5012 7067 5015
rect 7282 5012 7288 5024
rect 7055 4984 7288 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 8220 5012 8248 5052
rect 8604 5049 8616 5083
rect 8650 5080 8662 5083
rect 8754 5080 8760 5092
rect 8650 5052 8760 5080
rect 8650 5049 8662 5052
rect 8604 5043 8662 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 9030 5080 9036 5092
rect 8991 5052 9036 5080
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 9646 5052 9873 5080
rect 9646 5012 9674 5052
rect 9861 5049 9873 5052
rect 9907 5049 9919 5083
rect 9861 5043 9919 5049
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 12069 5083 12127 5089
rect 12069 5080 12081 5083
rect 12032 5052 12081 5080
rect 12032 5040 12038 5052
rect 12069 5049 12081 5052
rect 12115 5049 12127 5083
rect 12069 5043 12127 5049
rect 9950 5012 9956 5024
rect 8220 4984 9674 5012
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10781 5015 10839 5021
rect 10781 5012 10793 5015
rect 10459 4984 10793 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10781 4981 10793 4984
rect 10827 4981 10839 5015
rect 11146 5012 11152 5024
rect 11107 4984 11152 5012
rect 10781 4975 10839 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11241 5015 11299 5021
rect 11241 4981 11253 5015
rect 11287 5012 11299 5015
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11287 4984 11713 5012
rect 11287 4981 11299 4984
rect 11241 4975 11299 4981
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 12176 5012 12204 5108
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14921 5083 14979 5089
rect 14921 5080 14933 5083
rect 13688 5052 14933 5080
rect 13688 5040 13694 5052
rect 14921 5049 14933 5052
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 15470 5040 15476 5092
rect 15528 5080 15534 5092
rect 15626 5083 15684 5089
rect 15626 5080 15638 5083
rect 15528 5052 15638 5080
rect 15528 5040 15534 5052
rect 15626 5049 15638 5052
rect 15672 5080 15684 5083
rect 16408 5080 16436 5188
rect 17218 5176 17224 5188
rect 17276 5216 17282 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17276 5188 17509 5216
rect 17276 5176 17282 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 17310 5148 17316 5160
rect 17271 5120 17316 5148
rect 17310 5108 17316 5120
rect 17368 5148 17374 5160
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 17368 5120 17785 5148
rect 17368 5108 17374 5120
rect 17773 5117 17785 5120
rect 17819 5148 17831 5151
rect 18138 5148 18144 5160
rect 17819 5120 18144 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 19168 5157 19196 5324
rect 19153 5151 19211 5157
rect 19153 5117 19165 5151
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 15672 5052 16436 5080
rect 15672 5049 15684 5052
rect 15626 5043 15684 5049
rect 14274 5012 14280 5024
rect 12176 4984 14280 5012
rect 11701 4975 11759 4981
rect 14274 4972 14280 4984
rect 14332 4972 14338 5024
rect 14458 5012 14464 5024
rect 14419 4984 14464 5012
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14734 4972 14740 5024
rect 14792 5012 14798 5024
rect 14829 5015 14887 5021
rect 14829 5012 14841 5015
rect 14792 4984 14841 5012
rect 14792 4972 14798 4984
rect 14829 4981 14841 4984
rect 14875 4981 14887 5015
rect 15286 5012 15292 5024
rect 15247 4984 15292 5012
rect 14829 4975 14887 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17184 4984 17417 5012
rect 17184 4972 17190 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 17957 5015 18015 5021
rect 17957 5012 17969 5015
rect 17451 4984 17969 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 17957 4981 17969 4984
rect 18003 4981 18015 5015
rect 17957 4975 18015 4981
rect 19337 5015 19395 5021
rect 19337 4981 19349 5015
rect 19383 5012 19395 5015
rect 19978 5012 19984 5024
rect 19383 4984 19984 5012
rect 19383 4981 19395 4984
rect 19337 4975 19395 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4777 2099 4811
rect 2041 4771 2099 4777
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3142 4808 3148 4820
rect 3099 4780 3148 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 1026 4700 1032 4752
rect 1084 4740 1090 4752
rect 1489 4743 1547 4749
rect 1489 4740 1501 4743
rect 1084 4712 1501 4740
rect 1084 4700 1090 4712
rect 1489 4709 1501 4712
rect 1535 4740 1547 4743
rect 1670 4740 1676 4752
rect 1535 4712 1676 4740
rect 1535 4709 1547 4712
rect 1489 4703 1547 4709
rect 1670 4700 1676 4712
rect 1728 4700 1734 4752
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 2056 4672 2084 4771
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 3418 4808 3424 4820
rect 3375 4780 3424 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 4341 4743 4399 4749
rect 4341 4740 4353 4743
rect 3804 4712 4353 4740
rect 1811 4644 2084 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 2188 4644 2421 4672
rect 2188 4632 2194 4644
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 2861 4675 2919 4681
rect 2861 4641 2873 4675
rect 2907 4641 2919 4675
rect 2861 4635 2919 4641
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 1854 4604 1860 4616
rect 1719 4576 1860 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2498 4604 2504 4616
rect 2459 4576 2504 4604
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 2884 4604 2912 4635
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 3108 4644 3157 4672
rect 3108 4632 3114 4644
rect 3145 4641 3157 4644
rect 3191 4672 3203 4675
rect 3694 4672 3700 4684
rect 3191 4644 3700 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 3804 4616 3832 4712
rect 4341 4709 4353 4712
rect 4387 4709 4399 4743
rect 4341 4703 4399 4709
rect 4540 4684 4568 4771
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5408 4780 6285 4808
rect 5408 4768 5414 4780
rect 3878 4632 3884 4684
rect 3936 4632 3942 4684
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 4028 4644 4077 4672
rect 4028 4632 4034 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4522 4632 4528 4684
rect 4580 4632 4586 4684
rect 5626 4672 5632 4684
rect 5684 4681 5690 4684
rect 6196 4681 6224 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 7006 4808 7012 4820
rect 6967 4780 7012 4808
rect 6273 4771 6331 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 7374 4808 7380 4820
rect 7331 4780 7380 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7708 4780 8217 4808
rect 7708 4768 7714 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 8386 4768 8392 4820
rect 8444 4808 8450 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8444 4780 8585 4808
rect 8444 4768 8450 4780
rect 8573 4777 8585 4780
rect 8619 4777 8631 4811
rect 8573 4771 8631 4777
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9766 4808 9772 4820
rect 9088 4780 9772 4808
rect 9088 4768 9094 4780
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 9950 4808 9956 4820
rect 9911 4780 9956 4808
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10502 4808 10508 4820
rect 10091 4780 10508 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 11241 4811 11299 4817
rect 11241 4808 11253 4811
rect 11204 4780 11253 4808
rect 11204 4768 11210 4780
rect 11241 4777 11253 4780
rect 11287 4777 11299 4811
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 11241 4771 11299 4777
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12308 4780 13277 4808
rect 12308 4768 12314 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13265 4771 13323 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14792 4780 15117 4808
rect 14792 4768 14798 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 16807 4780 17141 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 17129 4777 17141 4780
rect 17175 4777 17187 4811
rect 17129 4771 17187 4777
rect 17221 4811 17279 4817
rect 17221 4777 17233 4811
rect 17267 4808 17279 4811
rect 17494 4808 17500 4820
rect 17267 4780 17500 4808
rect 17267 4777 17279 4780
rect 17221 4771 17279 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 7392 4712 7757 4740
rect 7392 4684 7420 4712
rect 7745 4709 7757 4712
rect 7791 4709 7803 4743
rect 9125 4743 9183 4749
rect 9125 4740 9137 4743
rect 7745 4703 7803 4709
rect 8312 4712 9137 4740
rect 8312 4684 8340 4712
rect 9125 4709 9137 4712
rect 9171 4709 9183 4743
rect 9125 4703 9183 4709
rect 9214 4700 9220 4752
rect 9272 4740 9278 4752
rect 9490 4740 9496 4752
rect 9272 4712 9496 4740
rect 9272 4700 9278 4712
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 12526 4700 12532 4752
rect 12584 4740 12590 4752
rect 12584 4712 12629 4740
rect 12584 4700 12590 4712
rect 14458 4700 14464 4752
rect 14516 4740 14522 4752
rect 15562 4740 15568 4752
rect 14516 4712 14872 4740
rect 15523 4712 15568 4740
rect 14516 4700 14522 4712
rect 5684 4675 5707 4681
rect 5559 4644 5632 4672
rect 5626 4632 5632 4644
rect 5695 4672 5707 4675
rect 6181 4675 6239 4681
rect 5695 4644 6040 4672
rect 5695 4641 5707 4644
rect 5684 4635 5707 4641
rect 5684 4632 5690 4635
rect 3605 4607 3663 4613
rect 3605 4604 3617 4607
rect 2648 4576 2693 4604
rect 2884 4576 3617 4604
rect 2648 4564 2654 4576
rect 3160 4548 3188 4576
rect 3605 4573 3617 4576
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 2314 4536 2320 4548
rect 1995 4508 2320 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 2314 4496 2320 4508
rect 2372 4496 2378 4548
rect 3142 4496 3148 4548
rect 3200 4496 3206 4548
rect 3896 4545 3924 4632
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 6012 4604 6040 4644
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7190 4672 7196 4684
rect 6963 4644 7196 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 7653 4635 7711 4641
rect 6822 4604 6828 4616
rect 6012 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7558 4604 7564 4616
rect 7064 4576 7564 4604
rect 7064 4564 7070 4576
rect 7558 4564 7564 4576
rect 7616 4604 7622 4616
rect 7668 4604 7696 4635
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 8444 4644 8677 4672
rect 8444 4632 8450 4644
rect 8665 4641 8677 4644
rect 8711 4672 8723 4675
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8711 4644 9321 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 10502 4632 10508 4684
rect 10560 4672 10566 4684
rect 10597 4675 10655 4681
rect 10597 4672 10609 4675
rect 10560 4644 10609 4672
rect 10560 4632 10566 4644
rect 10597 4641 10609 4644
rect 10643 4672 10655 4675
rect 10870 4672 10876 4684
rect 10643 4644 10876 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4672 11667 4675
rect 11974 4672 11980 4684
rect 11655 4644 11980 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4641 12495 4675
rect 12544 4672 12572 4700
rect 13173 4675 13231 4681
rect 13173 4672 13185 4675
rect 12544 4644 13185 4672
rect 12437 4635 12495 4641
rect 13173 4641 13185 4644
rect 13219 4641 13231 4675
rect 14550 4672 14556 4684
rect 13173 4635 13231 4641
rect 14476 4644 14556 4672
rect 7616 4576 7696 4604
rect 7837 4607 7895 4613
rect 7616 4564 7622 4576
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 3881 4539 3939 4545
rect 3881 4505 3893 4539
rect 3927 4505 3939 4539
rect 7282 4536 7288 4548
rect 3881 4499 3939 4505
rect 5920 4508 7288 4536
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 3476 4440 3521 4468
rect 3476 4428 3482 4440
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 4157 4471 4215 4477
rect 4157 4468 4169 4471
rect 3752 4440 4169 4468
rect 3752 4428 3758 4440
rect 4157 4437 4169 4440
rect 4203 4437 4215 4471
rect 4157 4431 4215 4437
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 5920 4468 5948 4508
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 7852 4536 7880 4567
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 8812 4576 9781 4604
rect 8812 4564 8818 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 9493 4539 9551 4545
rect 9493 4536 9505 4539
rect 7524 4508 7880 4536
rect 7944 4508 9505 4536
rect 7524 4496 7530 4508
rect 4396 4440 5948 4468
rect 5997 4471 6055 4477
rect 4396 4428 4402 4440
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6270 4468 6276 4480
rect 6043 4440 6276 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 6454 4468 6460 4480
rect 6415 4440 6460 4468
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 7944 4468 7972 4508
rect 9493 4505 9505 4508
rect 9539 4505 9551 4539
rect 9493 4499 9551 4505
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 10686 4536 10692 4548
rect 10192 4508 10692 4536
rect 10192 4496 10198 4508
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 11716 4536 11744 4567
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 11848 4576 11893 4604
rect 11848 4564 11854 4576
rect 12452 4548 12480 4635
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4604 13139 4607
rect 13630 4604 13636 4616
rect 13127 4576 13636 4604
rect 13127 4573 13139 4576
rect 13081 4567 13139 4573
rect 13630 4564 13636 4576
rect 13688 4604 13694 4616
rect 14476 4613 14504 4644
rect 14550 4632 14556 4644
rect 14608 4632 14614 4684
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13688 4576 14473 4604
rect 13688 4564 13694 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14642 4604 14648 4616
rect 14603 4576 14648 4604
rect 14461 4567 14519 4573
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 14844 4604 14872 4712
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 16301 4743 16359 4749
rect 16301 4709 16313 4743
rect 16347 4740 16359 4743
rect 16942 4740 16948 4752
rect 16347 4712 16948 4740
rect 16347 4709 16359 4712
rect 16301 4703 16359 4709
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 14976 4644 16405 4672
rect 14976 4632 14982 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 19978 4672 19984 4684
rect 19939 4644 19984 4672
rect 16393 4635 16451 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 14844 4576 15761 4604
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16482 4604 16488 4616
rect 16255 4576 16488 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 17402 4604 17408 4616
rect 17083 4576 17408 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 12066 4536 12072 4548
rect 11716 4508 12072 4536
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 12434 4496 12440 4548
rect 12492 4496 12498 4548
rect 13354 4496 13360 4548
rect 13412 4536 13418 4548
rect 15470 4536 15476 4548
rect 13412 4508 15476 4536
rect 13412 4496 13418 4508
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 8938 4468 8944 4480
rect 6604 4440 7972 4468
rect 8899 4440 8944 4468
rect 6604 4428 6610 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 10413 4471 10471 4477
rect 10413 4437 10425 4471
rect 10459 4468 10471 4471
rect 12526 4468 12532 4480
rect 10459 4440 12532 4468
rect 10459 4437 10471 4440
rect 10413 4431 10471 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15252 4440 15297 4468
rect 15252 4428 15258 4440
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17589 4471 17647 4477
rect 17589 4468 17601 4471
rect 17184 4440 17601 4468
rect 17184 4428 17190 4440
rect 17589 4437 17601 4440
rect 17635 4437 17647 4471
rect 17589 4431 17647 4437
rect 20165 4471 20223 4477
rect 20165 4437 20177 4471
rect 20211 4468 20223 4471
rect 20990 4468 20996 4480
rect 20211 4440 20996 4468
rect 20211 4437 20223 4440
rect 20165 4431 20223 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3418 4264 3424 4276
rect 2740 4236 3424 4264
rect 2740 4224 2746 4236
rect 3418 4224 3424 4236
rect 3476 4224 3482 4276
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4264 4031 4267
rect 4338 4264 4344 4276
rect 4019 4236 4344 4264
rect 4019 4233 4031 4236
rect 3973 4227 4031 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4433 4267 4491 4273
rect 4433 4233 4445 4267
rect 4479 4264 4491 4267
rect 5626 4264 5632 4276
rect 4479 4236 5632 4264
rect 4479 4233 4491 4236
rect 4433 4227 4491 4233
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6457 4267 6515 4273
rect 6457 4264 6469 4267
rect 5868 4236 6469 4264
rect 5868 4224 5874 4236
rect 6457 4233 6469 4236
rect 6503 4233 6515 4267
rect 6457 4227 6515 4233
rect 8110 4224 8116 4276
rect 8168 4264 8174 4276
rect 9030 4264 9036 4276
rect 8168 4236 9036 4264
rect 8168 4224 8174 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 11054 4264 11060 4276
rect 9140 4236 11060 4264
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 2924 4168 3157 4196
rect 2924 4156 2930 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 3697 4199 3755 4205
rect 3191 4168 3648 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 3620 4128 3648 4168
rect 3697 4165 3709 4199
rect 3743 4196 3755 4199
rect 3743 4168 4844 4196
rect 3743 4165 3755 4168
rect 3697 4159 3755 4165
rect 4614 4128 4620 4140
rect 3160 4100 3556 4128
rect 3620 4100 4620 4128
rect 3160 4072 3188 4100
rect 1210 4020 1216 4072
rect 1268 4060 1274 4072
rect 1489 4063 1547 4069
rect 1489 4060 1501 4063
rect 1268 4032 1501 4060
rect 1268 4020 1274 4032
rect 1489 4029 1501 4032
rect 1535 4060 1547 4063
rect 1578 4060 1584 4072
rect 1535 4032 1584 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 3050 4020 3056 4072
rect 3108 4020 3114 4072
rect 3142 4020 3148 4072
rect 3200 4020 3206 4072
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3418 4060 3424 4072
rect 3283 4032 3424 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 3528 4069 3556 4100
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3694 4060 3700 4072
rect 3559 4032 3700 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 4062 4060 4068 4072
rect 3844 4032 3889 4060
rect 3975 4032 4068 4060
rect 3844 4020 3850 4032
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4816 4060 4844 4168
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 6270 4196 6276 4208
rect 6052 4168 6276 4196
rect 6052 4156 6058 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 6840 4168 7512 4196
rect 6840 4128 6868 4168
rect 5736 4100 6868 4128
rect 5736 4060 5764 4100
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6972 4100 7021 4128
rect 6972 4088 6978 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 4816 4032 5764 4060
rect 5813 4063 5871 4069
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5902 4060 5908 4072
rect 5859 4032 5908 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 6788 4032 7297 4060
rect 6788 4020 6794 4032
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7484 4060 7512 4168
rect 7576 4168 8524 4196
rect 7576 4137 7604 4168
rect 8496 4140 8524 4168
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 9140 4196 9168 4236
rect 11054 4224 11060 4236
rect 11112 4264 11118 4276
rect 12250 4264 12256 4276
rect 11112 4236 12256 4264
rect 11112 4224 11118 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13630 4264 13636 4276
rect 13136 4236 13492 4264
rect 13591 4236 13636 4264
rect 13136 4224 13142 4236
rect 8812 4168 9168 4196
rect 8812 4156 8818 4168
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 12342 4196 12348 4208
rect 9732 4168 10732 4196
rect 9732 4156 9738 4168
rect 10704 4140 10732 4168
rect 11992 4168 12348 4196
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 8294 4128 8300 4140
rect 7708 4100 8300 4128
rect 7708 4088 7714 4100
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8478 4128 8484 4140
rect 8439 4100 8484 4128
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 10226 4128 10232 4140
rect 9539 4100 10232 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10594 4128 10600 4140
rect 10555 4100 10600 4128
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10744 4100 10837 4128
rect 10744 4088 10750 4100
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11992 4137 12020 4168
rect 12342 4156 12348 4168
rect 12400 4196 12406 4208
rect 13354 4196 13360 4208
rect 12400 4168 13360 4196
rect 12400 4156 12406 4168
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 13464 4196 13492 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 15102 4264 15108 4276
rect 14108 4236 15108 4264
rect 14108 4196 14136 4236
rect 13464 4168 14136 4196
rect 11425 4131 11483 4137
rect 11425 4128 11437 4131
rect 11020 4100 11437 4128
rect 11020 4088 11026 4100
rect 11425 4097 11437 4100
rect 11471 4097 11483 4131
rect 11425 4091 11483 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4097 12035 4131
rect 12434 4128 12440 4140
rect 11977 4091 12035 4097
rect 12176 4100 12440 4128
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7484 4032 7757 4060
rect 7285 4023 7343 4029
rect 7745 4029 7757 4032
rect 7791 4060 7803 4063
rect 8662 4060 8668 4072
rect 7791 4032 8432 4060
rect 8623 4032 8668 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 2038 4001 2044 4004
rect 2032 3955 2044 4001
rect 2096 3992 2102 4004
rect 3068 3992 3096 4020
rect 4080 3992 4108 4020
rect 2096 3964 2132 3992
rect 3068 3964 3464 3992
rect 2038 3952 2044 3955
rect 2096 3952 2102 3964
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 2590 3924 2596 3936
rect 1627 3896 2596 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3326 3924 3332 3936
rect 3108 3896 3332 3924
rect 3108 3884 3114 3896
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3436 3933 3464 3964
rect 3528 3964 4108 3992
rect 3528 3936 3556 3964
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5546 3995 5604 4001
rect 5546 3992 5558 3995
rect 4764 3964 5558 3992
rect 4764 3952 4770 3964
rect 5546 3961 5558 3964
rect 5592 3961 5604 3995
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 5546 3955 5604 3961
rect 5644 3964 6193 3992
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 3510 3884 3516 3936
rect 3568 3884 3574 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4982 3924 4988 3936
rect 4295 3896 4988 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5644 3924 5672 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 6270 3952 6276 4004
rect 6328 3992 6334 4004
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 6328 3964 6929 3992
rect 6328 3952 6334 3964
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 8110 3992 8116 4004
rect 7432 3964 8116 3992
rect 7432 3952 7438 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 5902 3924 5908 3936
rect 5132 3896 5672 3924
rect 5863 3896 5908 3924
rect 5132 3884 5138 3896
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 6822 3924 6828 3936
rect 6783 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7837 3927 7895 3933
rect 7837 3924 7849 3927
rect 7340 3896 7849 3924
rect 7340 3884 7346 3896
rect 7837 3893 7849 3896
rect 7883 3893 7895 3927
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 7837 3887 7895 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8404 3924 8432 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 12176 4069 12204 4100
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 13262 4128 13268 4140
rect 13223 4100 13268 4128
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 15028 4137 15056 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 8864 4032 12173 4060
rect 8573 3995 8631 4001
rect 8573 3961 8585 3995
rect 8619 3992 8631 3995
rect 8754 3992 8760 4004
rect 8619 3964 8760 3992
rect 8619 3961 8631 3964
rect 8573 3955 8631 3961
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 8864 3924 8892 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 12250 4020 12256 4072
rect 12308 4060 12314 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12308 4032 12817 4060
rect 12308 4020 12314 4032
rect 12805 4029 12817 4032
rect 12851 4060 12863 4063
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12851 4032 13093 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13081 4029 13093 4032
rect 13127 4029 13139 4063
rect 14918 4060 14924 4072
rect 13081 4023 13139 4029
rect 14476 4032 14924 4060
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 10505 3995 10563 4001
rect 9723 3964 10180 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 9030 3924 9036 3936
rect 8404 3896 8892 3924
rect 8991 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9585 3927 9643 3933
rect 9180 3896 9225 3924
rect 9180 3884 9186 3896
rect 9585 3893 9597 3927
rect 9631 3924 9643 3927
rect 9858 3924 9864 3936
rect 9631 3896 9864 3924
rect 9631 3893 9643 3896
rect 9585 3887 9643 3893
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10152 3933 10180 3964
rect 10505 3961 10517 3995
rect 10551 3992 10563 3995
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 10551 3964 10977 3992
rect 10551 3961 10563 3964
rect 10505 3955 10563 3961
rect 10965 3961 10977 3964
rect 11011 3961 11023 3995
rect 14476 3992 14504 4032
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 10965 3955 11023 3961
rect 12544 3964 14504 3992
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 11112 3896 11253 3924
rect 11112 3884 11118 3896
rect 11241 3893 11253 3896
rect 11287 3893 11299 3927
rect 11241 3887 11299 3893
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12544 3933 12572 3964
rect 14734 3952 14740 4004
rect 14792 4001 14798 4004
rect 14792 3992 14804 4001
rect 14792 3964 14837 3992
rect 14792 3955 14804 3964
rect 14792 3952 14798 3955
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 12032 3896 12081 3924
rect 12032 3884 12038 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12529 3927 12587 3933
rect 12529 3893 12541 3927
rect 12575 3893 12587 3927
rect 12529 3887 12587 3893
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 12710 3924 12716 3936
rect 12667 3896 12716 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14366 3884 14372 3936
rect 14424 3924 14430 3936
rect 15105 3927 15163 3933
rect 15105 3924 15117 3927
rect 14424 3896 15117 3924
rect 14424 3884 14430 3896
rect 15105 3893 15117 3896
rect 15151 3893 15163 3927
rect 15105 3887 15163 3893
rect 17313 3927 17371 3933
rect 17313 3893 17325 3927
rect 17359 3924 17371 3927
rect 18046 3924 18052 3936
rect 17359 3896 18052 3924
rect 17359 3893 17371 3896
rect 17313 3887 17371 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 2498 3720 2504 3732
rect 1627 3692 2504 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3786 3720 3792 3732
rect 3016 3692 3792 3720
rect 3016 3680 3022 3692
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4798 3720 4804 3732
rect 4028 3692 4804 3720
rect 4028 3680 4034 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5868 3692 6193 3720
rect 5868 3680 5874 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 6549 3723 6607 3729
rect 6549 3689 6561 3723
rect 6595 3720 6607 3723
rect 6914 3720 6920 3732
rect 6595 3692 6920 3720
rect 6595 3689 6607 3692
rect 6549 3683 6607 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7055 3692 7512 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 2774 3652 2780 3664
rect 2832 3661 2838 3664
rect 2832 3655 2866 3661
rect 2718 3624 2780 3652
rect 2774 3612 2780 3624
rect 2854 3652 2866 3655
rect 3050 3652 3056 3664
rect 2854 3624 3056 3652
rect 2854 3621 2866 3624
rect 2832 3615 2866 3621
rect 2832 3612 2838 3615
rect 3050 3612 3056 3624
rect 3108 3652 3114 3664
rect 3694 3652 3700 3664
rect 3108 3624 3700 3652
rect 3108 3612 3114 3624
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 4148 3655 4206 3661
rect 4148 3621 4160 3655
rect 4194 3652 4206 3655
rect 4614 3652 4620 3664
rect 4194 3624 4620 3652
rect 4194 3621 4206 3624
rect 4148 3615 4206 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 4706 3612 4712 3664
rect 4764 3652 4770 3664
rect 5353 3655 5411 3661
rect 5353 3652 5365 3655
rect 4764 3624 5365 3652
rect 4764 3612 4770 3624
rect 5353 3621 5365 3624
rect 5399 3621 5411 3655
rect 7484 3652 7512 3692
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7616 3692 7941 3720
rect 7616 3680 7622 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 8478 3720 8484 3732
rect 8352 3692 8484 3720
rect 8352 3680 8358 3692
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8628 3692 8769 3720
rect 8628 3680 8634 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 8757 3683 8815 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 9088 3692 9505 3720
rect 9088 3680 9094 3692
rect 9493 3689 9505 3692
rect 9539 3689 9551 3723
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 9493 3683 9551 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 11882 3720 11888 3732
rect 10100 3692 11888 3720
rect 10100 3680 10106 3692
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12066 3720 12072 3732
rect 12027 3692 12072 3720
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12158 3680 12164 3732
rect 12216 3680 12222 3732
rect 13357 3723 13415 3729
rect 13357 3689 13369 3723
rect 13403 3689 13415 3723
rect 14090 3720 14096 3732
rect 14051 3692 14096 3720
rect 13357 3683 13415 3689
rect 8018 3652 8024 3664
rect 7484 3624 8024 3652
rect 5353 3615 5411 3621
rect 8018 3612 8024 3624
rect 8076 3612 8082 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 9401 3655 9459 3661
rect 9401 3652 9413 3655
rect 8260 3624 9413 3652
rect 8260 3612 8266 3624
rect 9401 3621 9413 3624
rect 9447 3621 9459 3655
rect 9401 3615 9459 3621
rect 9646 3624 10548 3652
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1397 3587 1455 3593
rect 1397 3584 1409 3587
rect 1360 3556 1409 3584
rect 1360 3544 1366 3556
rect 1397 3553 1409 3556
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 3142 3584 3148 3596
rect 2556 3556 3148 3584
rect 2556 3544 2562 3556
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3584 3295 3587
rect 3326 3584 3332 3596
rect 3283 3556 3332 3584
rect 3283 3553 3295 3556
rect 3237 3547 3295 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3881 3587 3939 3593
rect 3881 3584 3893 3587
rect 3436 3556 3893 3584
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3436 3516 3464 3556
rect 3881 3553 3893 3556
rect 3927 3584 3939 3587
rect 4522 3584 4528 3596
rect 3927 3556 4528 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 4948 3556 5825 3584
rect 4948 3544 4954 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 6288 3556 6500 3584
rect 3099 3488 3464 3516
rect 3513 3519 3571 3525
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3513 3485 3525 3519
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5537 3479 5595 3485
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 6288 3516 6316 3556
rect 5767 3488 6316 3516
rect 6365 3519 6423 3525
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 3528 3448 3556 3479
rect 3786 3448 3792 3460
rect 3528 3420 3792 3448
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 5353 3451 5411 3457
rect 5353 3448 5365 3451
rect 5307 3420 5365 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 5353 3417 5365 3420
rect 5399 3448 5411 3451
rect 5552 3448 5580 3479
rect 5626 3448 5632 3460
rect 5399 3420 5632 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 5626 3408 5632 3420
rect 5684 3448 5690 3460
rect 6380 3448 6408 3479
rect 5684 3420 6408 3448
rect 6472 3448 6500 3556
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6604 3556 6653 3584
rect 6604 3544 6610 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 6641 3547 6699 3553
rect 6932 3556 7297 3584
rect 6730 3476 6736 3528
rect 6788 3516 6794 3528
rect 6932 3516 6960 3556
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 7285 3547 7343 3553
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7524 3556 8524 3584
rect 7524 3544 7530 3556
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 6788 3488 6960 3516
rect 7024 3488 8033 3516
rect 6788 3476 6794 3488
rect 6472 3420 6684 3448
rect 5684 3408 5690 3420
rect 1670 3380 1676 3392
rect 1631 3352 1676 3380
rect 1670 3340 1676 3352
rect 1728 3380 1734 3392
rect 1946 3380 1952 3392
rect 1728 3352 1952 3380
rect 1728 3340 1734 3352
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2866 3380 2872 3392
rect 2096 3352 2872 3380
rect 2096 3340 2102 3352
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3329 3383 3387 3389
rect 3329 3380 3341 3383
rect 3292 3352 3341 3380
rect 3292 3340 3298 3352
rect 3329 3349 3341 3352
rect 3375 3349 3387 3383
rect 6656 3380 6684 3420
rect 6822 3408 6828 3460
rect 6880 3448 6886 3460
rect 7024 3448 7052 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8294 3516 8300 3528
rect 8251 3488 8300 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 6880 3420 7052 3448
rect 7101 3451 7159 3457
rect 6880 3408 6886 3420
rect 7101 3417 7113 3451
rect 7147 3448 7159 3451
rect 7742 3448 7748 3460
rect 7147 3420 7748 3448
rect 7147 3417 7159 3420
rect 7101 3411 7159 3417
rect 7116 3380 7144 3411
rect 7742 3408 7748 3420
rect 7800 3408 7806 3460
rect 8036 3448 8064 3479
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8496 3516 8524 3556
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 8628 3556 8677 3584
rect 8628 3544 8634 3556
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 9646 3584 9674 3624
rect 10134 3584 10140 3596
rect 8665 3547 8723 3553
rect 9140 3556 9674 3584
rect 10095 3556 10140 3584
rect 9140 3516 9168 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 10393 3587 10451 3593
rect 10393 3584 10405 3587
rect 10284 3556 10405 3584
rect 10284 3544 10290 3556
rect 10393 3553 10405 3556
rect 10439 3553 10451 3587
rect 10520 3584 10548 3624
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 10520 3556 11989 3584
rect 10393 3547 10451 3553
rect 11977 3553 11989 3556
rect 12023 3584 12035 3587
rect 12176 3584 12204 3680
rect 13372 3652 13400 3683
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14642 3720 14648 3732
rect 14415 3692 14648 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 18325 3723 18383 3729
rect 18325 3720 18337 3723
rect 18196 3692 18337 3720
rect 18196 3680 18202 3692
rect 18325 3689 18337 3692
rect 18371 3689 18383 3723
rect 18325 3683 18383 3689
rect 12544 3624 13400 3652
rect 12434 3584 12440 3596
rect 12023 3556 12204 3584
rect 12395 3556 12440 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 8496 3488 9168 3516
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9272 3488 9321 3516
rect 9272 3476 9278 3488
rect 9309 3485 9321 3488
rect 9355 3516 9367 3519
rect 9582 3516 9588 3528
rect 9355 3488 9588 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11940 3488 12173 3516
rect 11940 3476 11946 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12544 3516 12572 3624
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14829 3655 14887 3661
rect 14829 3652 14841 3655
rect 14056 3624 14841 3652
rect 14056 3612 14062 3624
rect 14829 3621 14841 3624
rect 14875 3652 14887 3655
rect 15562 3652 15568 3664
rect 14875 3624 15568 3652
rect 14875 3621 14887 3624
rect 14829 3615 14887 3621
rect 15562 3612 15568 3624
rect 15620 3652 15626 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15620 3624 16037 3652
rect 15620 3612 15626 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 20162 3652 20168 3664
rect 16025 3615 16083 3621
rect 17880 3624 20168 3652
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12400 3488 12572 3516
rect 12636 3556 12817 3584
rect 12400 3476 12406 3488
rect 9766 3448 9772 3460
rect 8036 3420 9772 3448
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 12636 3457 12664 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 13078 3584 13084 3596
rect 13039 3556 13084 3584
rect 12805 3547 12863 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 13556 3516 13584 3547
rect 14090 3544 14096 3596
rect 14148 3584 14154 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14148 3556 14749 3584
rect 14148 3544 14154 3556
rect 14737 3553 14749 3556
rect 14783 3584 14795 3587
rect 15378 3584 15384 3596
rect 14783 3556 15240 3584
rect 15339 3556 15384 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 12820 3488 13829 3516
rect 12820 3460 12848 3488
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 14918 3516 14924 3528
rect 14879 3488 14924 3516
rect 13817 3479 13875 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 15212 3516 15240 3556
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 17880 3584 17908 3624
rect 20162 3612 20168 3624
rect 20220 3612 20226 3664
rect 18046 3584 18052 3596
rect 15580 3556 17908 3584
rect 18007 3556 18052 3584
rect 15580 3516 15608 3556
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 15212 3488 15608 3516
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 11164 3420 11621 3448
rect 11164 3392 11192 3420
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 12621 3451 12679 3457
rect 12621 3417 12633 3451
rect 12667 3417 12679 3451
rect 12621 3411 12679 3417
rect 12802 3408 12808 3460
rect 12860 3408 12866 3460
rect 14274 3408 14280 3460
rect 14332 3448 14338 3460
rect 15197 3451 15255 3457
rect 15197 3448 15209 3451
rect 14332 3420 15209 3448
rect 14332 3408 14338 3420
rect 15197 3417 15209 3420
rect 15243 3417 15255 3451
rect 15197 3411 15255 3417
rect 15378 3408 15384 3460
rect 15436 3448 15442 3460
rect 15565 3451 15623 3457
rect 15565 3448 15577 3451
rect 15436 3420 15577 3448
rect 15436 3408 15442 3420
rect 15565 3417 15577 3420
rect 15611 3417 15623 3451
rect 15565 3411 15623 3417
rect 18233 3451 18291 3457
rect 18233 3417 18245 3451
rect 18279 3448 18291 3451
rect 19150 3448 19156 3460
rect 18279 3420 19156 3448
rect 18279 3417 18291 3420
rect 18233 3411 18291 3417
rect 19150 3408 19156 3420
rect 19208 3408 19214 3460
rect 6656 3352 7144 3380
rect 3329 3343 3387 3349
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 7561 3383 7619 3389
rect 7561 3380 7573 3383
rect 7524 3352 7573 3380
rect 7524 3340 7530 3352
rect 7561 3349 7573 3352
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8570 3380 8576 3392
rect 8527 3352 8576 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9953 3383 10011 3389
rect 9953 3380 9965 3383
rect 9640 3352 9965 3380
rect 9640 3340 9646 3352
rect 9953 3349 9965 3352
rect 9999 3349 10011 3383
rect 9953 3343 10011 3349
rect 11146 3340 11152 3392
rect 11204 3340 11210 3392
rect 11517 3383 11575 3389
rect 11517 3349 11529 3383
rect 11563 3380 11575 3383
rect 12158 3380 12164 3392
rect 11563 3352 12164 3380
rect 11563 3349 11575 3352
rect 11517 3343 11575 3349
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12986 3380 12992 3392
rect 12947 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13262 3380 13268 3392
rect 13223 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 13633 3383 13691 3389
rect 13633 3380 13645 3383
rect 13596 3352 13645 3380
rect 13596 3340 13602 3352
rect 13633 3349 13645 3352
rect 13679 3349 13691 3383
rect 13633 3343 13691 3349
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 15841 3383 15899 3389
rect 15841 3380 15853 3383
rect 15804 3352 15853 3380
rect 15804 3340 15810 3352
rect 15841 3349 15853 3352
rect 15887 3349 15899 3383
rect 15841 3343 15899 3349
rect 19058 3340 19064 3392
rect 19116 3380 19122 3392
rect 19702 3380 19708 3392
rect 19116 3352 19708 3380
rect 19116 3340 19122 3352
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 2682 3176 2688 3188
rect 1636 3148 2688 3176
rect 1636 3136 1642 3148
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 3513 3179 3571 3185
rect 3513 3145 3525 3179
rect 3559 3176 3571 3179
rect 3559 3148 4108 3176
rect 3559 3145 3571 3148
rect 3513 3139 3571 3145
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 3970 3108 3976 3120
rect 1719 3080 3976 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 2406 3040 2412 3052
rect 1504 3012 2412 3040
rect 1504 2984 1532 3012
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2774 3040 2780 3052
rect 2639 3012 2780 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2774 3000 2780 3012
rect 2832 3040 2838 3052
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2832 3012 2881 3040
rect 2832 3000 2838 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 3068 3040 3096 3080
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 3068 3012 3188 3040
rect 2869 3003 2927 3009
rect 1486 2972 1492 2984
rect 1399 2944 1492 2972
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 2314 2972 2320 2984
rect 2275 2944 2320 2972
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 3160 2981 3188 3012
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 3844 3012 3889 3040
rect 3844 3000 3850 3012
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2941 3203 2975
rect 4080 2972 4108 3148
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4212 3148 5273 3176
rect 4212 3136 4218 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 6270 3176 6276 3188
rect 6227 3148 6276 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7469 3179 7527 3185
rect 7469 3176 7481 3179
rect 7432 3148 7481 3176
rect 7432 3136 7438 3148
rect 7469 3145 7481 3148
rect 7515 3176 7527 3179
rect 9214 3176 9220 3188
rect 7515 3148 9220 3176
rect 7515 3145 7527 3148
rect 7469 3139 7527 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10226 3176 10232 3188
rect 9732 3148 10232 3176
rect 9732 3136 9738 3148
rect 10226 3136 10232 3148
rect 10284 3176 10290 3188
rect 10321 3179 10379 3185
rect 10321 3176 10333 3179
rect 10284 3148 10333 3176
rect 10284 3136 10290 3148
rect 10321 3145 10333 3148
rect 10367 3145 10379 3179
rect 10321 3139 10379 3145
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10468 3148 10609 3176
rect 10468 3136 10474 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11756 3148 11897 3176
rect 11756 3136 11762 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 13633 3179 13691 3185
rect 13633 3145 13645 3179
rect 13679 3176 13691 3179
rect 14918 3176 14924 3188
rect 13679 3148 14924 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15749 3179 15807 3185
rect 15436 3148 15700 3176
rect 15436 3136 15442 3148
rect 4246 3068 4252 3120
rect 4304 3108 4310 3120
rect 4433 3111 4491 3117
rect 4433 3108 4445 3111
rect 4304 3080 4445 3108
rect 4304 3068 4310 3080
rect 4433 3077 4445 3080
rect 4479 3077 4491 3111
rect 4433 3071 4491 3077
rect 6086 3068 6092 3120
rect 6144 3108 6150 3120
rect 6457 3111 6515 3117
rect 6457 3108 6469 3111
rect 6144 3080 6469 3108
rect 6144 3068 6150 3080
rect 6457 3077 6469 3080
rect 6503 3077 6515 3111
rect 7282 3108 7288 3120
rect 6457 3071 6515 3077
rect 6840 3080 7288 3108
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5626 3040 5632 3052
rect 5040 3012 5085 3040
rect 5587 3012 5632 3040
rect 5040 3000 5046 3012
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3040 5779 3043
rect 6840 3040 6868 3080
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 14829 3111 14887 3117
rect 10192 3080 12296 3108
rect 10192 3068 10198 3080
rect 5767 3012 6868 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 6972 3012 7113 3040
rect 6972 3000 6978 3012
rect 7101 3009 7113 3012
rect 7147 3009 7159 3043
rect 8846 3040 8852 3052
rect 8759 3012 8852 3040
rect 7101 3003 7159 3009
rect 8846 3000 8852 3012
rect 8904 3040 8910 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8904 3012 8953 3040
rect 8904 3000 8910 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 10284 3012 11345 3040
rect 10284 3000 10290 3012
rect 11333 3009 11345 3012
rect 11379 3040 11391 3043
rect 11882 3040 11888 3052
rect 11379 3012 11888 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12268 3049 12296 3080
rect 14829 3077 14841 3111
rect 14875 3108 14887 3111
rect 15470 3108 15476 3120
rect 14875 3080 15476 3108
rect 14875 3077 14887 3080
rect 14829 3071 14887 3077
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 15672 3108 15700 3148
rect 15749 3145 15761 3179
rect 15795 3176 15807 3179
rect 16758 3176 16764 3188
rect 15795 3148 16764 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 20993 3179 21051 3185
rect 20993 3176 21005 3179
rect 16908 3148 21005 3176
rect 16908 3136 16914 3148
rect 20993 3145 21005 3148
rect 21039 3145 21051 3179
rect 20993 3139 21051 3145
rect 16025 3111 16083 3117
rect 15672 3080 15976 3108
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 13262 3000 13268 3052
rect 13320 3040 13326 3052
rect 13320 3012 14044 3040
rect 13320 3000 13326 3012
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 4080 2944 4813 2972
rect 3145 2935 3203 2941
rect 4801 2941 4813 2944
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 5994 2972 6000 2984
rect 5859 2944 6000 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 9214 2981 9220 2984
rect 9208 2972 9220 2981
rect 9175 2944 9220 2972
rect 9208 2935 9220 2944
rect 9214 2932 9220 2935
rect 9272 2932 9278 2984
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 10318 2972 10324 2984
rect 9640 2944 10324 2972
rect 9640 2932 9646 2944
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 11149 2975 11207 2981
rect 10560 2944 10605 2972
rect 10560 2932 10566 2944
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11238 2972 11244 2984
rect 11195 2944 11244 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11480 2944 12081 2972
rect 11480 2932 11486 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12342 2972 12348 2984
rect 12216 2944 12348 2972
rect 12216 2932 12222 2944
rect 12342 2932 12348 2944
rect 12400 2972 12406 2984
rect 12509 2975 12567 2981
rect 12509 2972 12521 2975
rect 12400 2944 12521 2972
rect 12400 2932 12406 2944
rect 12509 2941 12521 2944
rect 12555 2941 12567 2975
rect 12509 2935 12567 2941
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 14016 2981 14044 3012
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 15746 3040 15752 3052
rect 14424 3012 14964 3040
rect 14424 3000 14430 3012
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13412 2944 13737 2972
rect 13412 2932 13418 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2941 14059 2975
rect 14274 2972 14280 2984
rect 14235 2944 14280 2972
rect 14001 2935 14059 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14936 2981 14964 3012
rect 15304 3012 15752 3040
rect 15304 2981 15332 3012
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2941 15347 2975
rect 15562 2972 15568 2984
rect 15523 2944 15568 2972
rect 15289 2935 15347 2941
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 4356 2876 4905 2904
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1302 2836 1308 2848
rect 256 2808 1308 2836
rect 256 2796 262 2808
rect 1302 2796 1308 2808
rect 1360 2836 1366 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 1360 2808 1777 2836
rect 1360 2796 1366 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1946 2836 1952 2848
rect 1907 2808 1952 2836
rect 1765 2799 1823 2805
rect 1946 2796 1952 2808
rect 2004 2796 2010 2848
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3694 2836 3700 2848
rect 3099 2808 3700 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 3881 2839 3939 2845
rect 3881 2836 3893 2839
rect 3844 2808 3893 2836
rect 3844 2796 3850 2808
rect 3881 2805 3893 2808
rect 3927 2805 3939 2839
rect 3881 2799 3939 2805
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4246 2836 4252 2848
rect 4019 2808 4252 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 4356 2845 4384 2876
rect 4893 2873 4905 2876
rect 4939 2873 4951 2907
rect 4893 2867 4951 2873
rect 5442 2864 5448 2916
rect 5500 2904 5506 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 5500 2876 7297 2904
rect 5500 2864 5506 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 8018 2864 8024 2916
rect 8076 2864 8082 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8582 2907 8640 2913
rect 8582 2904 8594 2907
rect 8352 2876 8594 2904
rect 8352 2864 8358 2876
rect 8582 2873 8594 2876
rect 8628 2904 8640 2907
rect 8754 2904 8760 2916
rect 8628 2876 8760 2904
rect 8628 2873 8640 2876
rect 8582 2867 8640 2873
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 10226 2904 10232 2916
rect 9508 2876 10232 2904
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2805 4399 2839
rect 4341 2799 4399 2805
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 5534 2836 5540 2848
rect 4672 2808 5540 2836
rect 4672 2796 4678 2808
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6546 2796 6552 2848
rect 6604 2836 6610 2848
rect 6825 2839 6883 2845
rect 6825 2836 6837 2839
rect 6604 2808 6837 2836
rect 6604 2796 6610 2808
rect 6825 2805 6837 2808
rect 6871 2805 6883 2839
rect 6825 2799 6883 2805
rect 6917 2839 6975 2845
rect 6917 2805 6929 2839
rect 6963 2836 6975 2839
rect 8036 2836 8064 2864
rect 9508 2848 9536 2876
rect 10226 2864 10232 2876
rect 10284 2864 10290 2916
rect 10962 2904 10968 2916
rect 10520 2876 10968 2904
rect 10520 2848 10548 2876
rect 10962 2864 10968 2876
rect 11020 2904 11026 2916
rect 11793 2907 11851 2913
rect 11793 2904 11805 2907
rect 11020 2876 11805 2904
rect 11020 2864 11026 2876
rect 11793 2873 11805 2876
rect 11839 2873 11851 2907
rect 15304 2904 15332 2935
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 15654 2932 15660 2984
rect 15712 2972 15718 2984
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15712 2944 15853 2972
rect 15712 2932 15718 2944
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15948 2972 15976 3080
rect 16025 3077 16037 3111
rect 16071 3077 16083 3111
rect 16025 3071 16083 3077
rect 16393 3111 16451 3117
rect 16393 3077 16405 3111
rect 16439 3108 16451 3111
rect 16942 3108 16948 3120
rect 16439 3080 16948 3108
rect 16439 3077 16451 3080
rect 16393 3071 16451 3077
rect 16040 3040 16068 3071
rect 16942 3068 16948 3080
rect 17000 3068 17006 3120
rect 17313 3111 17371 3117
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 17954 3108 17960 3120
rect 17359 3080 17960 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18785 3111 18843 3117
rect 18785 3077 18797 3111
rect 18831 3108 18843 3111
rect 19518 3108 19524 3120
rect 18831 3080 19524 3108
rect 18831 3077 18843 3080
rect 18785 3071 18843 3077
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 19978 3108 19984 3120
rect 19659 3080 19984 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 20162 3108 20168 3120
rect 20123 3080 20168 3108
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 16040 3012 18736 3040
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 15948 2944 16221 2972
rect 15841 2935 15899 2941
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16209 2935 16267 2941
rect 16390 2932 16396 2984
rect 16448 2972 16454 2984
rect 16485 2975 16543 2981
rect 16485 2972 16497 2975
rect 16448 2944 16497 2972
rect 16448 2932 16454 2944
rect 16485 2941 16497 2944
rect 16531 2972 16543 2975
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 16531 2944 16957 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17129 2975 17187 2981
rect 17129 2972 17141 2975
rect 17092 2944 17141 2972
rect 17092 2932 17098 2944
rect 17129 2941 17141 2944
rect 17175 2941 17187 2975
rect 17681 2975 17739 2981
rect 17681 2972 17693 2975
rect 17129 2935 17187 2941
rect 17236 2944 17693 2972
rect 17236 2904 17264 2944
rect 17681 2941 17693 2944
rect 17727 2941 17739 2975
rect 17862 2972 17868 2984
rect 17823 2944 17868 2972
rect 17681 2935 17739 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 18196 2944 18337 2972
rect 18196 2932 18202 2944
rect 18325 2941 18337 2944
rect 18371 2941 18383 2975
rect 18598 2972 18604 2984
rect 18559 2944 18604 2972
rect 18325 2935 18383 2941
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 17494 2904 17500 2916
rect 11793 2867 11851 2873
rect 12406 2876 15332 2904
rect 16684 2876 17264 2904
rect 17455 2876 17500 2904
rect 6963 2808 8064 2836
rect 6963 2805 6975 2808
rect 6917 2799 6975 2805
rect 9490 2796 9496 2848
rect 9548 2796 9554 2848
rect 10502 2796 10508 2848
rect 10560 2796 10566 2848
rect 10778 2836 10784 2848
rect 10739 2808 10784 2836
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11241 2839 11299 2845
rect 11241 2836 11253 2839
rect 10928 2808 11253 2836
rect 10928 2796 10934 2808
rect 11241 2805 11253 2808
rect 11287 2836 11299 2839
rect 12406 2836 12434 2876
rect 13906 2836 13912 2848
rect 11287 2808 12434 2836
rect 13867 2808 13912 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14274 2836 14280 2848
rect 14231 2808 14280 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14458 2836 14464 2848
rect 14419 2808 14464 2836
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 15105 2839 15163 2845
rect 15105 2805 15117 2839
rect 15151 2836 15163 2839
rect 15378 2836 15384 2848
rect 15151 2808 15384 2836
rect 15151 2805 15163 2808
rect 15105 2799 15163 2805
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2836 15531 2839
rect 15654 2836 15660 2848
rect 15519 2808 15660 2836
rect 15519 2805 15531 2808
rect 15473 2799 15531 2805
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 16684 2845 16712 2876
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 17880 2904 17908 2932
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 17880 2876 18429 2904
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 18417 2867 18475 2873
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2805 16727 2839
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 16669 2799 16727 2805
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 18616 2836 18644 2932
rect 18708 2904 18736 3012
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 18932 3012 19196 3040
rect 18932 3000 18938 3012
rect 19058 2972 19064 2984
rect 19019 2944 19064 2972
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19168 2972 19196 3012
rect 19242 3000 19248 3052
rect 19300 3040 19306 3052
rect 22186 3040 22192 3052
rect 19300 3012 22192 3040
rect 19300 3000 19306 3012
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 19429 2975 19487 2981
rect 19429 2972 19441 2975
rect 19168 2944 19441 2972
rect 19429 2941 19441 2944
rect 19475 2972 19487 2975
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 19475 2944 19901 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 20349 2975 20407 2981
rect 20349 2972 20361 2975
rect 20220 2944 20361 2972
rect 20220 2932 20226 2944
rect 20349 2941 20361 2944
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 20901 2975 20959 2981
rect 20901 2941 20913 2975
rect 20947 2972 20959 2975
rect 21177 2975 21235 2981
rect 21177 2972 21189 2975
rect 20947 2944 21189 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 21177 2941 21189 2944
rect 21223 2972 21235 2975
rect 22646 2972 22652 2984
rect 21223 2944 22652 2972
rect 21223 2941 21235 2944
rect 21177 2935 21235 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 21361 2907 21419 2913
rect 21361 2904 21373 2907
rect 18708 2876 21373 2904
rect 21361 2873 21373 2876
rect 21407 2873 21419 2907
rect 21361 2867 21419 2873
rect 21545 2907 21603 2913
rect 21545 2873 21557 2907
rect 21591 2904 21603 2907
rect 21726 2904 21732 2916
rect 21591 2876 21732 2904
rect 21591 2873 21603 2876
rect 21545 2867 21603 2873
rect 21726 2864 21732 2876
rect 21784 2864 21790 2916
rect 18877 2839 18935 2845
rect 18877 2836 18889 2839
rect 18196 2808 18241 2836
rect 18616 2808 18889 2836
rect 18196 2796 18202 2808
rect 18877 2805 18889 2808
rect 18923 2805 18935 2839
rect 18877 2799 18935 2805
rect 19245 2839 19303 2845
rect 19245 2805 19257 2839
rect 19291 2836 19303 2839
rect 19426 2836 19432 2848
rect 19291 2808 19432 2836
rect 19291 2805 19303 2808
rect 19245 2799 19303 2805
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 19702 2836 19708 2848
rect 19663 2808 19708 2836
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 20533 2839 20591 2845
rect 20533 2805 20545 2839
rect 20579 2836 20591 2839
rect 20714 2836 20720 2848
rect 20579 2808 20720 2836
rect 20579 2805 20591 2808
rect 20533 2799 20591 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 1811 2604 2237 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 3510 2632 3516 2644
rect 2639 2604 3516 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3660 2604 3985 2632
rect 3660 2592 3666 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4062 2592 4068 2644
rect 4120 2592 4126 2644
rect 4246 2592 4252 2644
rect 4304 2592 4310 2644
rect 4614 2632 4620 2644
rect 4575 2604 4620 2632
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4948 2604 4997 2632
rect 4948 2592 4954 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 5258 2632 5264 2644
rect 5219 2604 5264 2632
rect 4985 2595 5043 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5902 2632 5908 2644
rect 5863 2604 5908 2632
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 6546 2632 6552 2644
rect 6319 2604 6552 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7561 2635 7619 2641
rect 7561 2601 7573 2635
rect 7607 2632 7619 2635
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7607 2604 8033 2632
rect 7607 2601 7619 2604
rect 7561 2595 7619 2601
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8021 2595 8079 2601
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 9214 2632 9220 2644
rect 9175 2604 9220 2632
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9398 2592 9404 2644
rect 9456 2592 9462 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10321 2635 10379 2641
rect 10321 2632 10333 2635
rect 9815 2604 10333 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10321 2601 10333 2604
rect 10367 2601 10379 2635
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10321 2595 10379 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11974 2632 11980 2644
rect 11287 2604 11980 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12253 2635 12311 2641
rect 12253 2632 12265 2635
rect 12216 2604 12265 2632
rect 12216 2592 12222 2604
rect 12253 2601 12265 2604
rect 12299 2601 12311 2635
rect 12253 2595 12311 2601
rect 12621 2635 12679 2641
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 13078 2632 13084 2644
rect 12667 2604 13084 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 14369 2635 14427 2641
rect 13228 2604 13273 2632
rect 13228 2592 13234 2604
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14642 2632 14648 2644
rect 14415 2604 14648 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17218 2632 17224 2644
rect 17083 2604 17224 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 18138 2632 18144 2644
rect 17696 2604 18144 2632
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 1946 2564 1952 2576
rect 1719 2536 1952 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 1946 2524 1952 2536
rect 2004 2524 2010 2576
rect 2685 2567 2743 2573
rect 2685 2533 2697 2567
rect 2731 2564 2743 2567
rect 3326 2564 3332 2576
rect 2731 2536 3332 2564
rect 2731 2533 2743 2536
rect 2685 2527 2743 2533
rect 3326 2524 3332 2536
rect 3384 2524 3390 2576
rect 3421 2567 3479 2573
rect 3421 2533 3433 2567
rect 3467 2564 3479 2567
rect 3694 2564 3700 2576
rect 3467 2536 3700 2564
rect 3467 2533 3479 2536
rect 3421 2527 3479 2533
rect 3694 2524 3700 2536
rect 3752 2564 3758 2576
rect 4080 2564 4108 2592
rect 3752 2536 4108 2564
rect 4264 2564 4292 2592
rect 4709 2567 4767 2573
rect 4264 2536 4384 2564
rect 3752 2524 3758 2536
rect 1118 2456 1124 2508
rect 1176 2496 1182 2508
rect 1176 2468 2774 2496
rect 1176 2456 1182 2468
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 1670 2428 1676 2440
rect 1627 2400 1676 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2130 2360 2136 2372
rect 2091 2332 2136 2360
rect 2130 2320 2136 2332
rect 2188 2320 2194 2372
rect 2746 2292 2774 2468
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 3200 2468 3249 2496
rect 3200 2456 3206 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3237 2459 3295 2465
rect 3605 2499 3663 2505
rect 3605 2465 3617 2499
rect 3651 2496 3663 2499
rect 3786 2496 3792 2508
rect 3651 2468 3792 2496
rect 3651 2465 3663 2468
rect 3605 2459 3663 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4062 2496 4068 2508
rect 4023 2468 4068 2496
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 4246 2496 4252 2508
rect 4207 2468 4252 2496
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 4356 2496 4384 2536
rect 4709 2533 4721 2567
rect 4755 2564 4767 2567
rect 5810 2564 5816 2576
rect 4755 2536 5672 2564
rect 5771 2536 5816 2564
rect 4755 2533 4767 2536
rect 4709 2527 4767 2533
rect 5074 2496 5080 2508
rect 4356 2468 4936 2496
rect 5035 2468 5080 2496
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 4798 2428 4804 2440
rect 3099 2400 4804 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4908 2360 4936 2468
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5644 2496 5672 2536
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 6822 2564 6828 2576
rect 6783 2536 6828 2564
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 9416 2564 9444 2592
rect 8435 2536 9444 2564
rect 10689 2567 10747 2573
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 10689 2533 10701 2567
rect 10735 2564 10747 2567
rect 11146 2564 11152 2576
rect 10735 2536 11152 2564
rect 10735 2533 10747 2536
rect 10689 2527 10747 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 12986 2524 12992 2576
rect 13044 2564 13050 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 13044 2536 13645 2564
rect 13044 2524 13050 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 13906 2524 13912 2576
rect 13964 2564 13970 2576
rect 14001 2567 14059 2573
rect 14001 2564 14013 2567
rect 13964 2536 14013 2564
rect 13964 2524 13970 2536
rect 14001 2533 14013 2536
rect 14047 2533 14059 2567
rect 14001 2527 14059 2533
rect 14274 2524 14280 2576
rect 14332 2564 14338 2576
rect 14737 2567 14795 2573
rect 14737 2564 14749 2567
rect 14332 2536 14749 2564
rect 14332 2524 14338 2536
rect 14737 2533 14749 2536
rect 14783 2533 14795 2567
rect 15470 2564 15476 2576
rect 15431 2536 15476 2564
rect 14737 2527 14795 2533
rect 15470 2524 15476 2536
rect 15528 2524 15534 2576
rect 15654 2524 15660 2576
rect 15712 2564 15718 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 15712 2536 16313 2564
rect 15712 2524 15718 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 16758 2564 16764 2576
rect 16719 2536 16764 2564
rect 16301 2527 16359 2533
rect 16758 2524 16764 2536
rect 16816 2524 16822 2576
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 17696 2573 17724 2604
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 17405 2567 17463 2573
rect 17405 2564 17417 2567
rect 17000 2536 17417 2564
rect 17000 2524 17006 2536
rect 17405 2533 17417 2536
rect 17451 2533 17463 2567
rect 17405 2527 17463 2533
rect 17681 2567 17739 2573
rect 17681 2533 17693 2567
rect 17727 2533 17739 2567
rect 17681 2527 17739 2533
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 18601 2567 18659 2573
rect 18601 2564 18613 2567
rect 18104 2536 18613 2564
rect 18104 2524 18110 2536
rect 18601 2533 18613 2536
rect 18647 2533 18659 2567
rect 19150 2564 19156 2576
rect 19111 2536 19156 2564
rect 18601 2527 18659 2533
rect 19150 2524 19156 2536
rect 19208 2524 19214 2576
rect 19518 2524 19524 2576
rect 19576 2564 19582 2576
rect 19613 2567 19671 2573
rect 19613 2564 19625 2567
rect 19576 2536 19625 2564
rect 19576 2524 19582 2536
rect 19613 2533 19625 2536
rect 19659 2533 19671 2567
rect 19613 2527 19671 2533
rect 19978 2524 19984 2576
rect 20036 2564 20042 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 20036 2536 20545 2564
rect 20036 2524 20042 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 20714 2524 20720 2576
rect 20772 2564 20778 2576
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 20772 2536 21465 2564
rect 20772 2524 20778 2536
rect 21453 2533 21465 2536
rect 21499 2533 21511 2567
rect 21453 2527 21511 2533
rect 6270 2496 6276 2508
rect 5644 2468 6276 2496
rect 6270 2456 6276 2468
rect 6328 2456 6334 2508
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 6641 2499 6699 2505
rect 6641 2496 6653 2499
rect 6512 2468 6653 2496
rect 6512 2456 6518 2468
rect 6641 2465 6653 2468
rect 6687 2465 6699 2499
rect 6641 2459 6699 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7098 2496 7104 2508
rect 6963 2468 7104 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8996 2468 9045 2496
rect 8996 2456 9002 2468
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9180 2468 9413 2496
rect 9180 2456 9186 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 5626 2428 5632 2440
rect 5587 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 8754 2428 8760 2440
rect 8711 2400 8760 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 8754 2388 8760 2400
rect 8812 2428 8818 2440
rect 9490 2428 9496 2440
rect 8812 2400 9496 2428
rect 8812 2388 8818 2400
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9732 2400 9777 2428
rect 9732 2388 9738 2400
rect 7929 2363 7987 2369
rect 4908 2332 7236 2360
rect 4154 2292 4160 2304
rect 2746 2264 4160 2292
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 6822 2292 6828 2304
rect 4479 2264 6828 2292
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7208 2292 7236 2332
rect 7929 2329 7941 2363
rect 7975 2360 7987 2363
rect 9876 2360 9904 2459
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 11330 2496 11336 2508
rect 10100 2468 11336 2496
rect 10100 2456 10106 2468
rect 11330 2456 11336 2468
rect 11388 2456 11394 2508
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2465 11759 2499
rect 12342 2496 12348 2508
rect 11701 2459 11759 2465
rect 12084 2468 12348 2496
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10836 2400 10885 2428
rect 10836 2388 10842 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11716 2428 11744 2459
rect 12084 2437 12112 2468
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 13265 2499 13323 2505
rect 13265 2465 13277 2499
rect 13311 2496 13323 2499
rect 13538 2496 13544 2508
rect 13311 2468 13544 2496
rect 13311 2465 13323 2468
rect 13265 2459 13323 2465
rect 11112 2400 11744 2428
rect 12069 2431 12127 2437
rect 11112 2388 11118 2400
rect 12069 2397 12081 2431
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2397 12219 2431
rect 13280 2428 13308 2459
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 14185 2499 14243 2505
rect 14185 2465 14197 2499
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 12161 2391 12219 2397
rect 12728 2400 13308 2428
rect 14200 2428 14228 2459
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 15105 2499 15163 2505
rect 15105 2496 15117 2499
rect 14516 2468 15117 2496
rect 14516 2456 14522 2468
rect 15105 2465 15117 2468
rect 15151 2465 15163 2499
rect 15105 2459 15163 2465
rect 15194 2456 15200 2508
rect 15252 2456 15258 2508
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15436 2468 15853 2496
rect 15436 2456 15442 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18141 2499 18199 2505
rect 18141 2496 18153 2499
rect 18012 2468 18153 2496
rect 18012 2456 18018 2468
rect 18141 2465 18153 2468
rect 18187 2465 18199 2499
rect 18141 2459 18199 2465
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 20073 2499 20131 2505
rect 20073 2496 20085 2499
rect 19484 2468 20085 2496
rect 19484 2456 19490 2468
rect 20073 2465 20085 2468
rect 20119 2465 20131 2499
rect 20990 2496 20996 2508
rect 20951 2468 20996 2496
rect 20073 2459 20131 2465
rect 20990 2456 20996 2468
rect 21048 2456 21054 2508
rect 15212 2428 15240 2456
rect 14200 2400 15240 2428
rect 17865 2431 17923 2437
rect 7975 2332 9904 2360
rect 10229 2363 10287 2369
rect 7975 2329 7987 2332
rect 7929 2323 7987 2329
rect 10229 2329 10241 2363
rect 10275 2360 10287 2363
rect 12176 2360 12204 2391
rect 10275 2332 12204 2360
rect 10275 2329 10287 2332
rect 10229 2323 10287 2329
rect 8849 2295 8907 2301
rect 8849 2292 8861 2295
rect 7208 2264 8861 2292
rect 8849 2261 8861 2264
rect 8895 2261 8907 2295
rect 8849 2255 8907 2261
rect 11238 2252 11244 2304
rect 11296 2292 11302 2304
rect 11517 2295 11575 2301
rect 11517 2292 11529 2295
rect 11296 2264 11529 2292
rect 11296 2252 11302 2264
rect 11517 2261 11529 2264
rect 11563 2261 11575 2295
rect 11517 2255 11575 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12728 2292 12756 2400
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 19242 2428 19248 2440
rect 17911 2400 19248 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13449 2363 13507 2369
rect 13449 2360 13461 2363
rect 13320 2332 13461 2360
rect 13320 2320 13326 2332
rect 13449 2329 13461 2332
rect 13495 2329 13507 2363
rect 13449 2323 13507 2329
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 13817 2363 13875 2369
rect 13817 2360 13829 2363
rect 13780 2332 13829 2360
rect 13780 2320 13786 2332
rect 13817 2329 13829 2332
rect 13863 2329 13875 2363
rect 13817 2323 13875 2329
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14332 2332 14565 2360
rect 14332 2320 14338 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 14734 2320 14740 2372
rect 14792 2360 14798 2372
rect 14921 2363 14979 2369
rect 14921 2360 14933 2363
rect 14792 2332 14933 2360
rect 14792 2320 14798 2332
rect 14921 2329 14933 2332
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 15289 2363 15347 2369
rect 15289 2360 15301 2363
rect 15252 2332 15301 2360
rect 15252 2320 15258 2332
rect 15289 2329 15301 2332
rect 15335 2329 15347 2363
rect 15654 2360 15660 2372
rect 15615 2332 15660 2360
rect 15289 2323 15347 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 16114 2360 16120 2372
rect 16075 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 16632 2332 16677 2360
rect 16632 2320 16638 2332
rect 17034 2320 17040 2372
rect 17092 2360 17098 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 17092 2332 17233 2360
rect 17092 2320 17098 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17954 2360 17960 2372
rect 17915 2332 17960 2360
rect 17221 2323 17279 2329
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 18966 2360 18972 2372
rect 18927 2332 18972 2360
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 19426 2360 19432 2372
rect 19387 2332 19432 2360
rect 19426 2320 19432 2332
rect 19484 2320 19490 2372
rect 19886 2360 19892 2372
rect 19847 2332 19892 2360
rect 19886 2320 19892 2332
rect 19944 2320 19950 2372
rect 20346 2360 20352 2372
rect 20307 2332 20352 2360
rect 20346 2320 20352 2332
rect 20404 2320 20410 2372
rect 20806 2360 20812 2372
rect 20767 2332 20812 2360
rect 20806 2320 20812 2332
rect 20864 2320 20870 2372
rect 21266 2360 21272 2372
rect 21227 2332 21272 2360
rect 21266 2320 21272 2332
rect 21324 2320 21330 2372
rect 11940 2264 12756 2292
rect 12805 2295 12863 2301
rect 11940 2252 11946 2264
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 15930 2292 15936 2304
rect 12851 2264 15936 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 18509 2295 18567 2301
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 18598 2292 18604 2304
rect 18555 2264 18604 2292
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 5718 2088 5724 2100
rect 3200 2060 5724 2088
rect 3200 2048 3206 2060
rect 5718 2048 5724 2060
rect 5776 2048 5782 2100
rect 7098 2048 7104 2100
rect 7156 2088 7162 2100
rect 13354 2088 13360 2100
rect 7156 2060 13360 2088
rect 7156 2048 7162 2060
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 3786 1980 3792 2032
rect 3844 2020 3850 2032
rect 6362 2020 6368 2032
rect 3844 1992 6368 2020
rect 3844 1980 3850 1992
rect 6362 1980 6368 1992
rect 6420 1980 6426 2032
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 12894 2020 12900 2032
rect 11480 1992 12900 2020
rect 11480 1980 11486 1992
rect 12894 1980 12900 1992
rect 12952 1980 12958 2032
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 6638 1952 6644 1964
rect 4120 1924 6644 1952
rect 4120 1912 4126 1924
rect 6638 1912 6644 1924
rect 6696 1912 6702 1964
rect 5166 1844 5172 1896
rect 5224 1884 5230 1896
rect 11238 1884 11244 1896
rect 5224 1856 11244 1884
rect 5224 1844 5230 1856
rect 11238 1844 11244 1856
rect 11296 1844 11302 1896
rect 658 1776 664 1828
rect 716 1816 722 1828
rect 4246 1816 4252 1828
rect 716 1788 4252 1816
rect 716 1776 722 1788
rect 4246 1776 4252 1788
rect 4304 1776 4310 1828
rect 5810 1776 5816 1828
rect 5868 1816 5874 1828
rect 6454 1816 6460 1828
rect 5868 1788 6460 1816
rect 5868 1776 5874 1788
rect 6454 1776 6460 1788
rect 6512 1776 6518 1828
rect 4154 1708 4160 1760
rect 4212 1748 4218 1760
rect 5442 1748 5448 1760
rect 4212 1720 5448 1748
rect 4212 1708 4218 1720
rect 5442 1708 5448 1720
rect 5500 1708 5506 1760
rect 4338 1640 4344 1692
rect 4396 1680 4402 1692
rect 8938 1680 8944 1692
rect 4396 1652 8944 1680
rect 4396 1640 4402 1652
rect 8938 1640 8944 1652
rect 8996 1640 9002 1692
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2780 20544 2832 20596
rect 3884 20544 3936 20596
rect 4068 20544 4120 20596
rect 2872 20519 2924 20528
rect 2872 20485 2881 20519
rect 2881 20485 2915 20519
rect 2915 20485 2924 20519
rect 2872 20476 2924 20485
rect 3240 20519 3292 20528
rect 3240 20485 3249 20519
rect 3249 20485 3283 20519
rect 3283 20485 3292 20519
rect 3240 20476 3292 20485
rect 3516 20476 3568 20528
rect 5172 20544 5224 20596
rect 4344 20476 4396 20528
rect 1124 20408 1176 20460
rect 3700 20408 3752 20460
rect 5816 20408 5868 20460
rect 6092 20408 6144 20460
rect 7196 20544 7248 20596
rect 6460 20476 6512 20528
rect 7472 20451 7524 20460
rect 204 20340 256 20392
rect 1584 20340 1636 20392
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 4344 20340 4396 20392
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 5724 20340 5776 20392
rect 6276 20340 6328 20392
rect 6920 20340 6972 20392
rect 7472 20417 7481 20451
rect 7481 20417 7515 20451
rect 7515 20417 7524 20451
rect 7472 20408 7524 20417
rect 10140 20544 10192 20596
rect 10600 20544 10652 20596
rect 21364 20544 21416 20596
rect 7656 20340 7708 20392
rect 8392 20340 8444 20392
rect 8484 20340 8536 20392
rect 8944 20340 8996 20392
rect 11796 20476 11848 20528
rect 13084 20519 13136 20528
rect 13084 20485 13093 20519
rect 13093 20485 13127 20519
rect 13127 20485 13136 20519
rect 13084 20476 13136 20485
rect 13544 20519 13596 20528
rect 13544 20485 13553 20519
rect 13553 20485 13587 20519
rect 13587 20485 13596 20519
rect 13544 20476 13596 20485
rect 14004 20519 14056 20528
rect 14004 20485 14013 20519
rect 14013 20485 14047 20519
rect 14047 20485 14056 20519
rect 14004 20476 14056 20485
rect 14464 20476 14516 20528
rect 14924 20519 14976 20528
rect 14924 20485 14933 20519
rect 14933 20485 14967 20519
rect 14967 20485 14976 20519
rect 14924 20476 14976 20485
rect 15384 20519 15436 20528
rect 15384 20485 15393 20519
rect 15393 20485 15427 20519
rect 15427 20485 15436 20519
rect 15384 20476 15436 20485
rect 15844 20519 15896 20528
rect 15844 20485 15853 20519
rect 15853 20485 15887 20519
rect 15887 20485 15896 20519
rect 15844 20476 15896 20485
rect 16304 20519 16356 20528
rect 16304 20485 16313 20519
rect 16313 20485 16347 20519
rect 16347 20485 16356 20519
rect 16304 20476 16356 20485
rect 16764 20519 16816 20528
rect 16764 20485 16773 20519
rect 16773 20485 16807 20519
rect 16807 20485 16816 20519
rect 16764 20476 16816 20485
rect 17684 20519 17736 20528
rect 17684 20485 17693 20519
rect 17693 20485 17727 20519
rect 17727 20485 17736 20519
rect 17684 20476 17736 20485
rect 18144 20519 18196 20528
rect 18144 20485 18153 20519
rect 18153 20485 18187 20519
rect 18187 20485 18196 20519
rect 18144 20476 18196 20485
rect 18604 20519 18656 20528
rect 18604 20485 18613 20519
rect 18613 20485 18647 20519
rect 18647 20485 18656 20519
rect 18604 20476 18656 20485
rect 19064 20519 19116 20528
rect 19064 20485 19073 20519
rect 19073 20485 19107 20519
rect 19107 20485 19116 20519
rect 19064 20476 19116 20485
rect 19524 20476 19576 20528
rect 19984 20476 20036 20528
rect 20444 20476 20496 20528
rect 20904 20476 20956 20528
rect 9128 20408 9180 20460
rect 11060 20408 11112 20460
rect 9404 20340 9456 20392
rect 10232 20383 10284 20392
rect 10232 20349 10241 20383
rect 10241 20349 10275 20383
rect 10275 20349 10284 20383
rect 10232 20340 10284 20349
rect 10324 20340 10376 20392
rect 11244 20340 11296 20392
rect 1676 20315 1728 20324
rect 1676 20281 1685 20315
rect 1685 20281 1719 20315
rect 1719 20281 1728 20315
rect 1676 20272 1728 20281
rect 1952 20315 2004 20324
rect 1952 20281 1961 20315
rect 1961 20281 1995 20315
rect 1995 20281 2004 20315
rect 1952 20272 2004 20281
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 2688 20315 2740 20324
rect 2688 20281 2697 20315
rect 2697 20281 2731 20315
rect 2731 20281 2740 20315
rect 2688 20272 2740 20281
rect 2964 20272 3016 20324
rect 3332 20272 3384 20324
rect 5356 20272 5408 20324
rect 7748 20315 7800 20324
rect 1860 20247 1912 20256
rect 1860 20213 1869 20247
rect 1869 20213 1903 20247
rect 1903 20213 1912 20247
rect 1860 20204 1912 20213
rect 2780 20204 2832 20256
rect 3516 20204 3568 20256
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 4160 20204 4212 20256
rect 5908 20204 5960 20256
rect 6276 20204 6328 20256
rect 6920 20247 6972 20256
rect 6920 20213 6929 20247
rect 6929 20213 6963 20247
rect 6963 20213 6972 20247
rect 6920 20204 6972 20213
rect 7288 20247 7340 20256
rect 7288 20213 7297 20247
rect 7297 20213 7331 20247
rect 7331 20213 7340 20247
rect 7288 20204 7340 20213
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7748 20281 7757 20315
rect 7757 20281 7791 20315
rect 7791 20281 7800 20315
rect 7748 20272 7800 20281
rect 7380 20204 7432 20213
rect 7656 20204 7708 20256
rect 9312 20272 9364 20324
rect 9864 20272 9916 20324
rect 10600 20315 10652 20324
rect 10600 20281 10609 20315
rect 10609 20281 10643 20315
rect 10643 20281 10652 20315
rect 10600 20272 10652 20281
rect 11060 20315 11112 20324
rect 11060 20281 11069 20315
rect 11069 20281 11103 20315
rect 11103 20281 11112 20315
rect 11060 20272 11112 20281
rect 11704 20272 11756 20324
rect 12072 20315 12124 20324
rect 12072 20281 12081 20315
rect 12081 20281 12115 20315
rect 12115 20281 12124 20315
rect 12072 20272 12124 20281
rect 12348 20340 12400 20392
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 21824 20408 21876 20460
rect 12440 20340 12492 20349
rect 13636 20340 13688 20392
rect 15384 20340 15436 20392
rect 17960 20340 18012 20392
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 22744 20340 22796 20392
rect 12900 20272 12952 20324
rect 13268 20315 13320 20324
rect 13268 20281 13277 20315
rect 13277 20281 13311 20315
rect 13311 20281 13320 20315
rect 13268 20272 13320 20281
rect 13728 20315 13780 20324
rect 13728 20281 13737 20315
rect 13737 20281 13771 20315
rect 13771 20281 13780 20315
rect 13728 20272 13780 20281
rect 14372 20272 14424 20324
rect 15200 20272 15252 20324
rect 15660 20272 15712 20324
rect 16212 20272 16264 20324
rect 16672 20272 16724 20324
rect 17868 20315 17920 20324
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 9220 20247 9272 20256
rect 9220 20213 9229 20247
rect 9229 20213 9263 20247
rect 9263 20213 9272 20247
rect 9220 20204 9272 20213
rect 9404 20204 9456 20256
rect 9772 20204 9824 20256
rect 10416 20204 10468 20256
rect 11244 20204 11296 20256
rect 11888 20204 11940 20256
rect 12164 20204 12216 20256
rect 12440 20204 12492 20256
rect 13544 20204 13596 20256
rect 13820 20204 13872 20256
rect 17868 20281 17877 20315
rect 17877 20281 17911 20315
rect 17911 20281 17920 20315
rect 17868 20272 17920 20281
rect 18144 20272 18196 20324
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 18880 20272 18932 20324
rect 19524 20315 19576 20324
rect 19524 20281 19533 20315
rect 19533 20281 19567 20315
rect 19567 20281 19576 20315
rect 19524 20272 19576 20281
rect 20076 20315 20128 20324
rect 20076 20281 20085 20315
rect 20085 20281 20119 20315
rect 20119 20281 20128 20315
rect 20076 20272 20128 20281
rect 20444 20315 20496 20324
rect 20444 20281 20453 20315
rect 20453 20281 20487 20315
rect 20487 20281 20496 20315
rect 20444 20272 20496 20281
rect 20536 20272 20588 20324
rect 21364 20247 21416 20256
rect 21364 20213 21373 20247
rect 21373 20213 21407 20247
rect 21407 20213 21416 20247
rect 21364 20204 21416 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1768 20000 1820 20052
rect 2688 20000 2740 20052
rect 6460 20000 6512 20052
rect 2044 19864 2096 19916
rect 664 19796 716 19848
rect 2412 19907 2464 19916
rect 2412 19873 2421 19907
rect 2421 19873 2455 19907
rect 2455 19873 2464 19907
rect 2872 19907 2924 19916
rect 2412 19864 2464 19873
rect 2872 19873 2881 19907
rect 2881 19873 2915 19907
rect 2915 19873 2924 19907
rect 2872 19864 2924 19873
rect 5172 19932 5224 19984
rect 8484 20000 8536 20052
rect 8944 20000 8996 20052
rect 11796 20000 11848 20052
rect 12624 20000 12676 20052
rect 12900 20000 12952 20052
rect 13544 20000 13596 20052
rect 17868 20000 17920 20052
rect 21548 20043 21600 20052
rect 21548 20009 21557 20043
rect 21557 20009 21591 20043
rect 21591 20009 21600 20043
rect 21548 20000 21600 20009
rect 3148 19864 3200 19916
rect 3424 19864 3476 19916
rect 3700 19864 3752 19916
rect 4896 19864 4948 19916
rect 5264 19864 5316 19916
rect 3516 19839 3568 19848
rect 1400 19771 1452 19780
rect 1400 19737 1409 19771
rect 1409 19737 1443 19771
rect 1443 19737 1452 19771
rect 1400 19728 1452 19737
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 8300 19932 8352 19984
rect 11060 19932 11112 19984
rect 6552 19864 6604 19916
rect 7104 19864 7156 19916
rect 7472 19864 7524 19916
rect 9128 19864 9180 19916
rect 12072 19907 12124 19916
rect 12072 19873 12081 19907
rect 12081 19873 12115 19907
rect 12115 19873 12124 19907
rect 12072 19864 12124 19873
rect 12624 19864 12676 19916
rect 17224 19975 17276 19984
rect 17224 19941 17233 19975
rect 17233 19941 17267 19975
rect 17267 19941 17276 19975
rect 17224 19932 17276 19941
rect 6460 19839 6512 19848
rect 3056 19728 3108 19780
rect 4252 19728 4304 19780
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 10508 19839 10560 19848
rect 5356 19728 5408 19780
rect 4804 19703 4856 19712
rect 4804 19669 4813 19703
rect 4813 19669 4847 19703
rect 4847 19669 4856 19703
rect 4804 19660 4856 19669
rect 5816 19660 5868 19712
rect 7012 19728 7064 19780
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 12348 19796 12400 19848
rect 12808 19796 12860 19848
rect 16580 19864 16632 19916
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 8760 19728 8812 19780
rect 11796 19728 11848 19780
rect 8484 19660 8536 19712
rect 8668 19660 8720 19712
rect 11980 19703 12032 19712
rect 11980 19669 11989 19703
rect 11989 19669 12023 19703
rect 12023 19669 12032 19703
rect 11980 19660 12032 19669
rect 12532 19660 12584 19712
rect 12992 19660 13044 19712
rect 13820 19660 13872 19712
rect 14280 19660 14332 19712
rect 16580 19703 16632 19712
rect 16580 19669 16589 19703
rect 16589 19669 16623 19703
rect 16623 19669 16632 19703
rect 16580 19660 16632 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19456 2004 19508
rect 2320 19456 2372 19508
rect 2872 19456 2924 19508
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 5356 19456 5408 19508
rect 7472 19456 7524 19508
rect 9128 19499 9180 19508
rect 9128 19465 9137 19499
rect 9137 19465 9171 19499
rect 9171 19465 9180 19499
rect 9128 19456 9180 19465
rect 10232 19456 10284 19508
rect 13268 19456 13320 19508
rect 13728 19456 13780 19508
rect 14372 19456 14424 19508
rect 15660 19456 15712 19508
rect 16212 19456 16264 19508
rect 17408 19456 17460 19508
rect 18144 19456 18196 19508
rect 18788 19456 18840 19508
rect 20536 19456 20588 19508
rect 9496 19388 9548 19440
rect 15384 19388 15436 19440
rect 20444 19388 20496 19440
rect 1400 19227 1452 19236
rect 1400 19193 1409 19227
rect 1409 19193 1443 19227
rect 1443 19193 1452 19227
rect 1400 19184 1452 19193
rect 1584 19227 1636 19236
rect 1584 19193 1593 19227
rect 1593 19193 1627 19227
rect 1627 19193 1636 19227
rect 1584 19184 1636 19193
rect 3516 19252 3568 19304
rect 4252 19295 4304 19304
rect 4252 19261 4270 19295
rect 4270 19261 4304 19295
rect 4252 19252 4304 19261
rect 3056 19116 3108 19168
rect 3792 19184 3844 19236
rect 5908 19320 5960 19372
rect 7288 19320 7340 19372
rect 8484 19363 8536 19372
rect 8484 19329 8493 19363
rect 8493 19329 8527 19363
rect 8527 19329 8536 19363
rect 8484 19320 8536 19329
rect 6920 19252 6972 19304
rect 6460 19116 6512 19168
rect 8668 19320 8720 19372
rect 9404 19320 9456 19372
rect 9220 19252 9272 19304
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 12992 19320 13044 19372
rect 11980 19295 12032 19304
rect 11980 19261 12014 19295
rect 12014 19261 12032 19295
rect 11980 19252 12032 19261
rect 12532 19252 12584 19304
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 13820 19252 13872 19304
rect 9956 19184 10008 19236
rect 14280 19252 14332 19304
rect 14556 19252 14608 19304
rect 15292 19252 15344 19304
rect 15568 19252 15620 19304
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 16120 19252 16172 19304
rect 16396 19252 16448 19304
rect 20076 19320 20128 19372
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 11704 19116 11756 19168
rect 17132 19227 17184 19236
rect 17132 19193 17141 19227
rect 17141 19193 17175 19227
rect 17175 19193 17184 19227
rect 17132 19184 17184 19193
rect 18144 19252 18196 19304
rect 18328 19295 18380 19304
rect 18328 19261 18337 19295
rect 18337 19261 18371 19295
rect 18371 19261 18380 19295
rect 18328 19252 18380 19261
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 22284 19184 22336 19236
rect 15200 19116 15252 19168
rect 16672 19116 16724 19168
rect 17960 19116 18012 19168
rect 18788 19159 18840 19168
rect 18788 19125 18797 19159
rect 18797 19125 18831 19159
rect 18831 19125 18840 19159
rect 18788 19116 18840 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1584 18912 1636 18964
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 2412 18912 2464 18964
rect 3240 18912 3292 18964
rect 3516 18912 3568 18964
rect 3608 18912 3660 18964
rect 4252 18887 4304 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 1768 18776 1820 18828
rect 2044 18776 2096 18828
rect 4252 18853 4261 18887
rect 4261 18853 4295 18887
rect 4295 18853 4304 18887
rect 4252 18844 4304 18853
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 2412 18708 2464 18760
rect 3240 18776 3292 18828
rect 3516 18776 3568 18828
rect 5540 18912 5592 18964
rect 7012 18955 7064 18964
rect 7012 18921 7021 18955
rect 7021 18921 7055 18955
rect 7055 18921 7064 18955
rect 7012 18912 7064 18921
rect 7380 18955 7432 18964
rect 7380 18921 7389 18955
rect 7389 18921 7423 18955
rect 7423 18921 7432 18955
rect 7380 18912 7432 18921
rect 7656 18912 7708 18964
rect 8392 18955 8444 18964
rect 8392 18921 8401 18955
rect 8401 18921 8435 18955
rect 8435 18921 8444 18955
rect 8392 18912 8444 18921
rect 9312 18955 9364 18964
rect 9312 18921 9321 18955
rect 9321 18921 9355 18955
rect 9355 18921 9364 18955
rect 9312 18912 9364 18921
rect 10324 18912 10376 18964
rect 10692 18912 10744 18964
rect 11152 18912 11204 18964
rect 11704 18955 11756 18964
rect 11704 18921 11713 18955
rect 11713 18921 11747 18955
rect 11747 18921 11756 18955
rect 11704 18912 11756 18921
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 12256 18912 12308 18964
rect 13728 18912 13780 18964
rect 14556 18912 14608 18964
rect 15936 18912 15988 18964
rect 18328 18912 18380 18964
rect 19616 18912 19668 18964
rect 5816 18844 5868 18896
rect 6460 18844 6512 18896
rect 8300 18844 8352 18896
rect 11796 18844 11848 18896
rect 15568 18887 15620 18896
rect 4988 18776 5040 18828
rect 6368 18776 6420 18828
rect 7288 18776 7340 18828
rect 8944 18776 8996 18828
rect 9220 18819 9272 18828
rect 9220 18785 9229 18819
rect 9229 18785 9263 18819
rect 9263 18785 9272 18819
rect 9220 18776 9272 18785
rect 10784 18776 10836 18828
rect 11152 18819 11204 18828
rect 11152 18785 11161 18819
rect 11161 18785 11195 18819
rect 11195 18785 11204 18819
rect 11152 18776 11204 18785
rect 12716 18776 12768 18828
rect 14004 18819 14056 18828
rect 14004 18785 14013 18819
rect 14013 18785 14047 18819
rect 14047 18785 14056 18819
rect 14004 18776 14056 18785
rect 14464 18819 14516 18828
rect 14464 18785 14473 18819
rect 14473 18785 14507 18819
rect 14507 18785 14516 18819
rect 14464 18776 14516 18785
rect 2964 18640 3016 18692
rect 3516 18640 3568 18692
rect 4344 18751 4396 18760
rect 4344 18717 4353 18751
rect 4353 18717 4387 18751
rect 4387 18717 4396 18751
rect 4344 18708 4396 18717
rect 3976 18640 4028 18692
rect 2596 18572 2648 18624
rect 3240 18572 3292 18624
rect 5172 18708 5224 18760
rect 6552 18708 6604 18760
rect 8668 18708 8720 18760
rect 9956 18751 10008 18760
rect 9956 18717 9965 18751
rect 9965 18717 9999 18751
rect 9999 18717 10008 18751
rect 9956 18708 10008 18717
rect 5356 18640 5408 18692
rect 6644 18640 6696 18692
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 6552 18572 6604 18624
rect 10692 18708 10744 18760
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 16672 18819 16724 18828
rect 16672 18785 16681 18819
rect 16681 18785 16715 18819
rect 16715 18785 16724 18819
rect 16672 18776 16724 18785
rect 18696 18819 18748 18828
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 17316 18708 17368 18760
rect 19524 18640 19576 18692
rect 11060 18572 11112 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 18144 18572 18196 18624
rect 18604 18572 18656 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 1952 18368 2004 18420
rect 2964 18368 3016 18420
rect 3240 18368 3292 18420
rect 3976 18411 4028 18420
rect 2504 18343 2556 18352
rect 2504 18309 2513 18343
rect 2513 18309 2547 18343
rect 2547 18309 2556 18343
rect 2504 18300 2556 18309
rect 3976 18377 3985 18411
rect 3985 18377 4019 18411
rect 4019 18377 4028 18411
rect 3976 18368 4028 18377
rect 4344 18411 4396 18420
rect 4344 18377 4353 18411
rect 4353 18377 4387 18411
rect 4387 18377 4396 18411
rect 4344 18368 4396 18377
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 6184 18368 6236 18420
rect 7104 18368 7156 18420
rect 7564 18368 7616 18420
rect 9220 18368 9272 18420
rect 10324 18368 10376 18420
rect 12072 18368 12124 18420
rect 5448 18300 5500 18352
rect 9680 18300 9732 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 1492 18232 1544 18284
rect 4252 18275 4304 18284
rect 1584 18139 1636 18148
rect 1584 18105 1593 18139
rect 1593 18105 1627 18139
rect 1627 18105 1636 18139
rect 1584 18096 1636 18105
rect 2136 18164 2188 18216
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2504 18096 2556 18148
rect 2228 18071 2280 18080
rect 2228 18037 2237 18071
rect 2237 18037 2271 18071
rect 2271 18037 2280 18071
rect 2228 18028 2280 18037
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 5080 18232 5132 18284
rect 5264 18232 5316 18284
rect 9128 18232 9180 18284
rect 9312 18232 9364 18284
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 12072 18232 12124 18284
rect 6000 18207 6052 18216
rect 6000 18173 6009 18207
rect 6009 18173 6043 18207
rect 6043 18173 6052 18207
rect 6000 18164 6052 18173
rect 3516 18096 3568 18148
rect 2872 18028 2924 18080
rect 2964 18028 3016 18080
rect 8576 18096 8628 18148
rect 10692 18164 10744 18216
rect 16672 18164 16724 18216
rect 13912 18096 13964 18148
rect 14832 18096 14884 18148
rect 3700 18028 3752 18080
rect 4620 18028 4672 18080
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 4896 18028 4948 18080
rect 5172 18028 5224 18080
rect 6460 18028 6512 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 11060 18028 11112 18080
rect 11796 18028 11848 18080
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1492 17867 1544 17876
rect 1492 17833 1501 17867
rect 1501 17833 1535 17867
rect 1535 17833 1544 17867
rect 1492 17824 1544 17833
rect 1584 17824 1636 17876
rect 2504 17824 2556 17876
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 3516 17867 3568 17876
rect 3516 17833 3525 17867
rect 3525 17833 3559 17867
rect 3559 17833 3568 17867
rect 3516 17824 3568 17833
rect 4160 17824 4212 17876
rect 4620 17824 4672 17876
rect 4896 17824 4948 17876
rect 8852 17824 8904 17876
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 7656 17756 7708 17808
rect 3332 17688 3384 17740
rect 3424 17731 3476 17740
rect 3424 17697 3433 17731
rect 3433 17697 3467 17731
rect 3467 17697 3476 17731
rect 3424 17688 3476 17697
rect 4252 17688 4304 17740
rect 2136 17552 2188 17604
rect 4804 17620 4856 17672
rect 5356 17620 5408 17672
rect 6552 17620 6604 17672
rect 2964 17552 3016 17604
rect 4344 17552 4396 17604
rect 3240 17484 3292 17536
rect 4252 17484 4304 17536
rect 5448 17484 5500 17536
rect 7380 17688 7432 17740
rect 7472 17620 7524 17672
rect 8668 17663 8720 17672
rect 7012 17552 7064 17604
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9864 17824 9916 17876
rect 12348 17824 12400 17876
rect 13636 17824 13688 17876
rect 9864 17688 9916 17740
rect 10968 17756 11020 17808
rect 15476 17756 15528 17808
rect 16396 17756 16448 17808
rect 10508 17688 10560 17740
rect 12072 17731 12124 17740
rect 12072 17697 12106 17731
rect 12106 17697 12124 17731
rect 12072 17688 12124 17697
rect 13360 17688 13412 17740
rect 11704 17620 11756 17672
rect 11060 17484 11112 17536
rect 11980 17484 12032 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1860 17323 1912 17332
rect 1860 17289 1869 17323
rect 1869 17289 1903 17323
rect 1903 17289 1912 17323
rect 1860 17280 1912 17289
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 2044 17212 2096 17264
rect 4344 17280 4396 17332
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 7472 17280 7524 17332
rect 1676 17144 1728 17196
rect 2228 17076 2280 17128
rect 2964 17144 3016 17196
rect 9864 17280 9916 17332
rect 10968 17323 11020 17332
rect 10968 17289 10977 17323
rect 10977 17289 11011 17323
rect 11011 17289 11020 17323
rect 10968 17280 11020 17289
rect 12072 17280 12124 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 9312 17255 9364 17264
rect 9312 17221 9321 17255
rect 9321 17221 9355 17255
rect 9355 17221 9364 17255
rect 9312 17212 9364 17221
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 1952 17051 2004 17060
rect 1952 17017 1961 17051
rect 1961 17017 1995 17051
rect 1995 17017 2004 17051
rect 1952 17008 2004 17017
rect 3056 17076 3108 17128
rect 3976 17076 4028 17128
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 10508 17119 10560 17128
rect 3792 17008 3844 17060
rect 6368 17008 6420 17060
rect 10508 17085 10526 17119
rect 10526 17085 10560 17119
rect 10508 17076 10560 17085
rect 11060 17076 11112 17128
rect 11152 17076 11204 17128
rect 11980 17119 12032 17128
rect 11980 17085 12014 17119
rect 12014 17085 12032 17119
rect 11980 17076 12032 17085
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 7104 17008 7156 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 3424 16940 3476 16992
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 12072 16940 12124 16992
rect 18144 16940 18196 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2228 16779 2280 16788
rect 2228 16745 2237 16779
rect 2237 16745 2271 16779
rect 2271 16745 2280 16779
rect 2228 16736 2280 16745
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 2964 16736 3016 16788
rect 5448 16736 5500 16788
rect 7380 16779 7432 16788
rect 2412 16668 2464 16720
rect 3424 16711 3476 16720
rect 1676 16600 1728 16652
rect 1860 16600 1912 16652
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 3424 16677 3433 16711
rect 3433 16677 3467 16711
rect 3467 16677 3476 16711
rect 3424 16668 3476 16677
rect 6828 16668 6880 16720
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 2964 16600 3016 16652
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 5264 16600 5316 16652
rect 3792 16464 3844 16516
rect 6460 16532 6512 16584
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 7104 16464 7156 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 3424 16396 3476 16448
rect 8668 16736 8720 16788
rect 10968 16736 11020 16788
rect 11336 16736 11388 16788
rect 11796 16736 11848 16788
rect 12164 16736 12216 16788
rect 11704 16668 11756 16720
rect 13452 16736 13504 16788
rect 14464 16736 14516 16788
rect 10784 16600 10836 16652
rect 10508 16532 10560 16584
rect 11980 16600 12032 16652
rect 11888 16532 11940 16584
rect 14556 16600 14608 16652
rect 10876 16396 10928 16448
rect 11704 16396 11756 16448
rect 13084 16396 13136 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1584 16192 1636 16244
rect 1860 16192 1912 16244
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 6368 16192 6420 16244
rect 6828 16192 6880 16244
rect 8484 16099 8536 16108
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 3424 15988 3476 16040
rect 3792 15988 3844 16040
rect 4160 16031 4212 16040
rect 4160 15997 4194 16031
rect 4194 15997 4212 16031
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 4160 15988 4212 15997
rect 7012 15988 7064 16040
rect 9864 16192 9916 16244
rect 10416 16192 10468 16244
rect 10784 16192 10836 16244
rect 11244 16192 11296 16244
rect 13176 16192 13228 16244
rect 11704 16124 11756 16176
rect 13820 16124 13872 16176
rect 11428 16056 11480 16108
rect 12532 16056 12584 16108
rect 14096 16056 14148 16108
rect 1400 15963 1452 15972
rect 1400 15929 1409 15963
rect 1409 15929 1443 15963
rect 1443 15929 1452 15963
rect 1400 15920 1452 15929
rect 1584 15963 1636 15972
rect 1584 15929 1593 15963
rect 1593 15929 1627 15963
rect 1627 15929 1636 15963
rect 1584 15920 1636 15929
rect 11704 15988 11756 16040
rect 12440 15988 12492 16040
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 5724 15852 5776 15904
rect 6460 15895 6512 15904
rect 6460 15861 6469 15895
rect 6469 15861 6503 15895
rect 6503 15861 6512 15895
rect 6460 15852 6512 15861
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11244 15852 11296 15904
rect 14188 15920 14240 15972
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1584 15648 1636 15700
rect 1952 15648 2004 15700
rect 4344 15648 4396 15700
rect 4804 15648 4856 15700
rect 5540 15648 5592 15700
rect 8484 15648 8536 15700
rect 9036 15648 9088 15700
rect 3608 15580 3660 15632
rect 5172 15623 5224 15632
rect 5172 15589 5181 15623
rect 5181 15589 5215 15623
rect 5215 15589 5224 15623
rect 5172 15580 5224 15589
rect 6920 15580 6972 15632
rect 9496 15648 9548 15700
rect 9956 15648 10008 15700
rect 10140 15648 10192 15700
rect 10416 15648 10468 15700
rect 13544 15648 13596 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 11428 15580 11480 15632
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 2228 15555 2280 15564
rect 2228 15521 2237 15555
rect 2237 15521 2271 15555
rect 2271 15521 2280 15555
rect 2228 15512 2280 15521
rect 2044 15444 2096 15496
rect 1400 15419 1452 15428
rect 1400 15385 1409 15419
rect 1409 15385 1443 15419
rect 1443 15385 1452 15419
rect 1400 15376 1452 15385
rect 4160 15512 4212 15564
rect 6368 15512 6420 15564
rect 11060 15512 11112 15564
rect 11796 15512 11848 15564
rect 12532 15512 12584 15564
rect 10968 15444 11020 15496
rect 5540 15376 5592 15428
rect 1676 15308 1728 15360
rect 6184 15308 6236 15360
rect 7380 15308 7432 15360
rect 8208 15351 8260 15360
rect 8208 15317 8217 15351
rect 8217 15317 8251 15351
rect 8251 15317 8260 15351
rect 8208 15308 8260 15317
rect 11060 15308 11112 15360
rect 11980 15308 12032 15360
rect 12992 15555 13044 15564
rect 12992 15521 13026 15555
rect 13026 15521 13044 15555
rect 12992 15512 13044 15521
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 12992 15308 13044 15360
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1952 15104 2004 15156
rect 2228 15104 2280 15156
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 6828 15104 6880 15156
rect 3700 15036 3752 15088
rect 7564 15104 7616 15156
rect 10600 15104 10652 15156
rect 11244 15147 11296 15156
rect 11244 15113 11253 15147
rect 11253 15113 11287 15147
rect 11287 15113 11296 15147
rect 11244 15104 11296 15113
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 12440 15104 12492 15113
rect 13084 15104 13136 15156
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 6828 14968 6880 15020
rect 1768 14832 1820 14884
rect 3792 14900 3844 14952
rect 6368 14900 6420 14952
rect 2780 14832 2832 14884
rect 3056 14832 3108 14884
rect 3792 14764 3844 14816
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 7472 14832 7524 14884
rect 12256 15036 12308 15088
rect 8208 14900 8260 14952
rect 9128 14900 9180 14952
rect 9680 14900 9732 14952
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 13176 15036 13228 15088
rect 19064 15036 19116 15088
rect 12992 14968 13044 15020
rect 15200 14968 15252 15020
rect 15752 14968 15804 15020
rect 9588 14832 9640 14884
rect 8300 14807 8352 14816
rect 8300 14773 8309 14807
rect 8309 14773 8343 14807
rect 8343 14773 8352 14807
rect 8300 14764 8352 14773
rect 11060 14900 11112 14952
rect 13544 14900 13596 14952
rect 10968 14832 11020 14884
rect 12808 14875 12860 14884
rect 12808 14841 12817 14875
rect 12817 14841 12851 14875
rect 12851 14841 12860 14875
rect 12808 14832 12860 14841
rect 11796 14764 11848 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 14740 14764 14792 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2044 14603 2096 14612
rect 2044 14569 2053 14603
rect 2053 14569 2087 14603
rect 2087 14569 2096 14603
rect 2044 14560 2096 14569
rect 3148 14560 3200 14612
rect 3700 14560 3752 14612
rect 6000 14560 6052 14612
rect 9772 14560 9824 14612
rect 10508 14560 10560 14612
rect 10692 14560 10744 14612
rect 11060 14560 11112 14612
rect 11152 14560 11204 14612
rect 12808 14560 12860 14612
rect 13268 14560 13320 14612
rect 15292 14560 15344 14612
rect 4068 14492 4120 14544
rect 8300 14492 8352 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 3700 14424 3752 14476
rect 2320 14356 2372 14408
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 2872 14220 2924 14272
rect 3516 14220 3568 14272
rect 4252 14220 4304 14272
rect 7564 14424 7616 14476
rect 10140 14492 10192 14544
rect 7472 14356 7524 14408
rect 9680 14424 9732 14476
rect 10048 14424 10100 14476
rect 10232 14424 10284 14476
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 15200 14492 15252 14544
rect 9220 14356 9272 14408
rect 10692 14356 10744 14408
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 14096 14424 14148 14476
rect 11060 14356 11112 14365
rect 12256 14356 12308 14408
rect 13084 14356 13136 14408
rect 13360 14356 13412 14408
rect 13820 14356 13872 14408
rect 14372 14356 14424 14408
rect 9496 14331 9548 14340
rect 9496 14297 9505 14331
rect 9505 14297 9539 14331
rect 9539 14297 9548 14331
rect 9496 14288 9548 14297
rect 12072 14288 12124 14340
rect 13728 14288 13780 14340
rect 5540 14220 5592 14272
rect 7288 14220 7340 14272
rect 9772 14220 9824 14272
rect 11888 14220 11940 14272
rect 12348 14220 12400 14272
rect 13268 14220 13320 14272
rect 15660 14220 15712 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1492 14059 1544 14068
rect 1492 14025 1501 14059
rect 1501 14025 1535 14059
rect 1535 14025 1544 14059
rect 1492 14016 1544 14025
rect 1952 14016 2004 14068
rect 2780 14016 2832 14068
rect 2320 13991 2372 14000
rect 2320 13957 2329 13991
rect 2329 13957 2363 13991
rect 2363 13957 2372 13991
rect 2320 13948 2372 13957
rect 10968 14016 11020 14068
rect 12440 14016 12492 14068
rect 12624 14059 12676 14068
rect 12624 14025 12633 14059
rect 12633 14025 12667 14059
rect 12667 14025 12676 14059
rect 12624 14016 12676 14025
rect 12900 14016 12952 14068
rect 7472 13948 7524 14000
rect 4068 13880 4120 13932
rect 4252 13880 4304 13932
rect 7656 13880 7708 13932
rect 9680 13948 9732 14000
rect 9312 13880 9364 13932
rect 10232 13880 10284 13932
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2044 13812 2096 13864
rect 2412 13812 2464 13864
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 3516 13855 3568 13864
rect 2872 13812 2924 13821
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 3700 13812 3752 13864
rect 6000 13812 6052 13864
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 6368 13744 6420 13796
rect 8392 13812 8444 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 5080 13719 5132 13728
rect 5080 13685 5089 13719
rect 5089 13685 5123 13719
rect 5123 13685 5132 13719
rect 5080 13676 5132 13685
rect 5172 13676 5224 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 10324 13812 10376 13864
rect 8576 13744 8628 13796
rect 9220 13744 9272 13796
rect 11152 13880 11204 13932
rect 12808 13880 12860 13932
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 11704 13812 11756 13864
rect 14740 13880 14792 13932
rect 15660 13880 15712 13932
rect 14096 13812 14148 13864
rect 21364 13812 21416 13864
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 9588 13676 9640 13728
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 12532 13676 12584 13728
rect 12624 13676 12676 13728
rect 13268 13676 13320 13728
rect 13544 13676 13596 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 14648 13719 14700 13728
rect 14648 13685 14657 13719
rect 14657 13685 14691 13719
rect 14691 13685 14700 13719
rect 14648 13676 14700 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 1492 13515 1544 13524
rect 1492 13481 1501 13515
rect 1501 13481 1535 13515
rect 1535 13481 1544 13515
rect 1492 13472 1544 13481
rect 4252 13472 4304 13524
rect 6000 13515 6052 13524
rect 6000 13481 6009 13515
rect 6009 13481 6043 13515
rect 6043 13481 6052 13515
rect 6000 13472 6052 13481
rect 8668 13515 8720 13524
rect 1768 13404 1820 13456
rect 5540 13404 5592 13456
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 5632 13379 5684 13388
rect 6460 13404 6512 13456
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9036 13472 9088 13524
rect 13176 13472 13228 13524
rect 13636 13472 13688 13524
rect 14648 13472 14700 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 16304 13472 16356 13524
rect 6920 13404 6972 13456
rect 5632 13345 5650 13379
rect 5650 13345 5684 13379
rect 5632 13336 5684 13345
rect 6828 13336 6880 13388
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 9312 13404 9364 13456
rect 9496 13447 9548 13456
rect 9496 13413 9505 13447
rect 9505 13413 9539 13447
rect 9539 13413 9548 13447
rect 9496 13404 9548 13413
rect 10232 13404 10284 13456
rect 7840 13336 7892 13388
rect 9220 13336 9272 13388
rect 9404 13336 9456 13388
rect 9956 13379 10008 13388
rect 9956 13345 9965 13379
rect 9965 13345 9999 13379
rect 9999 13345 10008 13379
rect 9956 13336 10008 13345
rect 11796 13404 11848 13456
rect 15476 13404 15528 13456
rect 16212 13404 16264 13456
rect 12072 13336 12124 13388
rect 14096 13336 14148 13388
rect 15844 13336 15896 13388
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 2688 13200 2740 13252
rect 6000 13200 6052 13252
rect 6368 13200 6420 13252
rect 1400 13132 1452 13184
rect 1860 13132 1912 13184
rect 5632 13132 5684 13184
rect 7472 13268 7524 13320
rect 6828 13200 6880 13252
rect 8484 13268 8536 13320
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 10140 13243 10192 13252
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 10140 13209 10149 13243
rect 10149 13209 10183 13243
rect 10183 13209 10192 13243
rect 10140 13200 10192 13209
rect 10232 13243 10284 13252
rect 10232 13209 10241 13243
rect 10241 13209 10275 13243
rect 10275 13209 10284 13243
rect 12808 13243 12860 13252
rect 10232 13200 10284 13209
rect 12808 13209 12817 13243
rect 12817 13209 12851 13243
rect 12851 13209 12860 13243
rect 12808 13200 12860 13209
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9312 13132 9364 13184
rect 17960 13200 18012 13252
rect 15292 13175 15344 13184
rect 15292 13141 15301 13175
rect 15301 13141 15335 13175
rect 15335 13141 15344 13175
rect 15292 13132 15344 13141
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2504 12928 2556 12980
rect 3332 12928 3384 12980
rect 3424 12792 3476 12844
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 3884 12724 3936 12776
rect 2688 12656 2740 12708
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4804 12928 4856 12980
rect 7656 12928 7708 12980
rect 6460 12835 6512 12844
rect 6460 12801 6469 12835
rect 6469 12801 6503 12835
rect 6503 12801 6512 12835
rect 6460 12792 6512 12801
rect 10508 12928 10560 12980
rect 11980 12928 12032 12980
rect 12256 12928 12308 12980
rect 13544 12928 13596 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 7840 12724 7892 12776
rect 6736 12699 6788 12708
rect 6736 12665 6770 12699
rect 6770 12665 6788 12699
rect 6736 12656 6788 12665
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 10692 12792 10744 12844
rect 11796 12792 11848 12844
rect 15660 12792 15712 12844
rect 9864 12724 9916 12776
rect 10048 12724 10100 12776
rect 12808 12724 12860 12776
rect 13728 12724 13780 12776
rect 16488 12724 16540 12776
rect 9404 12656 9456 12708
rect 14096 12656 14148 12708
rect 14648 12699 14700 12708
rect 14648 12665 14682 12699
rect 14682 12665 14700 12699
rect 14648 12656 14700 12665
rect 9496 12588 9548 12640
rect 10784 12588 10836 12640
rect 12716 12588 12768 12640
rect 13360 12588 13412 12640
rect 13636 12631 13688 12640
rect 13636 12597 13645 12631
rect 13645 12597 13679 12631
rect 13679 12597 13688 12631
rect 13636 12588 13688 12597
rect 16396 12656 16448 12708
rect 21364 12656 21416 12708
rect 15936 12588 15988 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 16304 12631 16356 12640
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 1952 12384 2004 12436
rect 2136 12384 2188 12436
rect 2688 12384 2740 12436
rect 5632 12384 5684 12436
rect 7104 12384 7156 12436
rect 7380 12384 7432 12436
rect 8668 12384 8720 12436
rect 11796 12384 11848 12436
rect 12164 12384 12216 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 14648 12384 14700 12436
rect 15292 12384 15344 12436
rect 3976 12316 4028 12368
rect 4252 12316 4304 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1860 12248 1912 12300
rect 2688 12248 2740 12300
rect 6920 12316 6972 12368
rect 9128 12316 9180 12368
rect 9496 12316 9548 12368
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 5356 12180 5408 12232
rect 7472 12248 7524 12300
rect 8208 12248 8260 12300
rect 13268 12316 13320 12368
rect 6828 12180 6880 12232
rect 10692 12180 10744 12232
rect 11796 12248 11848 12300
rect 8668 12112 8720 12164
rect 9312 12112 9364 12164
rect 12072 12112 12124 12164
rect 3056 12044 3108 12096
rect 3884 12044 3936 12096
rect 6828 12044 6880 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11060 12044 11112 12096
rect 13820 12248 13872 12300
rect 15476 12291 15528 12300
rect 15476 12257 15494 12291
rect 15494 12257 15528 12291
rect 15476 12248 15528 12257
rect 15660 12248 15712 12300
rect 16488 12316 16540 12368
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 14004 12044 14056 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2320 11883 2372 11892
rect 2320 11849 2329 11883
rect 2329 11849 2363 11883
rect 2363 11849 2372 11883
rect 2320 11840 2372 11849
rect 3240 11840 3292 11892
rect 7196 11840 7248 11892
rect 7380 11840 7432 11892
rect 3976 11772 4028 11824
rect 7012 11772 7064 11824
rect 11796 11840 11848 11892
rect 12164 11840 12216 11892
rect 12348 11840 12400 11892
rect 12532 11883 12584 11892
rect 12532 11849 12541 11883
rect 12541 11849 12575 11883
rect 12575 11849 12584 11883
rect 12532 11840 12584 11849
rect 16212 11840 16264 11892
rect 13176 11772 13228 11824
rect 2136 11704 2188 11756
rect 2688 11704 2740 11756
rect 4068 11704 4120 11756
rect 6828 11704 6880 11756
rect 6920 11704 6972 11756
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9220 11704 9272 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 10876 11704 10928 11756
rect 11060 11704 11112 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12072 11704 12124 11756
rect 14648 11704 14700 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 3884 11636 3936 11688
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 2320 11500 2372 11552
rect 3608 11568 3660 11620
rect 5264 11636 5316 11688
rect 6092 11636 6144 11688
rect 6276 11636 6328 11688
rect 4620 11568 4672 11620
rect 8944 11636 8996 11688
rect 9588 11636 9640 11688
rect 10232 11636 10284 11688
rect 7564 11568 7616 11620
rect 9680 11568 9732 11620
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 5264 11543 5316 11552
rect 5264 11509 5273 11543
rect 5273 11509 5307 11543
rect 5307 11509 5316 11543
rect 5264 11500 5316 11509
rect 5448 11500 5500 11552
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 8392 11500 8444 11552
rect 9588 11500 9640 11552
rect 10968 11568 11020 11620
rect 14280 11636 14332 11688
rect 16396 11636 16448 11688
rect 12624 11568 12676 11620
rect 12532 11500 12584 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 14740 11500 14792 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3240 11296 3292 11348
rect 4896 11296 4948 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 9588 11339 9640 11348
rect 9588 11305 9597 11339
rect 9597 11305 9631 11339
rect 9631 11305 9640 11339
rect 9588 11296 9640 11305
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 14556 11296 14608 11348
rect 1492 11160 1544 11212
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 4620 11160 4672 11212
rect 5908 11160 5960 11212
rect 6828 11203 6880 11212
rect 6828 11169 6862 11203
rect 6862 11169 6880 11203
rect 6828 11160 6880 11169
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 10324 11160 10376 11212
rect 11244 11160 11296 11212
rect 11888 11160 11940 11212
rect 12348 11160 12400 11212
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 1492 10956 1544 11008
rect 3148 11135 3200 11144
rect 2688 11024 2740 11076
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3884 11024 3936 11076
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5816 11092 5868 11144
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 5356 11024 5408 11076
rect 7564 11024 7616 11076
rect 9956 11092 10008 11144
rect 10876 11092 10928 11144
rect 10600 11024 10652 11076
rect 12716 11092 12768 11144
rect 14372 11228 14424 11280
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 15476 11092 15528 11144
rect 17132 11024 17184 11076
rect 3332 10999 3384 11008
rect 3332 10965 3341 10999
rect 3341 10965 3375 10999
rect 3375 10965 3384 10999
rect 3332 10956 3384 10965
rect 11796 10956 11848 11008
rect 12072 10956 12124 11008
rect 12348 10956 12400 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 12900 10956 12952 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 4988 10752 5040 10804
rect 5264 10752 5316 10804
rect 8576 10752 8628 10804
rect 10324 10752 10376 10804
rect 10968 10752 11020 10804
rect 2964 10684 3016 10736
rect 14464 10752 14516 10804
rect 16580 10684 16632 10736
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5356 10616 5408 10668
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 6552 10616 6604 10668
rect 6828 10616 6880 10668
rect 7564 10659 7616 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 3976 10548 4028 10600
rect 4344 10548 4396 10600
rect 5448 10548 5500 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 8392 10591 8444 10600
rect 2504 10480 2556 10532
rect 7012 10480 7064 10532
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 4160 10412 4212 10464
rect 4620 10455 4672 10464
rect 4620 10421 4629 10455
rect 4629 10421 4663 10455
rect 4663 10421 4672 10455
rect 4620 10412 4672 10421
rect 5264 10412 5316 10464
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 8484 10548 8536 10600
rect 9128 10548 9180 10600
rect 11244 10616 11296 10668
rect 15016 10616 15068 10668
rect 12624 10480 12676 10532
rect 12808 10480 12860 10532
rect 12900 10480 12952 10532
rect 13084 10480 13136 10532
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10968 10455 11020 10464
rect 10324 10412 10376 10421
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 11888 10412 11940 10464
rect 12440 10412 12492 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 14740 10412 14792 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2044 10208 2096 10260
rect 2228 10208 2280 10260
rect 2688 10208 2740 10260
rect 4252 10208 4304 10260
rect 4620 10208 4672 10260
rect 7656 10208 7708 10260
rect 10048 10208 10100 10260
rect 11244 10208 11296 10260
rect 3700 10140 3752 10192
rect 4896 10140 4948 10192
rect 6828 10140 6880 10192
rect 1492 10072 1544 10124
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 3608 10072 3660 10124
rect 5816 10072 5868 10124
rect 6460 10072 6512 10124
rect 3976 10004 4028 10056
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6736 9936 6788 9988
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 10232 10140 10284 10192
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9128 10004 9180 10056
rect 9772 10004 9824 10056
rect 10232 10004 10284 10056
rect 11060 10004 11112 10056
rect 12992 10140 13044 10192
rect 12440 10072 12492 10124
rect 13452 10072 13504 10124
rect 14096 10140 14148 10192
rect 16120 10072 16172 10124
rect 13176 10004 13228 10056
rect 14648 10004 14700 10056
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 9312 9936 9364 9988
rect 4896 9868 4948 9920
rect 5908 9868 5960 9920
rect 9220 9868 9272 9920
rect 11060 9868 11112 9920
rect 12348 9868 12400 9920
rect 12716 9868 12768 9920
rect 12900 9868 12952 9920
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 3700 9664 3752 9716
rect 9220 9664 9272 9716
rect 2320 9528 2372 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 1584 9460 1636 9512
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 3792 9596 3844 9648
rect 4896 9639 4948 9648
rect 4896 9605 4905 9639
rect 4905 9605 4939 9639
rect 4939 9605 4948 9639
rect 4896 9596 4948 9605
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 8484 9596 8536 9648
rect 10324 9664 10376 9716
rect 10968 9596 11020 9648
rect 4160 9528 4212 9580
rect 4804 9528 4856 9580
rect 5264 9528 5316 9580
rect 5724 9528 5776 9580
rect 4252 9460 4304 9512
rect 5908 9460 5960 9512
rect 6184 9503 6236 9512
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 8300 9528 8352 9580
rect 10692 9528 10744 9580
rect 11060 9571 11112 9580
rect 11060 9537 11069 9571
rect 11069 9537 11103 9571
rect 11103 9537 11112 9571
rect 11060 9528 11112 9537
rect 7472 9392 7524 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 2872 9324 2924 9376
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3516 9324 3568 9376
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5540 9324 5592 9376
rect 5816 9324 5868 9376
rect 8392 9460 8444 9512
rect 9956 9460 10008 9512
rect 12532 9596 12584 9648
rect 12900 9528 12952 9580
rect 13912 9596 13964 9648
rect 14096 9528 14148 9580
rect 9128 9392 9180 9444
rect 11060 9392 11112 9444
rect 11796 9392 11848 9444
rect 13452 9460 13504 9512
rect 13544 9460 13596 9512
rect 18696 9392 18748 9444
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 12164 9324 12216 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1676 9120 1728 9172
rect 3884 9120 3936 9172
rect 5080 9120 5132 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 7748 9120 7800 9172
rect 1584 9052 1636 9104
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 1400 8984 1452 8993
rect 2044 8984 2096 9036
rect 3516 8984 3568 9036
rect 4896 8984 4948 9036
rect 8300 9120 8352 9172
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 10140 9052 10192 9104
rect 10232 9095 10284 9104
rect 10232 9061 10250 9095
rect 10250 9061 10284 9095
rect 10508 9120 10560 9172
rect 12164 9163 12216 9172
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 13544 9120 13596 9172
rect 14556 9120 14608 9172
rect 10232 9052 10284 9061
rect 13268 9052 13320 9104
rect 2136 8916 2188 8968
rect 2596 8916 2648 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3976 8916 4028 8968
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 8116 8916 8168 8968
rect 3700 8823 3752 8832
rect 3700 8789 3709 8823
rect 3709 8789 3743 8823
rect 3743 8789 3752 8823
rect 3700 8780 3752 8789
rect 4252 8780 4304 8832
rect 7472 8848 7524 8900
rect 8392 8916 8444 8968
rect 8668 8916 8720 8968
rect 9404 8916 9456 8968
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 10324 8780 10376 8832
rect 10968 8984 11020 9036
rect 10876 8916 10928 8968
rect 12900 8984 12952 9036
rect 17132 9052 17184 9104
rect 13636 9027 13688 9036
rect 12164 8916 12216 8968
rect 12256 8848 12308 8900
rect 12716 8848 12768 8900
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 14004 8916 14056 8968
rect 13912 8848 13964 8900
rect 12440 8780 12492 8832
rect 13728 8780 13780 8832
rect 15292 8848 15344 8900
rect 15200 8780 15252 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 4896 8576 4948 8628
rect 5540 8619 5592 8628
rect 4436 8440 4488 8492
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5080 8440 5132 8492
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2688 8372 2740 8424
rect 3148 8372 3200 8424
rect 1492 8304 1544 8356
rect 2872 8304 2924 8356
rect 3976 8372 4028 8424
rect 3700 8304 3752 8356
rect 2596 8236 2648 8288
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 4252 8236 4304 8288
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 6184 8576 6236 8628
rect 6736 8576 6788 8628
rect 8668 8576 8720 8628
rect 7656 8508 7708 8560
rect 8852 8508 8904 8560
rect 9496 8576 9548 8628
rect 11152 8576 11204 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 10600 8508 10652 8560
rect 10784 8508 10836 8560
rect 6184 8440 6236 8492
rect 9128 8440 9180 8492
rect 9404 8440 9456 8492
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10232 8440 10284 8492
rect 10324 8440 10376 8492
rect 10968 8440 11020 8492
rect 12164 8508 12216 8560
rect 12256 8508 12308 8560
rect 14740 8508 14792 8560
rect 7656 8372 7708 8424
rect 9036 8372 9088 8424
rect 12716 8440 12768 8492
rect 12808 8440 12860 8492
rect 7012 8304 7064 8356
rect 4896 8236 4948 8288
rect 5264 8236 5316 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 7288 8304 7340 8356
rect 8208 8304 8260 8356
rect 10140 8304 10192 8356
rect 12992 8372 13044 8424
rect 13268 8372 13320 8424
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14556 8372 14608 8424
rect 15660 8372 15712 8424
rect 12716 8347 12768 8356
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 11060 8236 11112 8245
rect 11152 8236 11204 8288
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 13360 8304 13412 8356
rect 13820 8304 13872 8356
rect 14188 8304 14240 8356
rect 15200 8304 15252 8356
rect 16396 8304 16448 8356
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 13544 8236 13596 8245
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1584 8032 1636 8084
rect 12716 8032 12768 8084
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 2136 7964 2188 8016
rect 2596 7964 2648 8016
rect 4068 7964 4120 8016
rect 5264 7964 5316 8016
rect 6184 7964 6236 8016
rect 7104 7964 7156 8016
rect 7656 7964 7708 8016
rect 9772 7964 9824 8016
rect 10692 8007 10744 8016
rect 10692 7973 10726 8007
rect 10726 7973 10744 8007
rect 10692 7964 10744 7973
rect 11060 7964 11112 8016
rect 11796 7964 11848 8016
rect 2872 7896 2924 7948
rect 2964 7896 3016 7948
rect 5816 7939 5868 7948
rect 3148 7828 3200 7880
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 7288 7896 7340 7948
rect 7380 7896 7432 7948
rect 8944 7896 8996 7948
rect 9496 7896 9548 7948
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 12808 7939 12860 7948
rect 12808 7905 12842 7939
rect 12842 7905 12860 7939
rect 12808 7896 12860 7905
rect 13728 7896 13780 7948
rect 15844 7964 15896 8016
rect 4436 7803 4488 7812
rect 4436 7769 4445 7803
rect 4445 7769 4479 7803
rect 4479 7769 4488 7803
rect 4436 7760 4488 7769
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 3424 7692 3476 7744
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 6276 7828 6328 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 8300 7828 8352 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10324 7828 10376 7880
rect 5816 7760 5868 7812
rect 5908 7760 5960 7812
rect 7748 7760 7800 7812
rect 8668 7760 8720 7812
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 6092 7692 6144 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7104 7692 7156 7744
rect 7656 7692 7708 7744
rect 11152 7692 11204 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 15752 7735 15804 7744
rect 15752 7701 15761 7735
rect 15761 7701 15795 7735
rect 15795 7701 15804 7735
rect 15752 7692 15804 7701
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 17224 7692 17276 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 3240 7488 3292 7540
rect 3884 7488 3936 7540
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3148 7352 3200 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 3332 7284 3384 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 5816 7488 5868 7540
rect 7380 7488 7432 7540
rect 8484 7488 8536 7540
rect 10784 7488 10836 7540
rect 4712 7420 4764 7472
rect 5080 7420 5132 7472
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 6460 7352 6512 7404
rect 7196 7420 7248 7472
rect 6552 7284 6604 7336
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 12348 7352 12400 7404
rect 13912 7352 13964 7404
rect 14556 7352 14608 7404
rect 15752 7352 15804 7404
rect 6920 7284 6972 7336
rect 9496 7284 9548 7336
rect 12256 7284 12308 7336
rect 15292 7327 15344 7336
rect 3516 7216 3568 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 2228 7148 2280 7200
rect 2412 7148 2464 7200
rect 3240 7148 3292 7200
rect 4344 7148 4396 7200
rect 5540 7148 5592 7200
rect 8300 7216 8352 7268
rect 8668 7216 8720 7268
rect 11060 7216 11112 7268
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 6828 7148 6880 7200
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10876 7148 10928 7200
rect 12900 7216 12952 7268
rect 14280 7148 14332 7200
rect 15384 7148 15436 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 1676 6944 1728 6996
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 5080 6944 5132 6996
rect 5264 6987 5316 6996
rect 5264 6953 5273 6987
rect 5273 6953 5307 6987
rect 5307 6953 5316 6987
rect 5264 6944 5316 6953
rect 7196 6944 7248 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 9680 6944 9732 6996
rect 9864 6944 9916 6996
rect 10324 6944 10376 6996
rect 10692 6944 10744 6996
rect 3424 6876 3476 6928
rect 4988 6876 5040 6928
rect 1492 6808 1544 6860
rect 1308 6740 1360 6792
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 2872 6808 2924 6860
rect 3332 6808 3384 6860
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 3332 6604 3384 6656
rect 3700 6647 3752 6656
rect 3700 6613 3709 6647
rect 3709 6613 3743 6647
rect 3743 6613 3752 6647
rect 3700 6604 3752 6613
rect 4804 6808 4856 6860
rect 5632 6876 5684 6928
rect 6368 6876 6420 6928
rect 10968 6944 11020 6996
rect 14740 6987 14792 6996
rect 4988 6740 5040 6792
rect 5724 6808 5776 6860
rect 7472 6808 7524 6860
rect 11060 6876 11112 6928
rect 11796 6876 11848 6928
rect 14740 6953 14749 6987
rect 14749 6953 14783 6987
rect 14783 6953 14792 6987
rect 14740 6944 14792 6953
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 9772 6808 9824 6860
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 4804 6604 4856 6656
rect 7932 6672 7984 6724
rect 8668 6672 8720 6724
rect 9772 6672 9824 6724
rect 12164 6808 12216 6860
rect 14464 6808 14516 6860
rect 19064 6808 19116 6860
rect 9956 6740 10008 6792
rect 10968 6740 11020 6792
rect 12532 6740 12584 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 10692 6672 10744 6724
rect 10784 6604 10836 6656
rect 12440 6672 12492 6724
rect 16304 6672 16356 6724
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 15476 6604 15528 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 3332 6400 3384 6452
rect 3608 6400 3660 6452
rect 6828 6400 6880 6452
rect 7748 6400 7800 6452
rect 4160 6332 4212 6384
rect 1676 6196 1728 6248
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 1768 6128 1820 6180
rect 3148 6128 3200 6180
rect 4712 6264 4764 6316
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5080 6264 5132 6316
rect 4528 6196 4580 6248
rect 10508 6375 10560 6384
rect 10508 6341 10517 6375
rect 10517 6341 10551 6375
rect 10551 6341 10560 6375
rect 10508 6332 10560 6341
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 7196 6307 7248 6316
rect 5724 6239 5776 6248
rect 5724 6205 5733 6239
rect 5733 6205 5767 6239
rect 5767 6205 5776 6239
rect 5724 6196 5776 6205
rect 6000 6196 6052 6248
rect 6736 6239 6788 6248
rect 6736 6205 6745 6239
rect 6745 6205 6779 6239
rect 6779 6205 6788 6239
rect 6736 6196 6788 6205
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 7472 6264 7524 6316
rect 12256 6332 12308 6384
rect 7748 6196 7800 6248
rect 10784 6264 10836 6316
rect 12900 6332 12952 6384
rect 10692 6196 10744 6248
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 5264 6128 5316 6180
rect 6828 6128 6880 6180
rect 7288 6171 7340 6180
rect 7288 6137 7297 6171
rect 7297 6137 7331 6171
rect 7331 6137 7340 6171
rect 7288 6128 7340 6137
rect 1400 6060 1452 6112
rect 3608 6060 3660 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4896 6060 4948 6112
rect 6000 6060 6052 6112
rect 6184 6060 6236 6112
rect 6736 6060 6788 6112
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 10232 6128 10284 6180
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8760 6060 8812 6112
rect 9220 6060 9272 6112
rect 12256 6060 12308 6112
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 14464 6128 14516 6180
rect 17408 6128 17460 6180
rect 12808 6060 12860 6112
rect 14280 6060 14332 6112
rect 14648 6060 14700 6112
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 17868 6060 17920 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 3148 5856 3200 5908
rect 2412 5788 2464 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3792 5856 3844 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 5448 5856 5500 5908
rect 6000 5856 6052 5908
rect 7196 5856 7248 5908
rect 7288 5856 7340 5908
rect 10232 5856 10284 5908
rect 10876 5856 10928 5908
rect 10968 5856 11020 5908
rect 4344 5831 4396 5840
rect 4344 5797 4353 5831
rect 4353 5797 4387 5831
rect 4387 5797 4396 5831
rect 4344 5788 4396 5797
rect 5540 5788 5592 5840
rect 6644 5788 6696 5840
rect 7472 5788 7524 5840
rect 4988 5763 5040 5772
rect 3424 5720 3476 5729
rect 4528 5695 4580 5704
rect 4528 5661 4537 5695
rect 4537 5661 4571 5695
rect 4571 5661 4580 5695
rect 4528 5652 4580 5661
rect 4988 5729 5022 5763
rect 5022 5729 5040 5763
rect 4988 5720 5040 5729
rect 5724 5720 5776 5772
rect 7932 5720 7984 5772
rect 8116 5788 8168 5840
rect 9956 5788 10008 5840
rect 11060 5788 11112 5840
rect 7840 5695 7892 5704
rect 4252 5584 4304 5636
rect 3792 5516 3844 5568
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 12072 5856 12124 5908
rect 14372 5856 14424 5908
rect 11980 5788 12032 5840
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 11060 5652 11112 5704
rect 5908 5584 5960 5636
rect 6092 5516 6144 5568
rect 6644 5516 6696 5568
rect 6736 5516 6788 5568
rect 7840 5516 7892 5568
rect 7932 5516 7984 5568
rect 10784 5516 10836 5568
rect 12072 5720 12124 5772
rect 12532 5720 12584 5772
rect 13084 5788 13136 5840
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 15292 5788 15344 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 14832 5720 14884 5772
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14740 5652 14792 5704
rect 15200 5584 15252 5636
rect 21548 5763 21600 5772
rect 21548 5729 21557 5763
rect 21557 5729 21591 5763
rect 21591 5729 21600 5763
rect 21548 5720 21600 5729
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 17592 5584 17644 5636
rect 14372 5516 14424 5568
rect 15568 5516 15620 5568
rect 17500 5559 17552 5568
rect 17500 5525 17509 5559
rect 17509 5525 17543 5559
rect 17543 5525 17552 5559
rect 17500 5516 17552 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 1492 5151 1544 5160
rect 1492 5117 1501 5151
rect 1501 5117 1535 5151
rect 1535 5117 1544 5151
rect 4160 5312 4212 5364
rect 5356 5312 5408 5364
rect 5448 5312 5500 5364
rect 8208 5312 8260 5364
rect 1860 5244 1912 5296
rect 7472 5287 7524 5296
rect 3148 5176 3200 5228
rect 3332 5176 3384 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4528 5176 4580 5228
rect 4988 5176 5040 5228
rect 6184 5176 6236 5228
rect 7196 5176 7248 5228
rect 1492 5108 1544 5117
rect 1768 5108 1820 5160
rect 2136 5151 2188 5160
rect 2136 5117 2170 5151
rect 2170 5117 2188 5151
rect 2136 5108 2188 5117
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 3976 5040 4028 5092
rect 6000 5108 6052 5160
rect 6644 5108 6696 5160
rect 5816 5040 5868 5092
rect 6368 5040 6420 5092
rect 7196 5040 7248 5092
rect 7472 5253 7481 5287
rect 7481 5253 7515 5287
rect 7515 5253 7524 5287
rect 7472 5244 7524 5253
rect 9404 5244 9456 5296
rect 12532 5244 12584 5296
rect 16488 5244 16540 5296
rect 17592 5244 17644 5296
rect 10232 5176 10284 5228
rect 11060 5176 11112 5228
rect 11796 5176 11848 5228
rect 12716 5176 12768 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 15200 5176 15252 5228
rect 7840 5108 7892 5160
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 10876 5108 10928 5160
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 3332 4972 3384 5024
rect 4068 4972 4120 5024
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6092 4972 6144 5024
rect 7288 4972 7340 5024
rect 8760 5040 8812 5092
rect 9036 5083 9088 5092
rect 9036 5049 9045 5083
rect 9045 5049 9079 5083
rect 9079 5049 9088 5083
rect 9036 5040 9088 5049
rect 11980 5040 12032 5092
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 13636 5040 13688 5092
rect 15476 5040 15528 5092
rect 17224 5176 17276 5228
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 17316 5108 17368 5117
rect 18144 5108 18196 5160
rect 14280 4972 14332 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14740 4972 14792 5024
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17132 4972 17184 5024
rect 19984 4972 20036 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1032 4700 1084 4752
rect 1676 4700 1728 4752
rect 3148 4768 3200 4820
rect 3424 4768 3476 4820
rect 2136 4632 2188 4684
rect 1860 4564 1912 4616
rect 2504 4607 2556 4616
rect 2504 4573 2513 4607
rect 2513 4573 2547 4607
rect 2547 4573 2556 4607
rect 2504 4564 2556 4573
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 3056 4632 3108 4684
rect 3700 4632 3752 4684
rect 5356 4768 5408 4820
rect 3884 4632 3936 4684
rect 3976 4632 4028 4684
rect 4528 4632 4580 4684
rect 5632 4675 5684 4684
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7380 4768 7432 4820
rect 7656 4768 7708 4820
rect 8392 4768 8444 4820
rect 9036 4768 9088 4820
rect 9772 4768 9824 4820
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 10508 4768 10560 4820
rect 11152 4768 11204 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12256 4768 12308 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14740 4768 14792 4820
rect 15292 4768 15344 4820
rect 17500 4768 17552 4820
rect 9220 4700 9272 4752
rect 9496 4700 9548 4752
rect 12532 4743 12584 4752
rect 12532 4709 12541 4743
rect 12541 4709 12575 4743
rect 12575 4709 12584 4743
rect 12532 4700 12584 4709
rect 14464 4700 14516 4752
rect 15568 4743 15620 4752
rect 5632 4641 5661 4675
rect 5661 4641 5684 4675
rect 5632 4632 5684 4641
rect 2596 4564 2648 4573
rect 3792 4564 3844 4616
rect 2320 4496 2372 4548
rect 3148 4496 3200 4548
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6460 4632 6512 4684
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 7380 4632 7432 4684
rect 8300 4675 8352 4684
rect 6828 4564 6880 4616
rect 7012 4564 7064 4616
rect 7564 4564 7616 4616
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8392 4632 8444 4684
rect 10508 4632 10560 4684
rect 10876 4632 10928 4684
rect 11980 4632 12032 4684
rect 3424 4471 3476 4480
rect 3424 4437 3433 4471
rect 3433 4437 3467 4471
rect 3467 4437 3476 4471
rect 3424 4428 3476 4437
rect 3700 4428 3752 4480
rect 4344 4428 4396 4480
rect 7288 4496 7340 4548
rect 7472 4496 7524 4548
rect 8760 4564 8812 4616
rect 6276 4428 6328 4480
rect 6460 4471 6512 4480
rect 6460 4437 6469 4471
rect 6469 4437 6503 4471
rect 6503 4437 6512 4471
rect 6460 4428 6512 4437
rect 6552 4428 6604 4480
rect 10140 4496 10192 4548
rect 10692 4496 10744 4548
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 13636 4564 13688 4616
rect 14556 4632 14608 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 15568 4709 15577 4743
rect 15577 4709 15611 4743
rect 15611 4709 15620 4743
rect 15568 4700 15620 4709
rect 16948 4700 17000 4752
rect 14924 4632 14976 4684
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 16488 4564 16540 4616
rect 17408 4564 17460 4616
rect 12072 4496 12124 4548
rect 12440 4496 12492 4548
rect 13360 4496 13412 4548
rect 15476 4496 15528 4548
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 12532 4428 12584 4480
rect 15200 4471 15252 4480
rect 15200 4437 15209 4471
rect 15209 4437 15243 4471
rect 15243 4437 15252 4471
rect 15200 4428 15252 4437
rect 17132 4428 17184 4480
rect 20996 4428 21048 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2688 4224 2740 4276
rect 3424 4224 3476 4276
rect 4344 4224 4396 4276
rect 5632 4224 5684 4276
rect 5816 4224 5868 4276
rect 8116 4224 8168 4276
rect 9036 4224 9088 4276
rect 2872 4156 2924 4208
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 1216 4020 1268 4072
rect 1584 4020 1636 4072
rect 3056 4020 3108 4072
rect 3148 4020 3200 4072
rect 3424 4020 3476 4072
rect 4620 4088 4672 4140
rect 3700 4020 3752 4072
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 4068 4063 4120 4072
rect 3792 4020 3844 4029
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 6000 4156 6052 4208
rect 6276 4156 6328 4208
rect 6920 4088 6972 4140
rect 5908 4020 5960 4072
rect 6736 4020 6788 4072
rect 8760 4156 8812 4208
rect 11060 4224 11112 4276
rect 12256 4224 12308 4276
rect 13084 4224 13136 4276
rect 13636 4267 13688 4276
rect 9680 4156 9732 4208
rect 7656 4088 7708 4140
rect 8300 4088 8352 4140
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 10232 4088 10284 4140
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 10968 4088 11020 4140
rect 12348 4156 12400 4208
rect 13360 4156 13412 4208
rect 13636 4233 13645 4267
rect 13645 4233 13679 4267
rect 13679 4233 13688 4267
rect 13636 4224 13688 4233
rect 8668 4063 8720 4072
rect 2044 3995 2096 4004
rect 2044 3961 2078 3995
rect 2078 3961 2096 3995
rect 2044 3952 2096 3961
rect 2596 3884 2648 3936
rect 3056 3884 3108 3936
rect 3332 3884 3384 3936
rect 4712 3952 4764 4004
rect 3516 3884 3568 3936
rect 4988 3884 5040 3936
rect 5080 3884 5132 3936
rect 6276 3952 6328 4004
rect 7380 3952 7432 4004
rect 8116 3952 8168 4004
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7288 3884 7340 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 12440 4088 12492 4140
rect 13268 4131 13320 4140
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 15108 4224 15160 4276
rect 8760 3952 8812 4004
rect 12256 4020 12308 4072
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9864 3884 9916 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 14924 4020 14976 4072
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 11060 3884 11112 3936
rect 11980 3884 12032 3936
rect 14740 3995 14792 4004
rect 14740 3961 14758 3995
rect 14758 3961 14792 3995
rect 14740 3952 14792 3961
rect 12716 3884 12768 3936
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 14372 3884 14424 3936
rect 18052 3884 18104 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2504 3680 2556 3732
rect 2964 3680 3016 3732
rect 3792 3680 3844 3732
rect 3976 3680 4028 3732
rect 4804 3680 4856 3732
rect 5816 3680 5868 3732
rect 6920 3680 6972 3732
rect 2780 3655 2832 3664
rect 2780 3621 2820 3655
rect 2820 3621 2832 3655
rect 2780 3612 2832 3621
rect 3056 3612 3108 3664
rect 3700 3612 3752 3664
rect 4620 3612 4672 3664
rect 4712 3612 4764 3664
rect 7564 3680 7616 3732
rect 8300 3680 8352 3732
rect 8484 3680 8536 3732
rect 8576 3680 8628 3732
rect 9036 3680 9088 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 10048 3680 10100 3732
rect 11888 3680 11940 3732
rect 12072 3723 12124 3732
rect 12072 3689 12081 3723
rect 12081 3689 12115 3723
rect 12115 3689 12124 3723
rect 12072 3680 12124 3689
rect 12164 3680 12216 3732
rect 14096 3723 14148 3732
rect 8024 3612 8076 3664
rect 8208 3612 8260 3664
rect 1308 3544 1360 3596
rect 2504 3544 2556 3596
rect 3148 3544 3200 3596
rect 3332 3544 3384 3596
rect 4528 3544 4580 3596
rect 4896 3544 4948 3596
rect 3792 3408 3844 3460
rect 5632 3408 5684 3460
rect 6552 3544 6604 3596
rect 6736 3476 6788 3528
rect 7472 3544 7524 3596
rect 1676 3383 1728 3392
rect 1676 3349 1685 3383
rect 1685 3349 1719 3383
rect 1719 3349 1728 3383
rect 1676 3340 1728 3349
rect 1952 3340 2004 3392
rect 2044 3340 2096 3392
rect 2872 3340 2924 3392
rect 3240 3340 3292 3392
rect 6828 3408 6880 3460
rect 7748 3408 7800 3460
rect 8300 3476 8352 3528
rect 8576 3544 8628 3596
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 10232 3544 10284 3596
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 14648 3680 14700 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 18144 3680 18196 3732
rect 12440 3587 12492 3596
rect 12440 3553 12449 3587
rect 12449 3553 12483 3587
rect 12483 3553 12492 3587
rect 12440 3544 12492 3553
rect 9220 3476 9272 3528
rect 9588 3476 9640 3528
rect 11888 3476 11940 3528
rect 12348 3476 12400 3528
rect 14004 3612 14056 3664
rect 15568 3612 15620 3664
rect 9772 3408 9824 3460
rect 13084 3587 13136 3596
rect 13084 3553 13093 3587
rect 13093 3553 13127 3587
rect 13127 3553 13136 3587
rect 13084 3544 13136 3553
rect 14096 3544 14148 3596
rect 15384 3587 15436 3596
rect 14924 3519 14976 3528
rect 14924 3485 14933 3519
rect 14933 3485 14967 3519
rect 14967 3485 14976 3519
rect 14924 3476 14976 3485
rect 15384 3553 15393 3587
rect 15393 3553 15427 3587
rect 15427 3553 15436 3587
rect 15384 3544 15436 3553
rect 20168 3612 20220 3664
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 12808 3408 12860 3460
rect 14280 3408 14332 3460
rect 15384 3408 15436 3460
rect 19156 3408 19208 3460
rect 7472 3340 7524 3392
rect 8576 3340 8628 3392
rect 9588 3340 9640 3392
rect 11152 3340 11204 3392
rect 12164 3340 12216 3392
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 13544 3340 13596 3392
rect 15752 3340 15804 3392
rect 19064 3340 19116 3392
rect 19708 3340 19760 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 1584 3136 1636 3188
rect 2688 3136 2740 3188
rect 2412 3000 2464 3052
rect 2780 3000 2832 3052
rect 3976 3068 4028 3120
rect 1492 2975 1544 2984
rect 1492 2941 1501 2975
rect 1501 2941 1535 2975
rect 1535 2941 1544 2975
rect 1492 2932 1544 2941
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4160 3136 4212 3188
rect 6276 3136 6328 3188
rect 7380 3136 7432 3188
rect 9220 3136 9272 3188
rect 9680 3136 9732 3188
rect 10232 3136 10284 3188
rect 10416 3136 10468 3188
rect 11704 3136 11756 3188
rect 14924 3136 14976 3188
rect 15384 3136 15436 3188
rect 4252 3068 4304 3120
rect 6092 3068 6144 3120
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 5632 3043 5684 3052
rect 4988 3000 5040 3009
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 7288 3068 7340 3120
rect 10140 3068 10192 3120
rect 6920 3000 6972 3052
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 10232 3000 10284 3052
rect 11888 3000 11940 3052
rect 15476 3068 15528 3120
rect 16764 3136 16816 3188
rect 16856 3136 16908 3188
rect 13268 3000 13320 3052
rect 6000 2932 6052 2984
rect 9220 2975 9272 2984
rect 9220 2941 9254 2975
rect 9254 2941 9272 2975
rect 9220 2932 9272 2941
rect 9588 2932 9640 2984
rect 10324 2932 10376 2984
rect 10508 2975 10560 2984
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 11244 2932 11296 2984
rect 11428 2932 11480 2984
rect 12164 2932 12216 2984
rect 12348 2932 12400 2984
rect 13360 2932 13412 2984
rect 14372 3000 14424 3052
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 15752 3000 15804 3052
rect 15568 2975 15620 2984
rect 204 2796 256 2848
rect 1308 2796 1360 2848
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 3700 2796 3752 2848
rect 3792 2796 3844 2848
rect 4252 2796 4304 2848
rect 5448 2864 5500 2916
rect 8024 2864 8076 2916
rect 8300 2864 8352 2916
rect 8760 2864 8812 2916
rect 4620 2796 4672 2848
rect 5540 2796 5592 2848
rect 6552 2796 6604 2848
rect 10232 2864 10284 2916
rect 10968 2864 11020 2916
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 15660 2932 15712 2984
rect 16948 3068 17000 3120
rect 17960 3068 18012 3120
rect 19524 3068 19576 3120
rect 19984 3068 20036 3120
rect 20168 3111 20220 3120
rect 20168 3077 20177 3111
rect 20177 3077 20211 3111
rect 20211 3077 20220 3111
rect 20168 3068 20220 3077
rect 16396 2932 16448 2984
rect 17040 2932 17092 2984
rect 17868 2975 17920 2984
rect 17868 2941 17877 2975
rect 17877 2941 17911 2975
rect 17911 2941 17920 2975
rect 17868 2932 17920 2941
rect 18144 2932 18196 2984
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 17500 2907 17552 2916
rect 9496 2796 9548 2848
rect 10508 2796 10560 2848
rect 10784 2839 10836 2848
rect 10784 2805 10793 2839
rect 10793 2805 10827 2839
rect 10827 2805 10836 2839
rect 10784 2796 10836 2805
rect 10876 2796 10928 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14280 2796 14332 2848
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 15384 2796 15436 2848
rect 15660 2796 15712 2848
rect 17500 2873 17509 2907
rect 17509 2873 17543 2907
rect 17543 2873 17552 2907
rect 17500 2864 17552 2873
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18144 2839 18196 2848
rect 18144 2805 18153 2839
rect 18153 2805 18187 2839
rect 18187 2805 18196 2839
rect 18880 3000 18932 3052
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 19248 3000 19300 3052
rect 22192 3000 22244 3052
rect 20168 2932 20220 2984
rect 22652 2932 22704 2984
rect 21732 2864 21784 2916
rect 18144 2796 18196 2805
rect 19432 2796 19484 2848
rect 19708 2839 19760 2848
rect 19708 2805 19717 2839
rect 19717 2805 19751 2839
rect 19751 2805 19760 2839
rect 19708 2796 19760 2805
rect 20720 2796 20772 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 3516 2592 3568 2644
rect 3608 2592 3660 2644
rect 4068 2592 4120 2644
rect 4252 2592 4304 2644
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 4896 2592 4948 2644
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 6552 2592 6604 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 9220 2635 9272 2644
rect 9220 2601 9229 2635
rect 9229 2601 9263 2635
rect 9263 2601 9272 2635
rect 9220 2592 9272 2601
rect 9404 2592 9456 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 11980 2592 12032 2644
rect 12164 2592 12216 2644
rect 13084 2592 13136 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 14648 2592 14700 2644
rect 17224 2592 17276 2644
rect 1952 2524 2004 2576
rect 3332 2524 3384 2576
rect 3700 2524 3752 2576
rect 1124 2456 1176 2508
rect 1676 2388 1728 2440
rect 2136 2363 2188 2372
rect 2136 2329 2145 2363
rect 2145 2329 2179 2363
rect 2179 2329 2188 2363
rect 2136 2320 2188 2329
rect 3148 2456 3200 2508
rect 3792 2456 3844 2508
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 4252 2499 4304 2508
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 5816 2567 5868 2576
rect 5080 2499 5132 2508
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 4804 2388 4856 2440
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 6828 2567 6880 2576
rect 6828 2533 6837 2567
rect 6837 2533 6871 2567
rect 6871 2533 6880 2567
rect 6828 2524 6880 2533
rect 11152 2524 11204 2576
rect 12992 2524 13044 2576
rect 13912 2524 13964 2576
rect 14280 2524 14332 2576
rect 15476 2567 15528 2576
rect 15476 2533 15485 2567
rect 15485 2533 15519 2567
rect 15519 2533 15528 2567
rect 15476 2524 15528 2533
rect 15660 2524 15712 2576
rect 16764 2567 16816 2576
rect 16764 2533 16773 2567
rect 16773 2533 16807 2567
rect 16807 2533 16816 2567
rect 16764 2524 16816 2533
rect 16948 2524 17000 2576
rect 18144 2592 18196 2644
rect 18052 2524 18104 2576
rect 19156 2567 19208 2576
rect 19156 2533 19165 2567
rect 19165 2533 19199 2567
rect 19199 2533 19208 2567
rect 19156 2524 19208 2533
rect 19524 2524 19576 2576
rect 19984 2524 20036 2576
rect 20720 2524 20772 2576
rect 6276 2456 6328 2508
rect 6460 2456 6512 2508
rect 7104 2456 7156 2508
rect 8944 2456 8996 2508
rect 9128 2456 9180 2508
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 8760 2388 8812 2440
rect 9496 2388 9548 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 4160 2252 4212 2304
rect 6828 2252 6880 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 10048 2456 10100 2508
rect 11336 2499 11388 2508
rect 11336 2465 11345 2499
rect 11345 2465 11379 2499
rect 11379 2465 11388 2499
rect 11336 2456 11388 2465
rect 10784 2388 10836 2440
rect 11060 2388 11112 2440
rect 12348 2456 12400 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 13544 2456 13596 2508
rect 14464 2456 14516 2508
rect 15200 2456 15252 2508
rect 15384 2456 15436 2508
rect 17960 2456 18012 2508
rect 19432 2456 19484 2508
rect 20996 2499 21048 2508
rect 20996 2465 21005 2499
rect 21005 2465 21039 2499
rect 21039 2465 21048 2499
rect 20996 2456 21048 2465
rect 11244 2252 11296 2304
rect 11888 2252 11940 2304
rect 19248 2388 19300 2440
rect 13268 2320 13320 2372
rect 13728 2320 13780 2372
rect 14280 2320 14332 2372
rect 14740 2320 14792 2372
rect 15200 2320 15252 2372
rect 15660 2363 15712 2372
rect 15660 2329 15669 2363
rect 15669 2329 15703 2363
rect 15703 2329 15712 2363
rect 15660 2320 15712 2329
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 16580 2363 16632 2372
rect 16580 2329 16589 2363
rect 16589 2329 16623 2363
rect 16623 2329 16632 2363
rect 16580 2320 16632 2329
rect 17040 2320 17092 2372
rect 17960 2363 18012 2372
rect 17960 2329 17969 2363
rect 17969 2329 18003 2363
rect 18003 2329 18012 2363
rect 17960 2320 18012 2329
rect 18972 2363 19024 2372
rect 18972 2329 18981 2363
rect 18981 2329 19015 2363
rect 19015 2329 19024 2363
rect 18972 2320 19024 2329
rect 19432 2363 19484 2372
rect 19432 2329 19441 2363
rect 19441 2329 19475 2363
rect 19475 2329 19484 2363
rect 19432 2320 19484 2329
rect 19892 2363 19944 2372
rect 19892 2329 19901 2363
rect 19901 2329 19935 2363
rect 19935 2329 19944 2363
rect 19892 2320 19944 2329
rect 20352 2363 20404 2372
rect 20352 2329 20361 2363
rect 20361 2329 20395 2363
rect 20395 2329 20404 2363
rect 20352 2320 20404 2329
rect 20812 2363 20864 2372
rect 20812 2329 20821 2363
rect 20821 2329 20855 2363
rect 20855 2329 20864 2363
rect 20812 2320 20864 2329
rect 21272 2363 21324 2372
rect 21272 2329 21281 2363
rect 21281 2329 21315 2363
rect 21315 2329 21324 2363
rect 21272 2320 21324 2329
rect 15936 2252 15988 2304
rect 18604 2252 18656 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3148 2048 3200 2100
rect 5724 2048 5776 2100
rect 7104 2048 7156 2100
rect 13360 2048 13412 2100
rect 3792 1980 3844 2032
rect 6368 1980 6420 2032
rect 11428 1980 11480 2032
rect 12900 1980 12952 2032
rect 4068 1912 4120 1964
rect 6644 1912 6696 1964
rect 5172 1844 5224 1896
rect 11244 1844 11296 1896
rect 664 1776 716 1828
rect 4252 1776 4304 1828
rect 5816 1776 5868 1828
rect 6460 1776 6512 1828
rect 4160 1708 4212 1760
rect 5448 1708 5500 1760
rect 4344 1640 4396 1692
rect 8944 1640 8996 1692
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3238 22672 3294 22681
rect 3238 22607 3294 22616
rect 216 20398 244 22200
rect 204 20392 256 20398
rect 204 20334 256 20340
rect 676 19854 704 22200
rect 1136 20466 1164 22200
rect 1596 20482 1624 22200
rect 1766 21176 1822 21185
rect 1766 21111 1822 21120
rect 1124 20460 1176 20466
rect 1124 20402 1176 20408
rect 1504 20454 1624 20482
rect 664 19848 716 19854
rect 664 19790 716 19796
rect 1398 19816 1454 19825
rect 1398 19751 1400 19760
rect 1452 19751 1454 19760
rect 1400 19722 1452 19728
rect 1398 19272 1454 19281
rect 1398 19207 1400 19216
rect 1452 19207 1454 19216
rect 1400 19178 1452 19184
rect 1398 18864 1454 18873
rect 1398 18799 1400 18808
rect 1452 18799 1454 18808
rect 1400 18770 1452 18776
rect 1398 18320 1454 18329
rect 1504 18290 1532 20454
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19394 1624 20334
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1688 19825 1716 20266
rect 1780 20058 1808 21111
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1860 20256 1912 20262
rect 1858 20224 1860 20233
rect 1912 20224 1914 20233
rect 1858 20159 1914 20168
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1964 19514 1992 20266
rect 2056 20074 2084 22200
rect 2226 20768 2282 20777
rect 2226 20703 2282 20712
rect 2240 20602 2268 20703
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2056 20046 2176 20074
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1596 19366 1716 19394
rect 1584 19236 1636 19242
rect 1584 19178 1636 19184
rect 1596 18970 1624 19178
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1398 18255 1400 18264
rect 1452 18255 1454 18264
rect 1492 18284 1544 18290
rect 1400 18226 1452 18232
rect 1492 18226 1544 18232
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1490 17912 1546 17921
rect 1596 17882 1624 18090
rect 1490 17847 1492 17856
rect 1544 17847 1546 17856
rect 1584 17876 1636 17882
rect 1492 17818 1544 17824
rect 1584 17818 1636 17824
rect 1688 17202 1716 19366
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1780 18426 1808 18770
rect 1964 18426 1992 19246
rect 2056 18970 2084 19858
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2042 18864 2098 18873
rect 2042 18799 2044 18808
rect 2096 18799 2098 18808
rect 2044 18770 2096 18776
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2148 18222 2176 20046
rect 2332 19514 2360 20266
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2424 18970 2452 19858
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2516 18714 2544 22200
rect 2870 22128 2926 22137
rect 2870 22063 2926 22072
rect 2778 21720 2834 21729
rect 2778 21655 2834 21664
rect 2792 20602 2820 21655
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2884 20534 2912 22063
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2976 20482 3004 22200
rect 3252 20534 3280 22607
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 3240 20528 3292 20534
rect 2976 20454 3096 20482
rect 3240 20470 3292 20476
rect 2688 20324 2740 20330
rect 2688 20266 2740 20272
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2700 20058 2728 20266
rect 2780 20256 2832 20262
rect 2780 20198 2832 20204
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2792 18834 2820 20198
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2884 19514 2912 19858
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2136 18216 2188 18222
rect 2320 18216 2372 18222
rect 2136 18158 2188 18164
rect 2226 18184 2282 18193
rect 2320 18158 2372 18164
rect 2226 18119 2282 18128
rect 2240 18086 2268 18119
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 1858 17368 1914 17377
rect 2148 17338 2176 17546
rect 1858 17303 1860 17312
rect 1912 17303 1914 17312
rect 2136 17332 2188 17338
rect 1860 17274 1912 17280
rect 2136 17274 2188 17280
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1584 17060 1636 17066
rect 1584 17002 1636 17008
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1492 16992 1544 16998
rect 1490 16960 1492 16969
rect 1544 16960 1546 16969
rect 1490 16895 1546 16904
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1596 16250 1624 17002
rect 1964 16794 1992 17002
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2056 16658 2084 17206
rect 2228 17128 2280 17134
rect 2228 17070 2280 17076
rect 2240 16794 2268 17070
rect 2332 16794 2360 18158
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2424 16726 2452 18702
rect 2516 18686 2636 18714
rect 2976 18698 3004 20266
rect 3068 20040 3096 20454
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3068 20012 3280 20040
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 3068 19174 3096 19722
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2608 18630 2636 18686
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2504 18352 2556 18358
rect 2502 18320 2504 18329
rect 2556 18320 2558 18329
rect 2502 18255 2558 18264
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 17882 2544 18090
rect 2976 18086 3004 18362
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2884 17898 2912 18022
rect 2504 17876 2556 17882
rect 2884 17870 3096 17898
rect 3160 17882 3188 19858
rect 3252 18970 3280 20012
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3252 18630 3280 18770
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18426 3280 18566
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 2504 17818 2556 17824
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2976 17202 3004 17546
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3068 17134 3096 17870
rect 3148 17876 3200 17882
rect 3344 17864 3372 20266
rect 3436 20040 3464 22200
rect 3896 20602 3924 22200
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3528 20262 3556 20470
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3436 20012 3648 20040
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3148 17818 3200 17824
rect 3252 17836 3372 17864
rect 3252 17542 3280 17836
rect 3436 17746 3464 19858
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3528 19310 3556 19790
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3620 18970 3648 20012
rect 3712 19922 3740 20402
rect 4080 20398 4108 20538
rect 4356 20534 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4356 20398 4384 20470
rect 4816 20398 4844 22200
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3700 19916 3752 19922
rect 3700 19858 3752 19864
rect 3792 19236 3844 19242
rect 3792 19178 3844 19184
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3528 18834 3556 18906
rect 3516 18828 3568 18834
rect 3568 18788 3740 18816
rect 3516 18770 3568 18776
rect 3514 18728 3570 18737
rect 3514 18663 3516 18672
rect 3568 18663 3570 18672
rect 3516 18634 3568 18640
rect 3516 18148 3568 18154
rect 3516 18090 3568 18096
rect 3528 17882 3556 18090
rect 3712 18086 3740 18788
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3344 17338 3372 17682
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 3804 17066 3832 19178
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 2976 16794 3004 16934
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3436 16726 3464 16934
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1398 16008 1454 16017
rect 1398 15943 1400 15952
rect 1452 15943 1454 15952
rect 1584 15972 1636 15978
rect 1400 15914 1452 15920
rect 1584 15914 1636 15920
rect 1596 15706 1624 15914
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1398 15464 1454 15473
rect 1398 15399 1400 15408
rect 1452 15399 1454 15408
rect 1400 15370 1452 15376
rect 1688 15366 1716 16594
rect 1872 16250 1900 16594
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15706 1992 15982
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1964 15162 1992 15506
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1398 15056 1454 15065
rect 1398 14991 1400 15000
rect 1452 14991 1454 15000
rect 1400 14962 1452 14968
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1780 14618 1808 14826
rect 2056 14618 2084 15438
rect 2240 15162 2268 15506
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 1398 14512 1454 14521
rect 1398 14447 1400 14456
rect 1452 14447 1454 14456
rect 1952 14476 2004 14482
rect 1400 14418 1452 14424
rect 1952 14418 2004 14424
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 1490 14104 1546 14113
rect 1964 14074 1992 14418
rect 1490 14039 1492 14048
rect 1544 14039 1546 14048
rect 1952 14068 2004 14074
rect 1492 14010 1544 14016
rect 1952 14010 2004 14016
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1490 13560 1546 13569
rect 1490 13495 1492 13504
rect 1544 13495 1546 13504
rect 1492 13466 1544 13472
rect 1780 13462 1808 13670
rect 1768 13456 1820 13462
rect 1768 13398 1820 13404
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1412 12306 1440 13126
rect 1872 12306 1900 13126
rect 1964 12442 1992 13806
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1412 11665 1440 12242
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 10713 1440 11494
rect 1674 11248 1730 11257
rect 1492 11212 1544 11218
rect 1674 11183 1676 11192
rect 1492 11154 1544 11160
rect 1728 11183 1730 11192
rect 1676 11154 1728 11160
rect 1504 11121 1532 11154
rect 1490 11112 1546 11121
rect 1490 11047 1546 11056
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1412 10606 1440 10639
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1504 10169 1532 10950
rect 2056 10266 2084 13806
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2148 11762 2176 12378
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2240 10266 2268 14418
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 14006 2360 14350
rect 2792 14074 2820 14826
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2884 13870 2912 14214
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2332 11898 2360 13330
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 1490 10160 1546 10169
rect 1490 10095 1492 10104
rect 1544 10095 1546 10104
rect 1676 10124 1728 10130
rect 1492 10066 1544 10072
rect 1676 10066 1728 10072
rect 1504 10035 1532 10066
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9518 1624 9687
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1412 9217 1440 9454
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1596 9110 1624 9318
rect 1688 9178 1716 10066
rect 2240 9586 2360 9602
rect 2240 9580 2372 9586
rect 2240 9574 2320 9580
rect 1952 9512 2004 9518
rect 2240 9500 2268 9574
rect 2320 9522 2372 9528
rect 2004 9472 2268 9500
rect 1952 9454 2004 9460
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1412 8809 1440 8978
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 7857 1440 8366
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1398 7848 1454 7857
rect 1398 7783 1454 7792
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1412 7342 1440 7375
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1320 5953 1348 6734
rect 1412 6361 1440 7278
rect 1504 6866 1532 8298
rect 1964 8265 1992 9454
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1950 8256 2006 8265
rect 1950 8191 2006 8200
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1596 7546 1624 8026
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1676 7336 1728 7342
rect 1952 7336 2004 7342
rect 1676 7278 1728 7284
rect 1950 7304 1952 7313
rect 2004 7304 2006 7313
rect 1688 7002 1716 7278
rect 1950 7239 2006 7248
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1950 7168 2006 7177
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1688 6905 1716 6938
rect 1872 6905 1900 7142
rect 1950 7103 2006 7112
rect 1674 6896 1730 6905
rect 1492 6860 1544 6866
rect 1674 6831 1730 6840
rect 1858 6896 1914 6905
rect 1858 6831 1914 6840
rect 1492 6802 1544 6808
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1306 5944 1362 5953
rect 1306 5879 1362 5888
rect 1412 5778 1440 6054
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1032 4752 1084 4758
rect 1032 4694 1084 4700
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 1044 2553 1072 4694
rect 1216 4072 1268 4078
rect 1412 4049 1440 5714
rect 1504 5409 1532 6802
rect 1582 6760 1638 6769
rect 1582 6695 1584 6704
rect 1636 6695 1638 6704
rect 1584 6666 1636 6672
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1688 5545 1716 6190
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1780 5914 1808 6122
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1872 5760 1900 6190
rect 1780 5732 1900 5760
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 1490 5400 1546 5409
rect 1490 5335 1546 5344
rect 1780 5166 1808 5732
rect 1860 5296 1912 5302
rect 1964 5284 1992 7103
rect 2056 6662 2084 8978
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8022 2176 8910
rect 2136 8016 2188 8022
rect 2136 7958 2188 7964
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 1912 5256 1992 5284
rect 1860 5238 1912 5244
rect 2148 5166 2176 7958
rect 2424 7290 2452 13806
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12986 2544 13262
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2516 10538 2544 12922
rect 2700 12714 2728 13194
rect 2884 13161 2912 13806
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12442 2728 12650
rect 2884 12617 2912 12718
rect 2870 12608 2926 12617
rect 2870 12543 2926 12552
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2700 11762 2728 12242
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2700 11082 2728 11698
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2700 10266 2728 11018
rect 2976 10742 3004 16594
rect 3804 16522 3832 17002
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16046 3464 16390
rect 3804 16046 3832 16458
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 3068 14414 3096 14826
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3054 12744 3110 12753
rect 3054 12679 3110 12688
rect 3068 12646 3096 12679
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3160 12434 3188 14554
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 13870 3556 14214
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3068 12406 3188 12434
rect 3068 12102 3096 12406
rect 3146 12200 3202 12209
rect 3146 12135 3202 12144
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3160 11257 3188 12135
rect 3252 11898 3280 13330
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12986 3372 13262
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12238 3464 12786
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3620 11626 3648 15574
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 3712 14618 3740 15030
rect 3804 14958 3832 15982
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3712 13870 3740 14418
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11354 3280 11494
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3146 11248 3202 11257
rect 3146 11183 3202 11192
rect 3160 11150 3188 11183
rect 3620 11150 3648 11562
rect 3148 11144 3200 11150
rect 3608 11144 3660 11150
rect 3148 11086 3200 11092
rect 3436 11104 3608 11132
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2870 9480 2926 9489
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2608 8294 2636 8910
rect 2700 8430 2728 9454
rect 2870 9415 2926 9424
rect 2884 9382 2912 9415
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2608 8022 2636 8230
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2332 7262 2452 7290
rect 2228 7200 2280 7206
rect 2226 7168 2228 7177
rect 2280 7168 2282 7177
rect 2226 7103 2282 7112
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1216 4014 1268 4020
rect 1398 4040 1454 4049
rect 1030 2544 1086 2553
rect 1030 2479 1086 2488
rect 1124 2508 1176 2514
rect 1124 2450 1176 2456
rect 664 1828 716 1834
rect 664 1770 716 1776
rect 676 800 704 1770
rect 1136 800 1164 2450
rect 1228 1601 1256 4014
rect 1398 3975 1454 3984
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1320 2854 1348 3538
rect 1504 3505 1532 5102
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1688 4758 1716 4791
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1582 4584 1638 4593
rect 1582 4519 1638 4528
rect 1596 4078 1624 4519
rect 1780 4146 1808 5102
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 2136 4684 2188 4690
rect 1872 4622 1900 4655
rect 2136 4626 2188 4632
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 2044 4004 2096 4010
rect 1964 3964 2044 3992
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1964 3398 1992 3964
rect 2044 3946 2096 3952
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1214 1592 1270 1601
rect 1214 1527 1270 1536
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1504 241 1532 2926
rect 1596 800 1624 3130
rect 1688 2689 1716 3334
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1674 2680 1730 2689
rect 1674 2615 1730 2624
rect 1688 2446 1716 2615
rect 1964 2582 1992 2790
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2056 800 2084 3334
rect 2148 2378 2176 4626
rect 2332 4554 2360 7262
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 7002 2452 7142
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2608 6798 2636 7958
rect 2884 7954 2912 8298
rect 2976 7954 3004 9318
rect 3160 8430 3188 10406
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 7313 2820 7346
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2884 6866 2912 7686
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2424 3058 2452 5782
rect 2976 4729 3004 7890
rect 3160 7886 3188 8366
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3160 7410 3188 7822
rect 3252 7546 3280 8910
rect 3344 8537 3372 10950
rect 3330 8528 3386 8537
rect 3330 8463 3386 8472
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3344 7342 3372 8230
rect 3436 7834 3464 11104
rect 3608 11086 3660 11092
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3514 10024 3570 10033
rect 3514 9959 3570 9968
rect 3528 9382 3556 9959
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8634 3556 8978
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3436 7806 3556 7834
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6186 3188 6734
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3160 5710 3188 5850
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3160 5234 3188 5646
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3146 5128 3202 5137
rect 3146 5063 3202 5072
rect 3160 4826 3188 5063
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2516 4321 2544 4558
rect 2608 4434 2636 4558
rect 3068 4457 3096 4626
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3054 4448 3110 4457
rect 2608 4406 2820 4434
rect 2502 4312 2558 4321
rect 2792 4298 2820 4406
rect 3054 4383 3110 4392
rect 3160 4298 3188 4490
rect 2502 4247 2558 4256
rect 2688 4276 2740 4282
rect 2792 4270 2904 4298
rect 2688 4218 2740 4224
rect 2502 4176 2558 4185
rect 2502 4111 2558 4120
rect 2516 3738 2544 4111
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2608 3641 2636 3878
rect 2594 3632 2650 3641
rect 2504 3596 2556 3602
rect 2594 3567 2650 3576
rect 2504 3538 2556 3544
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2320 2984 2372 2990
rect 2318 2952 2320 2961
rect 2372 2952 2374 2961
rect 2318 2887 2374 2896
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2424 2553 2452 2790
rect 2410 2544 2466 2553
rect 2410 2479 2466 2488
rect 2136 2372 2188 2378
rect 2136 2314 2188 2320
rect 2516 800 2544 3538
rect 2700 3194 2728 4218
rect 2876 4214 2904 4270
rect 3068 4270 3188 4298
rect 2872 4208 2924 4214
rect 3068 4162 3096 4270
rect 2872 4150 2924 4156
rect 2976 4134 3096 4162
rect 2976 3890 3004 4134
rect 3056 4072 3108 4078
rect 3054 4040 3056 4049
rect 3148 4072 3200 4078
rect 3108 4040 3110 4049
rect 3148 4014 3200 4020
rect 3054 3975 3110 3984
rect 2884 3862 3004 3890
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2792 3058 2820 3606
rect 2884 3398 2912 3862
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2428 2820 2994
rect 2872 2440 2924 2446
rect 2792 2400 2872 2428
rect 2872 2382 2924 2388
rect 2976 800 3004 3674
rect 3068 3670 3096 3878
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3160 3602 3188 4014
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3252 3398 3280 7142
rect 3436 6934 3464 7686
rect 3528 7274 3556 7806
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3344 6662 3372 6802
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3344 5234 3372 6394
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3436 5545 3464 5714
rect 3422 5536 3478 5545
rect 3422 5471 3478 5480
rect 3422 5264 3478 5273
rect 3332 5228 3384 5234
rect 3422 5199 3478 5208
rect 3332 5170 3384 5176
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3344 3942 3372 4966
rect 3436 4826 3464 5199
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 4282 3464 4422
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3436 4078 3464 4218
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3528 4026 3556 7210
rect 3620 6458 3648 10066
rect 3712 9722 3740 10134
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3804 9654 3832 14758
rect 3896 12782 3924 20198
rect 3976 18692 4028 18698
rect 3976 18634 4028 18640
rect 3988 18426 4016 18634
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3988 17134 4016 18362
rect 4172 17882 4200 20198
rect 5184 19990 5212 20538
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5276 19922 5304 22200
rect 5736 20398 5764 22200
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5356 20324 5408 20330
rect 5408 20284 5488 20312
rect 5356 20266 5408 20272
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4264 19310 4292 19722
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4264 18290 4292 18838
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4356 18426 4384 18702
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4816 18290 4844 19654
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4908 18086 4936 19858
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4620 18080 4672 18086
rect 4712 18080 4764 18086
rect 4620 18022 4672 18028
rect 4710 18048 4712 18057
rect 4896 18080 4948 18086
rect 4764 18048 4766 18057
rect 4632 17882 4660 18022
rect 4896 18022 4948 18028
rect 4710 17983 4766 17992
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4724 17762 4752 17983
rect 5000 17898 5028 18770
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 18290 5120 18566
rect 5184 18306 5212 18702
rect 5276 18426 5304 19858
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5368 19514 5396 19722
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5368 18340 5396 18634
rect 5460 18442 5488 20284
rect 5552 18970 5580 20334
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5460 18414 5580 18442
rect 5736 18426 5764 20334
rect 5828 19718 5856 20402
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5828 18902 5856 19654
rect 5920 19378 5948 20198
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5448 18352 5500 18358
rect 5368 18312 5448 18340
rect 5184 18290 5304 18306
rect 5448 18294 5500 18300
rect 5080 18284 5132 18290
rect 5184 18284 5316 18290
rect 5184 18278 5264 18284
rect 5080 18226 5132 18232
rect 5264 18226 5316 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 4908 17882 5028 17898
rect 4896 17876 5028 17882
rect 4948 17870 5028 17876
rect 4896 17818 4948 17824
rect 4252 17740 4304 17746
rect 4724 17734 4936 17762
rect 4252 17682 4304 17688
rect 4264 17542 4292 17682
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4356 17338 4384 17546
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17338 4844 17614
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4172 15570 4200 15982
rect 4356 15706 4384 16594
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14550 4108 14758
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4080 13938 4108 14486
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13938 4292 14214
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4264 13530 4292 13874
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4816 12986 4844 15642
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11694 3924 12038
rect 3988 11830 4016 12310
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4080 11762 4108 12786
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3884 11688 3936 11694
rect 3936 11636 4108 11642
rect 3884 11630 4108 11636
rect 3896 11614 4108 11630
rect 3896 11565 3924 11614
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11076 3936 11082
rect 3988 11064 4016 11494
rect 3936 11036 4016 11064
rect 3884 11018 3936 11024
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3896 9178 3924 11018
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10062 4016 10542
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3988 8974 4016 9998
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3712 8362 3740 8774
rect 3988 8430 4016 8910
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 4080 8022 4108 11614
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10282 4200 10406
rect 4264 10305 4292 12310
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4528 11552 4580 11558
rect 4526 11520 4528 11529
rect 4580 11520 4582 11529
rect 4526 11455 4582 11464
rect 4632 11218 4660 11562
rect 4908 11354 4936 17734
rect 5184 15638 5212 18022
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5276 16250 5304 16594
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 5000 10810 5028 11086
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4141 10254 4200 10282
rect 4250 10296 4306 10305
rect 4141 9976 4169 10254
rect 4250 10231 4252 10240
rect 4304 10231 4306 10240
rect 4252 10202 4304 10208
rect 4264 10171 4292 10202
rect 4141 9948 4301 9976
rect 4158 9688 4214 9697
rect 4273 9674 4301 9948
rect 4158 9623 4214 9632
rect 4264 9646 4301 9674
rect 4172 9586 4200 9623
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4264 9518 4292 9646
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4356 8922 4384 10542
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10266 4660 10406
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4908 10198 4936 10610
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 5000 9874 5028 10746
rect 5092 9976 5120 13670
rect 5184 10554 5212 13670
rect 5368 12434 5396 17614
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 16794 5488 17478
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5276 12406 5396 12434
rect 5276 11694 5304 12406
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 10810 5304 11494
rect 5368 11082 5396 12174
rect 5460 11642 5488 16730
rect 5552 15706 5580 18414
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6012 18057 6040 18158
rect 5998 18048 6054 18057
rect 5998 17983 6054 17992
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15162 5580 15370
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13462 5580 14214
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5644 13190 5672 13330
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5644 12442 5672 13126
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5460 11614 5672 11642
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11354 5488 11494
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5368 10674 5396 11018
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5448 10600 5500 10606
rect 5184 10526 5396 10554
rect 5448 10542 5500 10548
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5092 9948 5192 9976
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4908 9654 4936 9862
rect 5000 9846 5120 9874
rect 5092 9704 5120 9846
rect 5164 9738 5192 9948
rect 5164 9710 5212 9738
rect 5000 9676 5120 9704
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4264 8894 4384 8922
rect 4264 8838 4292 8894
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4342 8528 4398 8537
rect 4342 8463 4398 8472
rect 4436 8492 4488 8498
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3896 7449 3924 7482
rect 3882 7440 3938 7449
rect 3882 7375 3938 7384
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 5234 3648 6054
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3712 5166 3740 6598
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5914 3832 6054
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3804 4706 3832 5510
rect 3712 4690 3832 4706
rect 3896 4690 3924 7278
rect 4080 5114 4108 7958
rect 4264 7750 4292 8230
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7449 4292 7686
rect 4250 7440 4306 7449
rect 4250 7375 4306 7384
rect 4356 7206 4384 8463
rect 4436 8434 4488 8440
rect 4448 7818 4476 8434
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4724 6644 4752 7414
rect 4816 7177 4844 9522
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4908 8634 4936 8978
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 8498 4936 8570
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4802 7168 4858 7177
rect 4802 7103 4858 7112
rect 4816 6866 4844 7103
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4804 6656 4856 6662
rect 4724 6616 4804 6644
rect 4804 6598 4856 6604
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4710 6352 4766 6361
rect 4172 5370 4200 6326
rect 4710 6287 4712 6296
rect 4764 6287 4766 6296
rect 4712 6258 4764 6264
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4264 5642 4292 5850
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3976 5092 4028 5098
rect 4080 5086 4200 5114
rect 3976 5034 4028 5040
rect 3988 4690 4016 5034
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3700 4684 3832 4690
rect 3752 4678 3832 4684
rect 3884 4684 3936 4690
rect 3700 4626 3752 4632
rect 3884 4626 3936 4632
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3712 4078 3740 4422
rect 3804 4078 3832 4558
rect 3988 4434 4016 4626
rect 3896 4406 4016 4434
rect 3700 4072 3752 4078
rect 3528 3998 3648 4026
rect 3700 4014 3752 4020
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 3720 3556 3878
rect 3436 3692 3556 3720
rect 3330 3632 3386 3641
rect 3330 3567 3332 3576
rect 3384 3567 3386 3576
rect 3332 3538 3384 3544
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3252 2564 3280 3334
rect 3344 3233 3372 3538
rect 3330 3224 3386 3233
rect 3330 3159 3386 3168
rect 3332 2576 3384 2582
rect 3252 2536 3332 2564
rect 3332 2518 3384 2524
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3160 2106 3188 2450
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 1490 232 1546 241
rect 1490 167 1546 176
rect 1582 0 1638 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3160 649 3188 2042
rect 3436 800 3464 3692
rect 3514 3360 3570 3369
rect 3514 3295 3570 3304
rect 3528 2650 3556 3295
rect 3620 2961 3648 3998
rect 3804 3738 3832 4014
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3712 3210 3740 3606
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3804 3369 3832 3402
rect 3790 3360 3846 3369
rect 3790 3295 3846 3304
rect 3712 3182 3832 3210
rect 3804 3058 3832 3182
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3606 2952 3662 2961
rect 3790 2952 3846 2961
rect 3606 2887 3662 2896
rect 3712 2910 3790 2938
rect 3620 2650 3648 2887
rect 3712 2854 3740 2910
rect 3790 2887 3846 2896
rect 3700 2848 3752 2854
rect 3792 2848 3844 2854
rect 3700 2790 3752 2796
rect 3790 2816 3792 2825
rect 3844 2816 3846 2825
rect 3790 2751 3846 2760
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3700 2576 3752 2582
rect 3698 2544 3700 2553
rect 3752 2544 3754 2553
rect 3698 2479 3754 2488
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3804 2038 3832 2450
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3804 1193 3832 1974
rect 3790 1184 3846 1193
rect 3790 1119 3846 1128
rect 3896 800 3924 4406
rect 4080 4078 4108 4966
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4172 3754 4200 5086
rect 4356 4486 4384 5782
rect 4540 5710 4568 6190
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4690 4568 5170
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4250 4312 4306 4321
rect 4356 4282 4384 4422
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4250 4247 4306 4256
rect 4344 4276 4396 4282
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3726 4200 3754
rect 3988 3126 4016 3674
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 4080 2650 4108 3726
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4172 2530 4200 3130
rect 4264 3126 4292 4247
rect 4344 4218 4396 4224
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4526 3904 4582 3913
rect 4526 3839 4582 3848
rect 4540 3602 4568 3839
rect 4632 3670 4660 4082
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4724 3670 4752 3946
rect 4816 3738 4844 6598
rect 4908 6118 4936 8230
rect 5000 6934 5028 9676
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5092 8498 5120 9114
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 7478 5120 8434
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5000 6322 5028 6734
rect 5092 6322 5120 6938
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4908 3602 4936 6054
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5000 5234 5028 5714
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 5000 4457 5028 4655
rect 4986 4448 5042 4457
rect 4986 4383 5042 4392
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4528 3596 4580 3602
rect 4896 3596 4948 3602
rect 4528 3538 4580 3544
rect 4816 3556 4896 3584
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4618 2952 4674 2961
rect 4618 2887 4674 2896
rect 4632 2854 4660 2887
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4264 2650 4292 2790
rect 4632 2650 4660 2790
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4172 2514 4292 2530
rect 4068 2508 4120 2514
rect 4172 2508 4304 2514
rect 4172 2502 4252 2508
rect 4068 2450 4120 2456
rect 4252 2450 4304 2456
rect 4080 2145 4108 2450
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4066 2136 4122 2145
rect 4066 2071 4122 2080
rect 4080 1970 4108 2071
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4172 1766 4200 2246
rect 4264 1834 4292 2450
rect 4816 2446 4844 3556
rect 4896 3538 4948 3544
rect 5000 3369 5028 3878
rect 4986 3360 5042 3369
rect 4986 3295 5042 3304
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4894 2952 4950 2961
rect 4894 2887 4950 2896
rect 4908 2650 4936 2887
rect 5000 2689 5028 2994
rect 4986 2680 5042 2689
rect 4896 2644 4948 2650
rect 4986 2615 5042 2624
rect 4896 2586 4948 2592
rect 5092 2514 5120 3878
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 5092 1850 5120 2450
rect 5184 1902 5212 9710
rect 5276 9586 5304 10406
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 8294 5304 9318
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5276 7002 5304 7958
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5276 2650 5304 6122
rect 5368 5370 5396 10526
rect 5460 5914 5488 10542
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8634 5580 9318
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5540 7200 5592 7206
rect 5538 7168 5540 7177
rect 5644 7188 5672 11614
rect 5736 10033 5764 15846
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14618 6040 14758
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6012 13530 6040 13806
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10130 5856 11086
rect 5920 10674 5948 11154
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9178 5764 9522
rect 5828 9382 5856 10066
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9518 5948 9862
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5828 8974 5856 9318
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5828 7954 5856 8910
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5920 7818 5948 8230
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5828 7546 5856 7754
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5592 7168 5672 7188
rect 5594 7160 5672 7168
rect 5538 7103 5594 7112
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4252 1828 4304 1834
rect 4252 1770 4304 1776
rect 4908 1822 5120 1850
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 4344 1692 4396 1698
rect 4344 1634 4396 1640
rect 4356 800 4384 1634
rect 4908 800 4936 1822
rect 5368 800 5396 4762
rect 5460 3641 5488 5306
rect 5446 3632 5502 3641
rect 5446 3567 5502 3576
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5460 2514 5488 2858
rect 5552 2854 5580 5782
rect 5644 5001 5672 6870
rect 5736 6866 5764 7346
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5722 6352 5778 6361
rect 5722 6287 5778 6296
rect 5736 6254 5764 6287
rect 6012 6254 6040 13194
rect 6104 11694 6132 20402
rect 6196 20380 6224 22200
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 6656 20482 6684 22200
rect 6276 20392 6328 20398
rect 6196 20352 6276 20380
rect 6196 18426 6224 20352
rect 6276 20334 6328 20340
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6196 9674 6224 15302
rect 6288 12434 6316 20198
rect 6472 20058 6500 20470
rect 6656 20454 6960 20482
rect 6932 20398 6960 20454
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6460 20052 6512 20058
rect 6460 19994 6512 20000
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6460 19848 6512 19854
rect 6380 19808 6460 19836
rect 6380 18834 6408 19808
rect 6460 19790 6512 19796
rect 6460 19168 6512 19174
rect 6564 19122 6592 19858
rect 6932 19310 6960 20198
rect 7116 19922 7144 22200
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6512 19116 6592 19122
rect 6460 19110 6592 19116
rect 6472 19094 6592 19110
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6380 17066 6408 18770
rect 6472 18086 6500 18838
rect 6564 18766 6592 19094
rect 7024 18970 7052 19722
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6642 18864 6698 18873
rect 6642 18799 6698 18808
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6656 18698 6684 18799
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6368 17060 6420 17066
rect 6368 17002 6420 17008
rect 6380 16250 6408 17002
rect 6472 16590 6500 18022
rect 6564 17678 6592 18566
rect 7116 18426 7144 19858
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6380 15570 6408 16186
rect 6472 15910 6500 16526
rect 6840 16250 6868 16662
rect 7024 16658 7052 17546
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7116 16522 7144 17002
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6380 14958 6408 15506
rect 6828 15156 6880 15162
rect 6932 15144 6960 15574
rect 6880 15116 6960 15144
rect 6828 15098 6880 15104
rect 6840 15026 6868 15098
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 7024 14226 7052 15982
rect 7208 14362 7236 20538
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7300 19378 7328 20198
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7392 18970 7420 20198
rect 7484 19922 7512 20402
rect 7576 20380 7604 22200
rect 7656 20392 7708 20398
rect 7576 20352 7656 20380
rect 7656 20334 7708 20340
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19514 7512 19858
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7668 18970 7696 20198
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7300 18086 7328 18770
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 15348 7328 18022
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 16794 7420 17682
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 17338 7512 17614
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7380 15360 7432 15366
rect 7300 15320 7380 15348
rect 7380 15302 7432 15308
rect 7576 15162 7604 18362
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 7668 16794 7696 17750
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7484 14414 7512 14826
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 14408 7524 14414
rect 7208 14334 7420 14362
rect 7472 14350 7524 14356
rect 7288 14272 7340 14278
rect 7024 14220 7288 14226
rect 7024 14214 7340 14220
rect 7024 14198 7328 14214
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6380 13258 6408 13738
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6472 12850 6500 13398
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 13258 6868 13330
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6748 12434 6776 12650
rect 6288 12406 6408 12434
rect 6748 12406 6868 12434
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6104 9646 6224 9674
rect 6104 7750 6132 9646
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 8634 6224 9454
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6196 8022 6224 8434
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 6322 6132 7686
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5736 5778 5764 6190
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5914 6040 6054
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5724 5024 5776 5030
rect 5630 4992 5686 5001
rect 5724 4966 5776 4972
rect 5630 4927 5686 4936
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5644 4282 5672 4626
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5644 3058 5672 3402
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5460 1766 5488 2450
rect 5644 2446 5672 2994
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5736 2106 5764 4966
rect 5828 4282 5856 5034
rect 5920 4622 5948 5578
rect 6104 5574 6132 6258
rect 6196 6118 6224 7958
rect 6288 7886 6316 11630
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6288 5953 6316 7822
rect 6380 6934 6408 12406
rect 6840 12238 6868 12406
rect 6932 12374 6960 13398
rect 7024 13394 7052 14198
rect 7392 14090 7420 14334
rect 7300 14062 7420 14090
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7116 12442 7144 13806
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 12102 6868 12174
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11762 6868 12038
rect 6932 11762 6960 12310
rect 7208 11898 7236 13670
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10674 6868 11154
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 9489 6500 10066
rect 6564 10062 6592 10610
rect 6932 10606 6960 11494
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7024 10538 7052 11766
rect 7012 10532 7064 10538
rect 7064 10492 7144 10520
rect 7012 10474 7064 10480
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6458 9480 6514 9489
rect 6458 9415 6514 9424
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6472 7410 6500 9415
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6564 7342 6592 7686
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6656 5846 6684 9415
rect 6748 8786 6776 9930
rect 6840 9654 6868 10134
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6748 8758 6868 8786
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6748 6254 6776 8570
rect 6840 7206 6868 8758
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6458 6868 7142
rect 6932 6798 6960 7278
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6748 5574 6776 6054
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6840 5522 6868 6122
rect 6932 6118 6960 6734
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6656 5250 6684 5510
rect 6840 5494 6960 5522
rect 6184 5228 6236 5234
rect 6656 5222 6776 5250
rect 6184 5170 6236 5176
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6012 4570 6040 5102
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4865 6132 4966
rect 6090 4856 6146 4865
rect 6090 4791 6146 4800
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5920 4078 5948 4558
rect 6012 4542 6132 4570
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5908 4072 5960 4078
rect 5828 4032 5908 4060
rect 5828 3913 5856 4032
rect 5908 4014 5960 4020
rect 5908 3936 5960 3942
rect 5814 3904 5870 3913
rect 5908 3878 5960 3884
rect 5814 3839 5870 3848
rect 5814 3768 5870 3777
rect 5814 3703 5816 3712
rect 5868 3703 5870 3712
rect 5816 3674 5868 3680
rect 5814 3224 5870 3233
rect 5814 3159 5870 3168
rect 5828 2582 5856 3159
rect 5920 2650 5948 3878
rect 6012 2990 6040 4150
rect 6104 3126 6132 4542
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6196 2774 6224 5170
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6288 4214 6316 4422
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6288 3194 6316 3946
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6196 2746 6316 2774
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 6288 2514 6316 2746
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5816 1828 5868 1834
rect 5816 1770 5868 1776
rect 5448 1760 5500 1766
rect 5448 1702 5500 1708
rect 5828 800 5856 1770
rect 6288 800 6316 2450
rect 6380 2038 6408 5034
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6472 4593 6500 4626
rect 6458 4584 6514 4593
rect 6458 4519 6514 4528
rect 6460 4480 6512 4486
rect 6552 4480 6604 4486
rect 6460 4422 6512 4428
rect 6550 4448 6552 4457
rect 6604 4448 6606 4457
rect 6472 2514 6500 4422
rect 6550 4383 6606 4392
rect 6564 3602 6592 4383
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2650 6592 2790
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6368 2032 6420 2038
rect 6368 1974 6420 1980
rect 6472 1834 6500 2450
rect 6656 1970 6684 5102
rect 6748 4162 6776 5222
rect 6932 4706 6960 5494
rect 7024 4826 7052 8298
rect 7116 8022 7144 10492
rect 7300 8362 7328 14062
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7484 13326 7512 13942
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12442 7420 13126
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7484 12306 7512 13262
rect 7576 12434 7604 14418
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7668 12986 7696 13874
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7576 12406 7696 12434
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7392 11529 7420 11834
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7378 11520 7434 11529
rect 7378 11455 7434 11464
rect 7576 11082 7604 11562
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 10674 7604 11018
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7668 10554 7696 12406
rect 7576 10526 7696 10554
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 8906 7512 9386
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6932 4678 7052 4706
rect 7024 4622 7052 4678
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6840 4264 6868 4558
rect 6840 4236 6960 4264
rect 6932 4162 6960 4236
rect 6748 4134 6868 4162
rect 6932 4146 7052 4162
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6840 4026 6868 4134
rect 6920 4140 7052 4146
rect 6972 4134 7052 4140
rect 6920 4082 6972 4088
rect 6748 3534 6776 4014
rect 6840 3998 6960 4026
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3777 6868 3878
rect 6826 3768 6882 3777
rect 6932 3738 6960 3998
rect 6826 3703 6882 3712
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6736 3528 6788 3534
rect 6932 3505 6960 3674
rect 6736 3470 6788 3476
rect 6918 3496 6974 3505
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 6460 1828 6512 1834
rect 6460 1770 6512 1776
rect 6748 800 6776 3470
rect 6828 3460 6880 3466
rect 6918 3431 6974 3440
rect 6828 3402 6880 3408
rect 6840 2774 6868 3402
rect 6920 3052 6972 3058
rect 7024 3040 7052 4134
rect 6972 3012 7052 3040
rect 6920 2994 6972 3000
rect 6840 2746 6960 2774
rect 6826 2680 6882 2689
rect 6826 2615 6882 2624
rect 6840 2582 6868 2615
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6932 2394 6960 2746
rect 7116 2514 7144 7686
rect 7208 7478 7236 7822
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7208 7002 7236 7414
rect 7300 7410 7328 7890
rect 7392 7546 7420 7890
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7208 6322 7236 6938
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 6322 7512 6802
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7208 5914 7236 6258
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7300 5914 7328 6122
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7208 5234 7236 5850
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7194 5128 7250 5137
rect 7194 5063 7196 5072
rect 7248 5063 7250 5072
rect 7196 5034 7248 5040
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 6840 2366 6960 2394
rect 6840 2310 6868 2366
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 2106 7144 2246
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7208 800 7236 4626
rect 7300 4554 7328 4966
rect 7392 4826 7420 6054
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7484 5302 7512 5782
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7300 3942 7328 4490
rect 7392 4185 7420 4626
rect 7484 4554 7512 5238
rect 7576 4706 7604 10526
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10266 7696 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7760 10146 7788 20266
rect 8036 20244 8064 22200
rect 8496 20398 8524 22200
rect 8956 20398 8984 22200
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8036 20216 8340 20244
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8312 19990 8340 20216
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8312 18902 8340 19926
rect 8404 18970 8432 20334
rect 8496 20058 8524 20334
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8496 19378 8524 19654
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8588 19258 8616 20198
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8680 19378 8708 19654
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8496 19230 8616 19258
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8496 16232 8524 19230
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8588 18154 8616 19110
rect 8680 18766 8708 19314
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 16794 8708 17614
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8404 16204 8524 16232
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 14958 8248 15302
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8312 14550 8340 14758
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8404 13870 8432 16204
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8496 15706 8524 16050
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 12782 7880 13330
rect 8484 13320 8536 13326
rect 8588 13308 8616 13738
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8536 13280 8616 13308
rect 8484 13262 8536 13268
rect 7840 12776 7892 12782
rect 7892 12736 8248 12764
rect 7840 12718 7892 12724
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12306 8248 12736
rect 8680 12442 8708 13466
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8404 11150 8432 11494
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8392 11144 8444 11150
rect 8444 11104 8524 11132
rect 8392 11086 8444 11092
rect 8496 10606 8524 11104
rect 8588 10810 8616 11154
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7668 10118 7788 10146
rect 7668 8566 7696 10118
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9178 7788 9998
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8312 9178 8340 9522
rect 8404 9518 8432 10542
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8392 8968 8444 8974
rect 8496 8956 8524 9590
rect 8680 8974 8708 12106
rect 8772 9110 8800 19722
rect 8956 18834 8984 19994
rect 9140 19922 9168 20402
rect 9416 20398 9444 22200
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9876 20330 9904 22200
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9034 19816 9090 19825
rect 9034 19751 9090 19760
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8864 17882 8892 18022
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 9048 15706 9076 19751
rect 9140 19514 9168 19858
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9232 19310 9260 20198
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9324 18970 9352 20266
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9416 19378 9444 20198
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18426 9260 18770
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9402 18320 9458 18329
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9312 18284 9364 18290
rect 9402 18255 9458 18264
rect 9312 18226 9364 18232
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 13530 9076 15642
rect 9140 14958 9168 18226
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17882 9260 18022
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9324 17270 9352 18226
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9416 14634 9444 18255
rect 9508 15706 9536 19382
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9324 14606 9444 14634
rect 9220 14408 9272 14414
rect 9324 14396 9352 14606
rect 9508 14498 9536 15642
rect 9692 14958 9720 18294
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9588 14884 9640 14890
rect 9588 14826 9640 14832
rect 9272 14368 9352 14396
rect 9220 14350 9272 14356
rect 9324 13938 9352 14368
rect 9416 14470 9536 14498
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9218 13832 9274 13841
rect 9218 13767 9220 13776
rect 9272 13767 9274 13776
rect 9220 13738 9272 13744
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9324 13462 9352 13670
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9416 13394 9444 14470
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9508 13462 9536 14282
rect 9600 13734 9628 14826
rect 9692 14482 9720 14894
rect 9784 14618 9812 20198
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18766 9996 19178
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9954 18184 10010 18193
rect 9954 18119 10010 18128
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9876 17746 9904 17818
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9876 17338 9904 17682
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9784 14278 9812 14554
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9678 14002 9734 14011
rect 9678 13937 9734 13946
rect 9876 13852 9904 16186
rect 9968 15706 9996 18119
rect 10152 15706 10180 20538
rect 10336 20398 10364 22200
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10244 19514 10272 20334
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10336 18970 10364 20334
rect 10612 20330 10640 20538
rect 10796 20482 10824 22200
rect 10796 20466 11100 20482
rect 10796 20460 11112 20466
rect 10796 20454 11060 20460
rect 11060 20402 11112 20408
rect 11256 20398 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11716 20330 11744 22200
rect 11796 20528 11848 20534
rect 12176 20516 12204 22200
rect 12176 20488 12480 20516
rect 11796 20470 11848 20476
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10230 18728 10286 18737
rect 10230 18663 10286 18672
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9784 13824 9904 13852
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9140 12374 9168 13126
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9232 11762 9260 13330
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12170 9352 13126
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9402 12744 9458 12753
rect 9402 12679 9404 12688
rect 9456 12679 9458 12688
rect 9404 12650 9456 12656
rect 9508 12646 9536 12786
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9508 12374 9536 12582
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8444 8928 8524 8956
rect 8668 8968 8720 8974
rect 8392 8910 8444 8916
rect 8668 8910 8720 8916
rect 8128 8820 8156 8910
rect 8404 8820 8432 8910
rect 8128 8792 8432 8820
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 8206 8392 8262 8401
rect 7668 8022 7696 8366
rect 8206 8327 8208 8336
rect 8260 8327 8262 8336
rect 8208 8298 8260 8304
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 4826 7696 7686
rect 7760 6458 7788 7754
rect 8312 7274 8340 7822
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8312 7002 8340 7210
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 7930 6760 7986 6769
rect 7930 6695 7932 6704
rect 7984 6695 7986 6704
rect 7932 6666 7984 6672
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7576 4678 7696 4706
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7378 4176 7434 4185
rect 7434 4134 7512 4162
rect 7378 4111 7434 4120
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7392 3754 7420 3946
rect 7300 3726 7420 3754
rect 7300 3126 7328 3726
rect 7484 3602 7512 4134
rect 7576 3738 7604 4558
rect 7668 4321 7696 4678
rect 7654 4312 7710 4321
rect 7654 4247 7710 4256
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7392 2446 7420 3130
rect 7484 2650 7512 3334
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7668 800 7696 4082
rect 7760 3466 7788 6190
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8116 5840 8168 5846
rect 8114 5808 8116 5817
rect 8168 5808 8170 5817
rect 7932 5772 7984 5778
rect 8114 5743 8170 5752
rect 7932 5714 7984 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7852 5574 7880 5646
rect 7944 5574 7972 5714
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7852 5166 7880 5510
rect 8220 5370 8248 6054
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8404 4826 8432 8792
rect 8680 8634 8708 8910
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8680 8378 8708 8570
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8588 8350 8708 8378
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8128 4010 8156 4218
rect 8312 4146 8340 4626
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3670 8248 3878
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 8036 2922 8064 3606
rect 8312 3534 8340 3674
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 2922 8340 3470
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8404 2774 8432 4626
rect 8496 4146 8524 7482
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8496 3738 8524 4082
rect 8588 3738 8616 8350
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7818 8708 8230
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 6905 8708 7210
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8680 4078 8708 6666
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5098 8800 6054
rect 8864 5658 8892 8502
rect 8956 7954 8984 11630
rect 9140 10606 9168 11698
rect 9600 11694 9628 13670
rect 9784 12628 9812 13824
rect 9968 13546 9996 15642
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9876 13518 9996 13546
rect 9876 12782 9904 13518
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9784 12600 9904 12628
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11354 9628 11494
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9450 9168 9998
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9232 9722 9260 9862
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8430 9076 9318
rect 9140 8838 9168 9386
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8498 9168 8774
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 8864 5630 9076 5658
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8772 4622 8800 5034
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8772 4010 8800 4150
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8220 2746 8432 2774
rect 8220 898 8248 2746
rect 8496 2650 8524 3431
rect 8588 3398 8616 3538
rect 8576 3392 8628 3398
rect 8772 3369 8800 3946
rect 8576 3334 8628 3340
rect 8758 3360 8814 3369
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8128 870 8248 898
rect 8128 800 8156 870
rect 8588 800 8616 3334
rect 8758 3295 8814 3304
rect 8864 3058 8892 5102
rect 9048 5098 9076 5630
rect 9232 5137 9260 6054
rect 9218 5128 9274 5137
rect 9036 5092 9088 5098
rect 9218 5063 9274 5072
rect 9036 5034 9088 5040
rect 9048 4826 9076 5034
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 2446 8800 2858
rect 8956 2514 8984 4422
rect 9048 4282 9076 4762
rect 9232 4758 9260 5063
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9048 3738 9076 3878
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9140 2774 9168 3878
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9232 3194 9260 3470
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9232 2990 9260 3130
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9324 2774 9352 9930
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8498 9444 8910
rect 9508 8634 9536 10066
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9692 8537 9720 11562
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10062 9812 10406
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9876 8650 9904 12600
rect 9968 11150 9996 13330
rect 10060 13002 10088 14418
rect 10152 13258 10180 14486
rect 10244 14482 10272 18663
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10244 13841 10272 13874
rect 10336 13870 10364 18362
rect 10428 16250 10456 20198
rect 11072 20074 11100 20266
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 10980 20046 11100 20074
rect 10980 20040 11008 20046
rect 10888 20012 11008 20040
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 19310 10548 19790
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10520 17746 10548 19246
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10704 18766 10732 18906
rect 10796 18834 10824 19110
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10520 16590 10548 17070
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 13864 10376 13870
rect 10230 13832 10286 13841
rect 10324 13806 10376 13812
rect 10230 13767 10286 13776
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10244 13258 10272 13398
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10232 13252 10284 13258
rect 10428 13240 10456 15642
rect 10520 14618 10548 15846
rect 10612 15162 10640 15846
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10704 14770 10732 18158
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10796 16250 10824 16594
rect 10888 16454 10916 20012
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11072 18630 11100 19926
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18970 11192 19110
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11164 18290 11192 18770
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10980 17338 11008 17750
rect 11072 17542 11100 18022
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10980 16794 11008 17274
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11072 16998 11100 17070
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10612 14742 10732 14770
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10428 13212 10548 13240
rect 10232 13194 10284 13200
rect 10244 13138 10272 13194
rect 10244 13110 10456 13138
rect 10060 12974 10272 13002
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9968 9518 9996 11086
rect 10060 10266 10088 12718
rect 10244 11694 10272 12974
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10244 10198 10272 11630
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10336 10810 10364 11154
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10244 9110 10272 9998
rect 10336 9722 10364 10406
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9876 8622 9996 8650
rect 9678 8528 9734 8537
rect 9404 8492 9456 8498
rect 9678 8463 9734 8472
rect 9864 8492 9916 8498
rect 9404 8434 9456 8440
rect 9864 8434 9916 8440
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7342 9536 7890
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9600 6798 9628 8230
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 7002 9720 7346
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6866 9812 7958
rect 9876 7886 9904 8434
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 7002 9904 7142
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9968 6798 9996 8622
rect 10152 8362 10180 9046
rect 10244 8498 10272 9046
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 8498 10364 8774
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7002 10364 7822
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 9588 6792 9640 6798
rect 9956 6792 10008 6798
rect 9588 6734 9640 6740
rect 9770 6760 9826 6769
rect 9404 5296 9456 5302
rect 9600 5273 9628 6734
rect 9956 6734 10008 6740
rect 9770 6695 9772 6704
rect 9824 6695 9826 6704
rect 9772 6666 9824 6672
rect 9968 5846 9996 6734
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10244 5914 10272 6122
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9404 5238 9456 5244
rect 9586 5264 9642 5273
rect 9416 4049 9444 5238
rect 10244 5234 10272 5850
rect 9586 5199 9642 5208
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9770 4856 9826 4865
rect 9968 4826 9996 4966
rect 9770 4791 9772 4800
rect 9824 4791 9826 4800
rect 9956 4820 10008 4826
rect 9772 4762 9824 4768
rect 9956 4762 10008 4768
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9416 3505 9444 3975
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9508 3346 9536 4694
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 3528 9640 3534
rect 9692 3482 9720 4150
rect 9864 3936 9916 3942
rect 9770 3904 9826 3913
rect 9864 3878 9916 3884
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9770 3839 9826 3848
rect 9640 3476 9720 3482
rect 9588 3470 9720 3476
rect 9600 3454 9720 3470
rect 9784 3466 9812 3839
rect 9876 3738 9904 3878
rect 10060 3738 10088 3878
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10152 3602 10180 4490
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10244 3602 10272 4082
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9048 2746 9168 2774
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8956 1698 8984 2450
rect 8944 1692 8996 1698
rect 8944 1634 8996 1640
rect 9048 800 9076 2746
rect 9140 2514 9168 2746
rect 9232 2746 9352 2774
rect 9416 3318 9536 3346
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9232 2650 9260 2746
rect 9416 2650 9444 3318
rect 9600 2990 9628 3334
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9508 2446 9536 2790
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9600 800 9628 2926
rect 9692 2446 9720 3130
rect 10152 3126 10180 3538
rect 10244 3194 10272 3538
rect 10428 3194 10456 13110
rect 10520 12986 10548 13212
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10612 11082 10640 14742
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10704 14414 10732 14554
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10704 12238 10732 12786
rect 10796 12646 10824 14418
rect 10888 14226 10916 16390
rect 11072 15570 11100 16934
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 14890 11008 15438
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14958 11100 15302
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10980 14396 11008 14826
rect 11058 14648 11114 14657
rect 11164 14618 11192 17070
rect 11256 16250 11284 20198
rect 11808 20058 11836 20470
rect 12452 20398 12480 20488
rect 12348 20392 12400 20398
rect 12084 20330 12296 20346
rect 12348 20334 12400 20340
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12072 20324 12296 20330
rect 12124 20318 12296 20324
rect 12072 20266 12124 20272
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18970 11744 19110
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11808 18902 11836 19722
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17202 11744 17614
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11348 16794 11376 16934
rect 11808 16794 11836 18022
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11716 16454 11744 16662
rect 11900 16590 11928 20198
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11992 19310 12020 19654
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12084 18426 12112 19858
rect 12176 18970 12204 20198
rect 12268 18970 12296 20318
rect 12360 19854 12388 20334
rect 12452 20262 12480 20334
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12636 20058 12664 22200
rect 13096 20534 13124 22200
rect 13556 20534 13584 22200
rect 14016 20534 14044 22200
rect 14476 20534 14504 22200
rect 14936 20534 14964 22200
rect 15396 20534 15424 22200
rect 15856 20534 15884 22200
rect 16316 20534 16344 22200
rect 16776 20534 16804 22200
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14924 20528 14976 20534
rect 14924 20470 14976 20476
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 12912 20058 12940 20266
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12084 17746 12112 18226
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 17134 12020 17478
rect 12084 17338 12112 17682
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11992 16658 12020 17070
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11256 15910 11284 16186
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11440 15638 11468 16050
rect 11716 16046 11744 16118
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11440 15416 11468 15574
rect 11256 15388 11468 15416
rect 11256 15162 11284 15388
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11716 15042 11744 15982
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11256 15014 11744 15042
rect 11058 14583 11060 14592
rect 11112 14583 11114 14592
rect 11152 14612 11204 14618
rect 11060 14554 11112 14560
rect 11152 14554 11204 14560
rect 11060 14408 11112 14414
rect 10980 14368 11060 14396
rect 11060 14350 11112 14356
rect 10888 14198 11100 14226
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10980 12594 11008 14010
rect 11072 13818 11100 14198
rect 11164 13938 11192 14554
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11072 13790 11192 13818
rect 10796 12434 10824 12582
rect 10980 12566 11100 12594
rect 10796 12406 11008 12434
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 12102 10732 12174
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11762 10732 12038
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10888 11150 10916 11698
rect 10980 11626 11008 12406
rect 11072 12102 11100 12566
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10980 10470 11008 10746
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 11072 10062 11100 11698
rect 11060 10056 11112 10062
rect 10980 10016 11060 10044
rect 10980 9654 11008 10016
rect 11060 9998 11112 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10968 9648 11020 9654
rect 10888 9608 10968 9636
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 9382 10732 9522
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10520 6769 10548 9114
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10520 4826 10548 6326
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10506 4720 10562 4729
rect 10506 4655 10508 4664
rect 10560 4655 10562 4664
rect 10508 4626 10560 4632
rect 10612 4146 10640 8502
rect 10704 8022 10732 9318
rect 10888 8974 10916 9608
rect 10968 9590 11020 9596
rect 11072 9586 11100 9862
rect 11164 9674 11192 13790
rect 11256 11218 11284 15014
rect 11808 14822 11836 15506
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 15026 12020 15302
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 12084 14346 12112 16934
rect 12176 16794 12204 18022
rect 12360 17882 12388 18702
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 15162 12480 15982
rect 12544 15570 12572 16050
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12268 14414 12296 15030
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11794 13968 11850 13977
rect 11794 13903 11850 13912
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10266 11284 10610
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11164 9646 11284 9674
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10796 7546 10824 8502
rect 10980 8498 11008 8978
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11072 8294 11100 9386
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11164 8634 11192 9318
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 11072 7274 11100 7958
rect 11164 7750 11192 8230
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10704 6730 10732 6938
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10704 6254 10732 6666
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10888 6254 10916 7142
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10980 6798 11008 6938
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10704 5710 10732 6190
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 4554 10732 5646
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2922 10272 2994
rect 10324 2984 10376 2990
rect 10508 2984 10560 2990
rect 10376 2944 10508 2972
rect 10324 2926 10376 2932
rect 10508 2926 10560 2932
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10060 800 10088 2450
rect 10520 800 10548 2790
rect 10704 2530 10732 4082
rect 10796 3097 10824 5510
rect 10888 5166 10916 5850
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10980 5114 11008 5850
rect 11072 5846 11100 6870
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5710 11100 5782
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5234 11100 5646
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10980 5086 11100 5114
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10782 3088 10838 3097
rect 10782 3023 10838 3032
rect 10888 2854 10916 4626
rect 11072 4282 11100 5086
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 4706 11284 9646
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11164 4678 11284 4706
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 4185 11192 4678
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11150 4176 11206 4185
rect 10968 4140 11020 4146
rect 11150 4111 11206 4120
rect 10968 4082 11020 4088
rect 10980 2922 11008 4082
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10796 2650 10824 2790
rect 11072 2774 11100 3878
rect 11164 3516 11192 4111
rect 11164 3488 11284 3516
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10980 2746 11100 2774
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10704 2502 10824 2530
rect 10796 2446 10824 2502
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10980 2394 11008 2746
rect 11164 2582 11192 3334
rect 11256 2990 11284 3488
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 3194 11744 13806
rect 11808 13462 11836 13903
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11808 12889 11836 13398
rect 11794 12880 11850 12889
rect 11794 12815 11796 12824
rect 11848 12815 11850 12824
rect 11796 12786 11848 12792
rect 11808 12442 11836 12786
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11808 11898 11836 12242
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 11665 11836 11698
rect 11794 11656 11850 11665
rect 11794 11591 11850 11600
rect 11900 11336 11928 14214
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11992 11762 12020 12922
rect 12084 12170 12112 13330
rect 12176 12442 12204 13670
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11762 12112 12106
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11900 11308 12020 11336
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 9450 11836 10950
rect 11900 10470 11928 11154
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11794 9344 11850 9353
rect 11794 9279 11850 9288
rect 11808 8022 11836 9279
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 6934 11836 7686
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11808 5234 11836 6870
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11808 4622 11836 5170
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11900 4434 11928 10406
rect 11992 5846 12020 11308
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 9353 12112 10950
rect 12176 9489 12204 11834
rect 12162 9480 12218 9489
rect 12162 9415 12218 9424
rect 12164 9376 12216 9382
rect 12070 9344 12126 9353
rect 12164 9318 12216 9324
rect 12070 9279 12126 9288
rect 12176 9178 12204 9318
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12268 9058 12296 12922
rect 12360 11898 12388 14214
rect 12636 14074 12664 19858
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12820 19334 12848 19790
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 19378 13032 19654
rect 13280 19514 13308 20266
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 20058 13584 20198
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 12728 19306 12848 19334
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12728 18834 12756 19306
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12452 13954 12480 14010
rect 12452 13926 12664 13954
rect 12636 13734 12664 13926
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12544 11898 12572 13670
rect 12728 13546 12756 18770
rect 13648 17882 13676 20334
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 14372 20324 14424 20330
rect 14372 20266 14424 20272
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 13740 19514 13768 20266
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19718 13860 20198
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14292 19310 14320 19654
rect 14384 19514 14412 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 13740 18970 13768 19246
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17338 13400 17682
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 16130 13124 16390
rect 13188 16250 13216 17070
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13096 16102 13216 16130
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13004 15366 13032 15506
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 15026 13032 15302
rect 13096 15162 13124 15982
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13188 15094 13216 16102
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 14618 12848 14826
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12912 14074 12940 14758
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12636 13518 12756 13546
rect 12636 12050 12664 13518
rect 12820 13258 12848 13874
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12820 12782 12848 13194
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12442 12756 12582
rect 13096 12442 13124 14350
rect 13188 13938 13216 15030
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13280 14278 13308 14554
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13372 13938 13400 14350
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12636 12022 12848 12050
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12360 11014 12388 11154
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10130 12480 10406
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12084 9030 12296 9058
rect 12084 5914 12112 9030
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8566 12204 8910
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12268 8566 12296 8842
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12176 6866 12204 8502
rect 12360 7528 12388 9862
rect 12452 8838 12480 10066
rect 12544 9654 12572 11494
rect 12636 11014 12664 11562
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12268 7500 12388 7528
rect 12268 7342 12296 7500
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12268 6390 12296 6695
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12072 5908 12124 5914
rect 12124 5868 12204 5896
rect 12072 5850 12124 5856
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11992 5137 12020 5782
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11978 5128 12034 5137
rect 11978 5063 11980 5072
rect 12032 5063 12034 5072
rect 11980 5034 12032 5040
rect 11992 5003 12020 5034
rect 12084 4826 12112 5714
rect 12176 5166 12204 5868
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12268 4978 12296 6054
rect 12176 4950 12296 4978
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11808 4406 11928 4434
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11440 2774 11468 2926
rect 11348 2746 11468 2774
rect 11808 2774 11836 4406
rect 11992 3942 12020 4626
rect 12070 4584 12126 4593
rect 12070 4519 12072 4528
rect 12124 4519 12126 4528
rect 12072 4490 12124 4496
rect 11980 3936 12032 3942
rect 11978 3904 11980 3913
rect 12032 3904 12034 3913
rect 11978 3839 12034 3848
rect 12084 3738 12112 4490
rect 12176 3738 12204 4950
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12268 4282 12296 4762
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12360 4214 12388 7346
rect 12544 6798 12572 7890
rect 12532 6792 12584 6798
rect 12438 6760 12494 6769
rect 12532 6734 12584 6740
rect 12438 6695 12440 6704
rect 12492 6695 12494 6704
rect 12440 6666 12492 6672
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5778 12572 6598
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12544 4758 12572 5238
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12452 4146 12480 4490
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12346 4040 12402 4049
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11900 3618 11928 3674
rect 11900 3590 12112 3618
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 3058 11928 3470
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12084 2774 12112 3590
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 2990 12204 3334
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11808 2746 12020 2774
rect 12084 2746 12204 2774
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11348 2514 11376 2746
rect 11992 2650 12020 2746
rect 12176 2650 12204 2746
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11060 2440 11112 2446
rect 10980 2388 11060 2394
rect 10980 2382 11112 2388
rect 10980 2366 11100 2382
rect 10980 800 11008 2366
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11256 1902 11284 2246
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11440 800 11468 1974
rect 11900 800 11928 2246
rect 12268 1442 12296 4014
rect 12346 3975 12402 3984
rect 12360 3534 12388 3975
rect 12440 3596 12492 3602
rect 12544 3584 12572 4422
rect 12636 4060 12664 10474
rect 12728 9926 12756 11086
rect 12820 10538 12848 12022
rect 13188 11830 13216 13466
rect 13280 12434 13308 13670
rect 13372 12646 13400 13874
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13280 12406 13400 12434
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11014 12940 11494
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 13096 10538 13124 11154
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12912 9926 12940 10474
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9586 12940 9862
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 9042 12940 9522
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8498 12756 8842
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 8090 12756 8298
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12820 7954 12848 8434
rect 13004 8430 13032 10134
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12820 6118 12848 7890
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 6390 12940 7210
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13096 5234 13124 5782
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12728 4622 12756 5170
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 13096 4282 13124 5170
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12636 4032 12756 4060
rect 12728 3942 12756 4032
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12492 3556 12572 3584
rect 12440 3538 12492 3544
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 2514 12388 2926
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12268 1414 12388 1442
rect 12360 800 12388 1414
rect 12820 800 12848 3402
rect 12912 2514 12940 3878
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 2582 13032 3334
rect 13096 2650 13124 3538
rect 13188 2650 13216 9998
rect 13280 9110 13308 12310
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13280 8430 13308 9046
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13372 8362 13400 12406
rect 13464 10130 13492 16730
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13556 14958 13584 15642
rect 13544 14952 13596 14958
rect 13740 14906 13768 18906
rect 13832 16182 13860 19246
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13544 14894 13596 14900
rect 13648 14878 13768 14906
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 13326 13584 13670
rect 13648 13530 13676 14878
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14346 13768 14758
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13728 13728 13780 13734
rect 13832 13716 13860 14350
rect 13780 13688 13860 13716
rect 13728 13670 13780 13676
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12986 13584 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13740 12889 13768 13670
rect 13726 12880 13782 12889
rect 13726 12815 13782 12824
rect 13740 12782 13768 12815
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12238 13676 12582
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9518 13492 9862
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 9178 13584 9454
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13556 8294 13584 8910
rect 13648 8634 13676 8978
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13740 7954 13768 8774
rect 13832 8362 13860 12242
rect 13924 9654 13952 18090
rect 14016 12102 14044 18770
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14108 15706 14136 16050
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 13870 14136 14418
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 13394 14136 13806
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14108 11354 14136 12650
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10198 14136 10406
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14108 9586 14136 10134
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13924 8090 13952 8842
rect 14016 8430 14044 8910
rect 14200 8514 14228 15914
rect 14292 11694 14320 19246
rect 14568 18970 14596 19246
rect 15212 19174 15240 20266
rect 15396 19446 15424 20334
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 16212 20324 16264 20330
rect 16212 20266 16264 20272
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 15672 19514 15700 20266
rect 16224 19514 16252 20266
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16592 19718 16620 19858
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14476 16794 14504 18770
rect 14844 18154 14872 18770
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14384 14414 14412 15438
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14568 11642 14596 16594
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14660 14657 14688 14758
rect 14646 14648 14702 14657
rect 14646 14583 14702 14592
rect 14752 13938 14780 14758
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15212 14550 15240 14962
rect 15304 14618 15332 19246
rect 15580 18902 15608 19246
rect 15948 18970 15976 19246
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14660 13530 14688 13670
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 15488 13462 15516 17750
rect 15580 13530 15608 18838
rect 16132 18630 16160 19246
rect 16408 18630 16436 19246
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15026 15792 15302
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13938 15700 14214
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 12714 14688 13262
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14660 12442 14688 12650
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15304 12442 15332 13126
rect 15672 12850 15700 13874
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 12986 15884 13330
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14660 11762 14688 12378
rect 15672 12306 15700 12786
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14738 11656 14794 11665
rect 14568 11614 14688 11642
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14108 8486 14228 8514
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13924 7410 13952 8026
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 4826 13676 5034
rect 14002 4856 14058 4865
rect 13636 4820 13688 4826
rect 14002 4791 14004 4800
rect 13636 4762 13688 4768
rect 14056 4791 14058 4800
rect 14004 4762 14056 4768
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13372 4214 13400 4490
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13360 4208 13412 4214
rect 13266 4176 13322 4185
rect 13360 4150 13412 4156
rect 13266 4111 13268 4120
rect 13320 4111 13322 4120
rect 13268 4082 13320 4088
rect 14016 3670 14044 4762
rect 14108 3738 14136 8486
rect 14186 8392 14242 8401
rect 14186 8327 14188 8336
rect 14240 8327 14242 8336
rect 14188 8298 14240 8304
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6118 14320 7142
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14384 5914 14412 11222
rect 14476 10810 14504 11494
rect 14568 11354 14596 11494
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14660 10656 14688 11614
rect 14738 11591 14794 11600
rect 14752 11558 14780 11591
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14568 10628 14688 10656
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 6866 14504 10406
rect 14568 9178 14596 10628
rect 14752 10554 14780 11494
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15488 11150 15516 12242
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15028 10674 15056 11086
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14660 10526 14780 10554
rect 14660 10062 14688 10526
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14568 8430 14596 9114
rect 14752 8566 14780 10406
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7410 14596 8230
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14752 7002 14780 8502
rect 15212 8362 15240 8774
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15304 7342 15332 8842
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14108 3602 14136 3674
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14292 3466 14320 4966
rect 14384 3942 14412 5510
rect 14476 5030 14504 6122
rect 14568 5710 14596 6734
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5794 14688 6054
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14660 5778 14872 5794
rect 14660 5772 14884 5778
rect 14660 5766 14832 5772
rect 14832 5714 14884 5720
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4758 14504 4966
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14568 4690 14596 5646
rect 14752 5234 14780 5646
rect 15212 5642 15240 6190
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5846 15332 6054
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15212 5234 15240 5578
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4826 14780 4966
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14740 4820 14792 4826
rect 15212 4808 15240 5170
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15304 4826 15332 4966
rect 14740 4762 14792 4768
rect 15120 4780 15240 4808
rect 15292 4820 15344 4826
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14648 4616 14700 4622
rect 14752 4593 14780 4626
rect 14648 4558 14700 4564
rect 14738 4584 14794 4593
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13280 3058 13308 3334
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12912 2038 12940 2450
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 13280 800 13308 2314
rect 13372 2106 13400 2926
rect 13556 2514 13584 3334
rect 14292 2990 14320 3402
rect 14384 3058 14412 3878
rect 14660 3738 14688 4558
rect 14738 4519 14794 4528
rect 14936 4078 14964 4626
rect 15120 4282 15148 4780
rect 15292 4762 15344 4768
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14752 3516 14780 3946
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14924 3528 14976 3534
rect 14752 3488 14924 3516
rect 14924 3470 14976 3476
rect 14936 3194 14964 3470
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 13924 2582 13952 2790
rect 14292 2582 14320 2790
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 14280 2576 14332 2582
rect 14280 2518 14332 2524
rect 14476 2514 14504 2790
rect 14660 2650 14688 2926
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 15212 2514 15240 4422
rect 15396 3602 15424 7142
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 5846 15516 6598
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15488 4554 15516 5034
rect 15580 4758 15608 5510
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15672 3738 15700 8366
rect 15856 8022 15884 9998
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7886 15884 7958
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7410 15792 7686
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15396 3194 15424 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15396 2514 15424 2790
rect 15488 2582 15516 3062
rect 15580 2990 15608 3606
rect 15672 2990 15700 3674
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 3058 15792 3334
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15672 2582 15700 2790
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13740 800 13768 2314
rect 14292 800 14320 2314
rect 14752 800 14780 2314
rect 15212 800 15240 2314
rect 15672 800 15700 2314
rect 15948 2310 15976 12582
rect 16132 10130 16160 18566
rect 16408 17814 16436 18566
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16224 12646 16252 13398
rect 16316 12646 16344 13466
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16224 11898 16252 12242
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16316 6730 16344 12582
rect 16408 12238 16436 12650
rect 16500 12374 16528 12718
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16408 11694 16436 12174
rect 16500 11762 16528 12310
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16592 10742 16620 19654
rect 16684 19174 16712 20266
rect 17236 19990 17264 22200
rect 17696 20534 17724 22200
rect 18156 20534 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18616 20534 18644 22200
rect 19076 20534 19104 22200
rect 19536 20534 19564 22200
rect 19996 20534 20024 22200
rect 20456 20534 20484 22200
rect 20916 20534 20944 22200
rect 21376 20602 21404 22200
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20904 20528 20956 20534
rect 20904 20470 20956 20476
rect 21836 20466 21864 22200
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17880 20058 17908 20266
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17420 19514 17448 19858
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 16684 18222 16712 18770
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 17144 11082 17172 19178
rect 17972 19174 18000 20334
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 20076 20324 20128 20330
rect 20076 20266 20128 20272
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 18156 19514 18184 20266
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18800 19514 18828 20266
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18604 19304 18656 19310
rect 18892 19292 18920 20266
rect 18604 19246 18656 19252
rect 18800 19264 18920 19292
rect 19064 19304 19116 19310
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17316 18760 17368 18766
rect 18156 18714 18184 19246
rect 18340 18970 18368 19246
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 17316 18702 17368 18708
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16408 2990 16436 8298
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16500 4622 16528 5238
rect 17144 5030 17172 9046
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 5234 17264 7686
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17328 5166 17356 18702
rect 17972 18686 18184 18714
rect 17972 18630 18000 18686
rect 18616 18630 18644 19246
rect 18800 19174 18828 19264
rect 19064 19246 19116 19252
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 17972 13258 18000 18566
rect 18156 16998 18184 18566
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18708 9450 18736 18770
rect 19076 15094 19104 19246
rect 19536 18698 19564 20266
rect 20088 19378 20116 20266
rect 20456 19446 20484 20266
rect 20548 19514 20576 20266
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 18970 19656 19246
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 21376 13870 21404 20198
rect 21560 20058 21588 20334
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 22296 19242 22324 22200
rect 22756 20398 22784 22200
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 21546 17232 21602 17241
rect 21546 17167 21548 17176
rect 21600 17167 21602 17176
rect 21548 17138 21600 17144
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17420 5642 17448 6122
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5914 17908 6054
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 16948 5024 17000 5030
rect 17132 5024 17184 5030
rect 16948 4966 17000 4972
rect 17052 4984 17132 5012
rect 16960 4758 16988 4966
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 16868 3194 16896 4519
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16776 2582 16804 3130
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16960 2582 16988 3062
rect 17052 2990 17080 4984
rect 17132 4966 17184 4972
rect 17420 4622 17448 5578
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 4826 17540 5510
rect 17604 5302 17632 5578
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18602 5128 18658 5137
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17144 4078 17172 4422
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3602 18092 3878
rect 18156 3738 18184 5102
rect 18602 5063 18658 5072
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17960 3120 18012 3126
rect 17866 3088 17922 3097
rect 17960 3062 18012 3068
rect 17866 3023 17922 3032
rect 17880 2990 17908 3023
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17052 2774 17080 2926
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17052 2746 17264 2774
rect 17236 2650 17264 2746
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 16764 2576 16816 2582
rect 16764 2518 16816 2524
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 16132 800 16160 2314
rect 16592 800 16620 2314
rect 17052 800 17080 2314
rect 17512 800 17540 2858
rect 17972 2514 18000 3062
rect 18156 2990 18184 3674
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 2990 18644 5063
rect 18878 4176 18934 4185
rect 18878 4111 18934 4120
rect 18892 3058 18920 4111
rect 19076 3398 19104 6802
rect 21376 5914 21404 12650
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21546 5808 21602 5817
rect 21546 5743 21548 5752
rect 21600 5743 21602 5752
rect 21548 5714 21600 5720
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4690 20024 4966
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 19076 2990 19104 3334
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18064 2582 18092 2790
rect 18156 2650 18184 2790
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 19168 2582 19196 3402
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 19260 2446 19288 2994
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19444 2514 19472 2790
rect 19536 2582 19564 3062
rect 19720 2854 19748 3334
rect 20180 3126 20208 3606
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19996 2582 20024 3062
rect 20180 2990 20208 3062
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20720 2848 20772 2854
rect 20720 2790 20772 2796
rect 20732 2582 20760 2790
rect 19524 2576 19576 2582
rect 19524 2518 19576 2524
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 21008 2514 21036 4422
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 19892 2372 19944 2378
rect 19892 2314 19944 2320
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 17972 800 18000 2314
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18616 1170 18644 2246
rect 18432 1142 18644 1170
rect 18432 800 18460 1142
rect 18984 800 19012 2314
rect 19444 800 19472 2314
rect 19904 800 19932 2314
rect 20364 800 20392 2314
rect 20824 800 20852 2314
rect 21284 800 21312 2314
rect 21744 800 21772 2858
rect 22204 800 22232 2994
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22664 800 22692 2926
rect 3146 640 3202 649
rect 3146 575 3202 584
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22190 0 22246 800
rect 22650 0 22706 800
<< via2 >>
rect 3238 22616 3294 22672
rect 1766 21120 1822 21176
rect 1398 19780 1454 19816
rect 1398 19760 1400 19780
rect 1400 19760 1452 19780
rect 1452 19760 1454 19780
rect 1398 19236 1454 19272
rect 1398 19216 1400 19236
rect 1400 19216 1452 19236
rect 1452 19216 1454 19236
rect 1398 18828 1454 18864
rect 1398 18808 1400 18828
rect 1400 18808 1452 18828
rect 1452 18808 1454 18828
rect 1398 18284 1454 18320
rect 1858 20204 1860 20224
rect 1860 20204 1912 20224
rect 1912 20204 1914 20224
rect 1858 20168 1914 20204
rect 1674 19760 1730 19816
rect 2226 20712 2282 20768
rect 1398 18264 1400 18284
rect 1400 18264 1452 18284
rect 1452 18264 1454 18284
rect 1490 17876 1546 17912
rect 1490 17856 1492 17876
rect 1492 17856 1544 17876
rect 1544 17856 1546 17876
rect 2042 18828 2098 18864
rect 2042 18808 2044 18828
rect 2044 18808 2096 18828
rect 2096 18808 2098 18828
rect 2870 22072 2926 22128
rect 2778 21664 2834 21720
rect 2226 18128 2282 18184
rect 1858 17332 1914 17368
rect 1858 17312 1860 17332
rect 1860 17312 1912 17332
rect 1912 17312 1914 17332
rect 1490 16940 1492 16960
rect 1492 16940 1544 16960
rect 1544 16940 1546 16960
rect 1490 16904 1546 16940
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 2502 18300 2504 18320
rect 2504 18300 2556 18320
rect 2556 18300 2558 18320
rect 2502 18264 2558 18300
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 3514 18692 3570 18728
rect 3514 18672 3516 18692
rect 3516 18672 3568 18692
rect 3568 18672 3570 18692
rect 1398 15972 1454 16008
rect 1398 15952 1400 15972
rect 1400 15952 1452 15972
rect 1452 15952 1454 15972
rect 1398 15428 1454 15464
rect 1398 15408 1400 15428
rect 1400 15408 1452 15428
rect 1452 15408 1454 15428
rect 1398 15020 1454 15056
rect 1398 15000 1400 15020
rect 1400 15000 1452 15020
rect 1452 15000 1454 15020
rect 1398 14476 1454 14512
rect 1398 14456 1400 14476
rect 1400 14456 1452 14476
rect 1452 14456 1454 14476
rect 1490 14068 1546 14104
rect 1490 14048 1492 14068
rect 1492 14048 1544 14068
rect 1544 14048 1546 14068
rect 1490 13524 1546 13560
rect 1490 13504 1492 13524
rect 1492 13504 1544 13524
rect 1544 13504 1546 13524
rect 1398 11600 1454 11656
rect 1674 11212 1730 11248
rect 1674 11192 1676 11212
rect 1676 11192 1728 11212
rect 1728 11192 1730 11212
rect 1490 11056 1546 11112
rect 1398 10648 1454 10704
rect 1490 10124 1546 10160
rect 1490 10104 1492 10124
rect 1492 10104 1544 10124
rect 1544 10104 1546 10124
rect 1582 9696 1638 9752
rect 1398 9152 1454 9208
rect 1398 8744 1454 8800
rect 1398 7792 1454 7848
rect 1398 7384 1454 7440
rect 1950 8200 2006 8256
rect 1950 7284 1952 7304
rect 1952 7284 2004 7304
rect 2004 7284 2006 7304
rect 1950 7248 2006 7284
rect 1950 7112 2006 7168
rect 1674 6840 1730 6896
rect 1858 6840 1914 6896
rect 1398 6296 1454 6352
rect 1306 5888 1362 5944
rect 1582 6724 1638 6760
rect 1582 6704 1584 6724
rect 1584 6704 1636 6724
rect 1636 6704 1638 6724
rect 1674 5480 1730 5536
rect 1490 5344 1546 5400
rect 2870 13096 2926 13152
rect 2870 12552 2926 12608
rect 3054 12688 3110 12744
rect 3146 12144 3202 12200
rect 3146 11192 3202 11248
rect 2870 9424 2926 9480
rect 2226 7148 2228 7168
rect 2228 7148 2280 7168
rect 2280 7148 2282 7168
rect 2226 7112 2282 7148
rect 1030 2488 1086 2544
rect 1398 3984 1454 4040
rect 1674 4800 1730 4856
rect 1582 4528 1638 4584
rect 1858 4664 1914 4720
rect 1490 3440 1546 3496
rect 1214 1536 1270 1592
rect 1674 2624 1730 2680
rect 2778 7248 2834 7304
rect 3330 8472 3386 8528
rect 3514 9968 3570 10024
rect 3146 5072 3202 5128
rect 2962 4664 3018 4720
rect 2502 4256 2558 4312
rect 3054 4392 3110 4448
rect 2502 4120 2558 4176
rect 2594 3576 2650 3632
rect 2318 2932 2320 2952
rect 2320 2932 2372 2952
rect 2372 2932 2374 2952
rect 2318 2896 2374 2932
rect 2410 2488 2466 2544
rect 3054 4020 3056 4040
rect 3056 4020 3108 4040
rect 3108 4020 3110 4040
rect 3054 3984 3110 4020
rect 3422 5480 3478 5536
rect 3422 5208 3478 5264
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4710 18028 4712 18048
rect 4712 18028 4764 18048
rect 4764 18028 4766 18048
rect 4710 17992 4766 18028
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4526 11500 4528 11520
rect 4528 11500 4580 11520
rect 4580 11500 4582 11520
rect 4526 11464 4582 11500
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4250 10260 4306 10296
rect 4250 10240 4252 10260
rect 4252 10240 4304 10260
rect 4304 10240 4306 10260
rect 4158 9632 4214 9688
rect 5998 17992 6054 18048
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4342 8472 4398 8528
rect 3882 7384 3938 7440
rect 4250 7384 4306 7440
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4802 7112 4858 7168
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4710 6316 4766 6352
rect 4710 6296 4712 6316
rect 4712 6296 4764 6316
rect 4764 6296 4766 6316
rect 3330 3596 3386 3632
rect 3330 3576 3332 3596
rect 3332 3576 3384 3596
rect 3384 3576 3386 3596
rect 3330 3168 3386 3224
rect 1490 176 1546 232
rect 3514 3304 3570 3360
rect 3790 3304 3846 3360
rect 3606 2896 3662 2952
rect 3790 2896 3846 2952
rect 3790 2796 3792 2816
rect 3792 2796 3844 2816
rect 3844 2796 3846 2816
rect 3790 2760 3846 2796
rect 3698 2524 3700 2544
rect 3700 2524 3752 2544
rect 3752 2524 3754 2544
rect 3698 2488 3754 2524
rect 3790 1128 3846 1184
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4250 4256 4306 4312
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4526 3848 4582 3904
rect 4986 4664 5042 4720
rect 4986 4392 5042 4448
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4618 2896 4674 2952
rect 4066 2080 4122 2136
rect 4986 3304 5042 3360
rect 4894 2896 4950 2952
rect 4986 2624 5042 2680
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5722 9968 5778 10024
rect 5538 7148 5540 7168
rect 5540 7148 5592 7168
rect 5592 7148 5594 7168
rect 5538 7112 5594 7148
rect 5446 3576 5502 3632
rect 5722 6296 5778 6352
rect 6642 18808 6698 18864
rect 5630 4936 5686 4992
rect 6458 9424 6514 9480
rect 6642 9424 6698 9480
rect 6274 5888 6330 5944
rect 6090 4800 6146 4856
rect 5814 3848 5870 3904
rect 5814 3732 5870 3768
rect 5814 3712 5816 3732
rect 5816 3712 5868 3732
rect 5868 3712 5870 3732
rect 5814 3168 5870 3224
rect 6458 4528 6514 4584
rect 6550 4428 6552 4448
rect 6552 4428 6604 4448
rect 6604 4428 6606 4448
rect 6550 4392 6606 4428
rect 7378 11464 7434 11520
rect 6826 3712 6882 3768
rect 6918 3440 6974 3496
rect 6826 2624 6882 2680
rect 7194 5092 7250 5128
rect 7194 5072 7196 5092
rect 7196 5072 7248 5092
rect 7248 5072 7250 5092
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 9034 19760 9090 19816
rect 9402 18264 9458 18320
rect 9218 13796 9274 13832
rect 9218 13776 9220 13796
rect 9220 13776 9272 13796
rect 9272 13776 9274 13796
rect 9954 18128 10010 18184
rect 9678 14000 9734 14002
rect 9678 13948 9680 14000
rect 9680 13948 9732 14000
rect 9732 13948 9734 14000
rect 9678 13946 9734 13948
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10230 18672 10286 18728
rect 9402 12708 9458 12744
rect 9402 12688 9404 12708
rect 9404 12688 9456 12708
rect 9456 12688 9458 12708
rect 8206 8356 8262 8392
rect 8206 8336 8208 8356
rect 8208 8336 8260 8356
rect 8260 8336 8262 8356
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7930 6724 7986 6760
rect 7930 6704 7932 6724
rect 7932 6704 7984 6724
rect 7984 6704 7986 6724
rect 7378 4120 7434 4176
rect 7654 4256 7710 4312
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 8114 5788 8116 5808
rect 8116 5788 8168 5808
rect 8168 5788 8170 5808
rect 8114 5752 8170 5788
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8666 6840 8722 6896
rect 8482 3440 8538 3496
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8758 3304 8814 3360
rect 9218 5072 9274 5128
rect 10230 13776 10286 13832
rect 9678 8472 9734 8528
rect 9770 6724 9826 6760
rect 9770 6704 9772 6724
rect 9772 6704 9824 6724
rect 9824 6704 9826 6724
rect 9586 5208 9642 5264
rect 9770 4820 9826 4856
rect 9770 4800 9772 4820
rect 9772 4800 9824 4820
rect 9824 4800 9826 4820
rect 9402 3984 9458 4040
rect 9402 3440 9458 3496
rect 9770 3848 9826 3904
rect 11058 14612 11114 14648
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11058 14592 11060 14612
rect 11060 14592 11112 14612
rect 11112 14592 11114 14612
rect 10506 6704 10562 6760
rect 10506 4684 10562 4720
rect 10506 4664 10508 4684
rect 10508 4664 10560 4684
rect 10560 4664 10562 4684
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11794 13912 11850 13968
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10782 3032 10838 3088
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11150 4120 11206 4176
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11794 12844 11850 12880
rect 11794 12824 11796 12844
rect 11796 12824 11848 12844
rect 11848 12824 11850 12844
rect 11794 11600 11850 11656
rect 11794 9288 11850 9344
rect 12162 9424 12218 9480
rect 12070 9288 12126 9344
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 12254 6704 12310 6760
rect 11978 5092 12034 5128
rect 11978 5072 11980 5092
rect 11980 5072 12032 5092
rect 12032 5072 12034 5092
rect 12070 4548 12126 4584
rect 12070 4528 12072 4548
rect 12072 4528 12124 4548
rect 12124 4528 12126 4548
rect 11978 3884 11980 3904
rect 11980 3884 12032 3904
rect 12032 3884 12034 3904
rect 11978 3848 12034 3884
rect 12438 6724 12494 6760
rect 12438 6704 12440 6724
rect 12440 6704 12492 6724
rect 12492 6704 12494 6724
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12346 3984 12402 4040
rect 13726 12824 13782 12880
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14646 14592 14702 14648
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14002 4820 14058 4856
rect 14002 4800 14004 4820
rect 14004 4800 14056 4820
rect 14056 4800 14058 4820
rect 13266 4140 13322 4176
rect 13266 4120 13268 4140
rect 13268 4120 13320 4140
rect 13320 4120 13322 4140
rect 14186 8356 14242 8392
rect 14186 8336 14188 8356
rect 14188 8336 14240 8356
rect 14240 8336 14242 8356
rect 14738 11600 14794 11656
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14738 4528 14794 4584
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 21546 17196 21602 17232
rect 21546 17176 21548 17196
rect 21548 17176 21600 17196
rect 21600 17176 21602 17196
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 16854 4528 16910 4584
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18602 5072 18658 5128
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 17866 3032 17922 3088
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18878 4120 18934 4176
rect 21546 5772 21602 5808
rect 21546 5752 21548 5772
rect 21548 5752 21600 5772
rect 21600 5752 21602 5772
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 3146 584 3202 640
<< metal3 >>
rect 0 22674 800 22704
rect 3233 22674 3299 22677
rect 0 22672 3299 22674
rect 0 22616 3238 22672
rect 3294 22616 3299 22672
rect 0 22614 3299 22616
rect 0 22584 800 22614
rect 3233 22611 3299 22614
rect 0 22130 800 22160
rect 2865 22130 2931 22133
rect 0 22128 2931 22130
rect 0 22072 2870 22128
rect 2926 22072 2931 22128
rect 0 22070 2931 22072
rect 0 22040 800 22070
rect 2865 22067 2931 22070
rect 0 21722 800 21752
rect 2773 21722 2839 21725
rect 0 21720 2839 21722
rect 0 21664 2778 21720
rect 2834 21664 2839 21720
rect 0 21662 2839 21664
rect 0 21632 800 21662
rect 2773 21659 2839 21662
rect 0 21178 800 21208
rect 1761 21178 1827 21181
rect 0 21176 1827 21178
rect 0 21120 1766 21176
rect 1822 21120 1827 21176
rect 0 21118 1827 21120
rect 0 21088 800 21118
rect 1761 21115 1827 21118
rect 0 20770 800 20800
rect 2221 20770 2287 20773
rect 0 20768 2287 20770
rect 0 20712 2226 20768
rect 2282 20712 2287 20768
rect 0 20710 2287 20712
rect 0 20680 800 20710
rect 2221 20707 2287 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20226 800 20256
rect 1853 20226 1919 20229
rect 0 20224 1919 20226
rect 0 20168 1858 20224
rect 1914 20168 1919 20224
rect 0 20166 1919 20168
rect 0 20136 800 20166
rect 1853 20163 1919 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 1669 19818 1735 19821
rect 9029 19818 9095 19821
rect 1669 19816 9095 19818
rect 1669 19760 1674 19816
rect 1730 19760 9034 19816
rect 9090 19760 9095 19816
rect 1669 19758 9095 19760
rect 1669 19755 1735 19758
rect 9029 19755 9095 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19274 800 19304
rect 1393 19274 1459 19277
rect 0 19272 1459 19274
rect 0 19216 1398 19272
rect 1454 19216 1459 19272
rect 0 19214 1459 19216
rect 0 19184 800 19214
rect 1393 19211 1459 19214
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 800 18806
rect 1393 18803 1459 18806
rect 2037 18866 2103 18869
rect 6637 18866 6703 18869
rect 2037 18864 6703 18866
rect 2037 18808 2042 18864
rect 2098 18808 6642 18864
rect 6698 18808 6703 18864
rect 2037 18806 6703 18808
rect 2037 18803 2103 18806
rect 6637 18803 6703 18806
rect 3509 18730 3575 18733
rect 10225 18730 10291 18733
rect 3509 18728 10291 18730
rect 3509 18672 3514 18728
rect 3570 18672 10230 18728
rect 10286 18672 10291 18728
rect 3509 18670 10291 18672
rect 3509 18667 3575 18670
rect 10225 18667 10291 18670
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 0 18322 800 18352
rect 1393 18322 1459 18325
rect 0 18320 1459 18322
rect 0 18264 1398 18320
rect 1454 18264 1459 18320
rect 0 18262 1459 18264
rect 0 18232 800 18262
rect 1393 18259 1459 18262
rect 2497 18322 2563 18325
rect 9397 18322 9463 18325
rect 2497 18320 9463 18322
rect 2497 18264 2502 18320
rect 2558 18264 9402 18320
rect 9458 18264 9463 18320
rect 2497 18262 9463 18264
rect 2497 18259 2563 18262
rect 9397 18259 9463 18262
rect 2221 18186 2287 18189
rect 9949 18186 10015 18189
rect 2221 18184 10015 18186
rect 2221 18128 2226 18184
rect 2282 18128 9954 18184
rect 10010 18128 10015 18184
rect 2221 18126 10015 18128
rect 2221 18123 2287 18126
rect 9949 18123 10015 18126
rect 4705 18050 4771 18053
rect 5993 18050 6059 18053
rect 4705 18048 6059 18050
rect 4705 17992 4710 18048
rect 4766 17992 5998 18048
rect 6054 17992 6059 18048
rect 4705 17990 6059 17992
rect 4705 17987 4771 17990
rect 5993 17987 6059 17990
rect 7874 17984 8194 17985
rect 0 17914 800 17944
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 1485 17914 1551 17917
rect 0 17912 1551 17914
rect 0 17856 1490 17912
rect 1546 17856 1551 17912
rect 0 17854 1551 17856
rect 0 17824 800 17854
rect 1485 17851 1551 17854
rect 4409 17440 4729 17441
rect 0 17370 800 17400
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 1853 17370 1919 17373
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 800 17310
rect 1853 17307 1919 17310
rect 21541 17234 21607 17237
rect 22200 17234 23000 17264
rect 21541 17232 23000 17234
rect 21541 17176 21546 17232
rect 21602 17176 23000 17232
rect 21541 17174 23000 17176
rect 21541 17171 21607 17174
rect 22200 17144 23000 17174
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16010 800 16040
rect 1393 16010 1459 16013
rect 0 16008 1459 16010
rect 0 15952 1398 16008
rect 1454 15952 1459 16008
rect 0 15950 1459 15952
rect 0 15920 800 15950
rect 1393 15947 1459 15950
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15466 800 15496
rect 1393 15466 1459 15469
rect 0 15464 1459 15466
rect 0 15408 1398 15464
rect 1454 15408 1459 15464
rect 0 15406 1459 15408
rect 0 15376 800 15406
rect 1393 15403 1459 15406
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 11053 14650 11119 14653
rect 14641 14650 14707 14653
rect 11053 14648 14707 14650
rect 11053 14592 11058 14648
rect 11114 14592 14646 14648
rect 14702 14592 14707 14648
rect 11053 14590 14707 14592
rect 11053 14587 11119 14590
rect 14641 14587 14707 14590
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 4409 14176 4729 14177
rect 0 14106 800 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 1485 14106 1551 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 800 14046
rect 1485 14043 1551 14046
rect 9673 14004 9739 14007
rect 9630 14002 9739 14004
rect 9630 13946 9678 14002
rect 9734 13970 9739 14002
rect 11789 13970 11855 13973
rect 9734 13968 11855 13970
rect 9734 13946 11794 13968
rect 9630 13912 11794 13946
rect 11850 13912 11855 13968
rect 9630 13910 11855 13912
rect 11789 13907 11855 13910
rect 9213 13834 9279 13837
rect 10225 13834 10291 13837
rect 9213 13832 10291 13834
rect 9213 13776 9218 13832
rect 9274 13776 10230 13832
rect 10286 13776 10291 13832
rect 9213 13774 10291 13776
rect 9213 13771 9279 13774
rect 10225 13771 10291 13774
rect 7874 13632 8194 13633
rect 0 13562 800 13592
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 0 13154 800 13184
rect 2865 13154 2931 13157
rect 0 13152 2931 13154
rect 0 13096 2870 13152
rect 2926 13096 2931 13152
rect 0 13094 2931 13096
rect 0 13064 800 13094
rect 2865 13091 2931 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 11789 12882 11855 12885
rect 13721 12882 13787 12885
rect 11789 12880 13787 12882
rect 11789 12824 11794 12880
rect 11850 12824 13726 12880
rect 13782 12824 13787 12880
rect 11789 12822 13787 12824
rect 11789 12819 11855 12822
rect 13721 12819 13787 12822
rect 3049 12746 3115 12749
rect 9397 12746 9463 12749
rect 3049 12744 9463 12746
rect 3049 12688 3054 12744
rect 3110 12688 9402 12744
rect 9458 12688 9463 12744
rect 3049 12686 9463 12688
rect 3049 12683 3115 12686
rect 9397 12683 9463 12686
rect 0 12610 800 12640
rect 2865 12610 2931 12613
rect 0 12608 2931 12610
rect 0 12552 2870 12608
rect 2926 12552 2931 12608
rect 0 12550 2931 12552
rect 0 12520 800 12550
rect 2865 12547 2931 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12202 800 12232
rect 3141 12202 3207 12205
rect 0 12200 3207 12202
rect 0 12144 3146 12200
rect 3202 12144 3207 12200
rect 0 12142 3207 12144
rect 0 12112 800 12142
rect 3141 12139 3207 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 11789 11658 11855 11661
rect 14733 11658 14799 11661
rect 11789 11656 14799 11658
rect 11789 11600 11794 11656
rect 11850 11600 14738 11656
rect 14794 11600 14799 11656
rect 11789 11598 14799 11600
rect 11789 11595 11855 11598
rect 14733 11595 14799 11598
rect 4521 11522 4587 11525
rect 4838 11522 4844 11524
rect 4521 11520 4844 11522
rect 4521 11464 4526 11520
rect 4582 11464 4844 11520
rect 4521 11462 4844 11464
rect 4521 11459 4587 11462
rect 4838 11460 4844 11462
rect 4908 11522 4914 11524
rect 7373 11522 7439 11525
rect 4908 11520 7439 11522
rect 4908 11464 7378 11520
rect 7434 11464 7439 11520
rect 4908 11462 7439 11464
rect 4908 11460 4914 11462
rect 7373 11459 7439 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 1669 11250 1735 11253
rect 3141 11250 3207 11253
rect 1669 11248 3207 11250
rect 1669 11192 1674 11248
rect 1730 11192 3146 11248
rect 3202 11192 3207 11248
rect 1669 11190 3207 11192
rect 1669 11187 1735 11190
rect 3141 11187 3207 11190
rect 0 11114 800 11144
rect 1485 11114 1551 11117
rect 0 11112 1551 11114
rect 0 11056 1490 11112
rect 1546 11056 1551 11112
rect 0 11054 1551 11056
rect 0 11024 800 11054
rect 1485 11051 1551 11054
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 0 10706 800 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 800 10646
rect 1393 10643 1459 10646
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 4102 10236 4108 10300
rect 4172 10298 4178 10300
rect 4245 10298 4311 10301
rect 4172 10296 4311 10298
rect 4172 10240 4250 10296
rect 4306 10240 4311 10296
rect 4172 10238 4311 10240
rect 4172 10236 4178 10238
rect 4245 10235 4311 10238
rect 0 10162 800 10192
rect 1485 10162 1551 10165
rect 0 10160 1551 10162
rect 0 10104 1490 10160
rect 1546 10104 1551 10160
rect 0 10102 1551 10104
rect 0 10072 800 10102
rect 1485 10099 1551 10102
rect 3509 10026 3575 10029
rect 5717 10026 5783 10029
rect 3509 10024 5783 10026
rect 3509 9968 3514 10024
rect 3570 9968 5722 10024
rect 5778 9968 5783 10024
rect 3509 9966 5783 9968
rect 3509 9963 3575 9966
rect 5717 9963 5783 9966
rect 4409 9824 4729 9825
rect 0 9754 800 9784
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 1577 9754 1643 9757
rect 0 9752 1643 9754
rect 0 9696 1582 9752
rect 1638 9696 1643 9752
rect 0 9694 1643 9696
rect 0 9664 800 9694
rect 1577 9691 1643 9694
rect 4102 9692 4108 9756
rect 4172 9693 4178 9756
rect 4172 9692 4219 9693
rect 4110 9688 4219 9692
rect 4110 9632 4158 9688
rect 4214 9632 4219 9688
rect 4110 9630 4219 9632
rect 4153 9627 4219 9630
rect 2865 9482 2931 9485
rect 6453 9482 6519 9485
rect 2865 9480 6519 9482
rect 2865 9424 2870 9480
rect 2926 9424 6458 9480
rect 6514 9424 6519 9480
rect 2865 9422 6519 9424
rect 2865 9419 2931 9422
rect 6453 9419 6519 9422
rect 6637 9482 6703 9485
rect 12157 9482 12223 9485
rect 6637 9480 12223 9482
rect 6637 9424 6642 9480
rect 6698 9424 12162 9480
rect 12218 9424 12223 9480
rect 6637 9422 12223 9424
rect 6637 9419 6703 9422
rect 12157 9419 12223 9422
rect 11789 9346 11855 9349
rect 12065 9346 12131 9349
rect 11789 9344 12131 9346
rect 11789 9288 11794 9344
rect 11850 9288 12070 9344
rect 12126 9288 12131 9344
rect 11789 9286 12131 9288
rect 11789 9283 11855 9286
rect 12065 9283 12131 9286
rect 7874 9280 8194 9281
rect 0 9210 800 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 0 8802 800 8832
rect 1393 8802 1459 8805
rect 0 8800 1459 8802
rect 0 8744 1398 8800
rect 1454 8744 1459 8800
rect 0 8742 1459 8744
rect 0 8712 800 8742
rect 1393 8739 1459 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 3325 8530 3391 8533
rect 4337 8530 4403 8533
rect 9673 8530 9739 8533
rect 3325 8528 4403 8530
rect 3325 8472 3330 8528
rect 3386 8472 4342 8528
rect 4398 8472 4403 8528
rect 3325 8470 4403 8472
rect 3325 8467 3391 8470
rect 4337 8467 4403 8470
rect 6870 8528 9739 8530
rect 6870 8472 9678 8528
rect 9734 8472 9739 8528
rect 6870 8470 9739 8472
rect 0 8258 800 8288
rect 1945 8258 2011 8261
rect 6870 8260 6930 8470
rect 9673 8467 9739 8470
rect 8201 8394 8267 8397
rect 14181 8394 14247 8397
rect 8201 8392 14247 8394
rect 8201 8336 8206 8392
rect 8262 8336 14186 8392
rect 14242 8336 14247 8392
rect 8201 8334 14247 8336
rect 8201 8331 8267 8334
rect 14181 8331 14247 8334
rect 0 8256 2011 8258
rect 0 8200 1950 8256
rect 2006 8200 2011 8256
rect 0 8198 2011 8200
rect 0 8168 800 8198
rect 1945 8195 2011 8198
rect 6862 8196 6868 8260
rect 6932 8196 6938 8260
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 0 7850 800 7880
rect 1393 7850 1459 7853
rect 0 7848 1459 7850
rect 0 7792 1398 7848
rect 1454 7792 1459 7848
rect 0 7790 1459 7792
rect 0 7760 800 7790
rect 1393 7787 1459 7790
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 1393 7442 1459 7445
rect 3877 7442 3943 7445
rect 1393 7440 3943 7442
rect 1393 7384 1398 7440
rect 1454 7384 3882 7440
rect 3938 7384 3943 7440
rect 1393 7382 3943 7384
rect 1393 7379 1459 7382
rect 3877 7379 3943 7382
rect 4245 7442 4311 7445
rect 6862 7442 6868 7444
rect 4245 7440 6868 7442
rect 4245 7384 4250 7440
rect 4306 7384 6868 7440
rect 4245 7382 6868 7384
rect 4245 7379 4311 7382
rect 6862 7380 6868 7382
rect 6932 7380 6938 7444
rect 0 7306 800 7336
rect 1945 7306 2011 7309
rect 2773 7306 2839 7309
rect 0 7304 2011 7306
rect 0 7248 1950 7304
rect 2006 7248 2011 7304
rect 0 7246 2011 7248
rect 0 7216 800 7246
rect 1945 7243 2011 7246
rect 2086 7304 5596 7306
rect 2086 7248 2778 7304
rect 2834 7248 5596 7304
rect 2086 7246 5596 7248
rect 1945 7170 2011 7173
rect 2086 7170 2146 7246
rect 2773 7243 2839 7246
rect 5536 7173 5596 7246
rect 1945 7168 2146 7170
rect 1945 7112 1950 7168
rect 2006 7112 2146 7168
rect 1945 7110 2146 7112
rect 2221 7170 2287 7173
rect 4797 7170 4863 7173
rect 5533 7172 5599 7173
rect 5533 7170 5580 7172
rect 2221 7168 4863 7170
rect 2221 7112 2226 7168
rect 2282 7112 4802 7168
rect 4858 7112 4863 7168
rect 2221 7110 4863 7112
rect 5488 7168 5580 7170
rect 5488 7112 5538 7168
rect 5488 7110 5580 7112
rect 1945 7107 2011 7110
rect 2221 7107 2287 7110
rect 4797 7107 4863 7110
rect 5533 7108 5580 7110
rect 5644 7108 5650 7172
rect 5533 7107 5599 7108
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6898 800 6928
rect 1669 6898 1735 6901
rect 0 6896 1735 6898
rect 0 6840 1674 6896
rect 1730 6840 1735 6896
rect 0 6838 1735 6840
rect 0 6808 800 6838
rect 1669 6835 1735 6838
rect 1853 6898 1919 6901
rect 8661 6898 8727 6901
rect 1853 6896 8727 6898
rect 1853 6840 1858 6896
rect 1914 6840 8666 6896
rect 8722 6840 8727 6896
rect 1853 6838 8727 6840
rect 1853 6835 1919 6838
rect 8661 6835 8727 6838
rect 1577 6762 1643 6765
rect 7925 6762 7991 6765
rect 1577 6760 7991 6762
rect 1577 6704 1582 6760
rect 1638 6704 7930 6760
rect 7986 6704 7991 6760
rect 1577 6702 7991 6704
rect 1577 6699 1643 6702
rect 7925 6699 7991 6702
rect 9765 6762 9831 6765
rect 10501 6762 10567 6765
rect 9765 6760 10567 6762
rect 9765 6704 9770 6760
rect 9826 6704 10506 6760
rect 10562 6704 10567 6760
rect 9765 6702 10567 6704
rect 9765 6699 9831 6702
rect 10501 6699 10567 6702
rect 12249 6762 12315 6765
rect 12433 6762 12499 6765
rect 12249 6760 12499 6762
rect 12249 6704 12254 6760
rect 12310 6704 12438 6760
rect 12494 6704 12499 6760
rect 12249 6702 12499 6704
rect 12249 6699 12315 6702
rect 12433 6699 12499 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6354 800 6384
rect 1393 6354 1459 6357
rect 0 6352 1459 6354
rect 0 6296 1398 6352
rect 1454 6296 1459 6352
rect 0 6294 1459 6296
rect 0 6264 800 6294
rect 1393 6291 1459 6294
rect 4705 6354 4771 6357
rect 5717 6354 5783 6357
rect 4705 6352 5783 6354
rect 4705 6296 4710 6352
rect 4766 6296 5722 6352
rect 5778 6296 5783 6352
rect 4705 6294 5783 6296
rect 4705 6291 4771 6294
rect 5717 6291 5783 6294
rect 7874 6016 8194 6017
rect 0 5946 800 5976
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 1301 5946 1367 5949
rect 0 5944 1367 5946
rect 0 5888 1306 5944
rect 1362 5888 1367 5944
rect 0 5886 1367 5888
rect 0 5856 800 5886
rect 1301 5883 1367 5886
rect 6269 5946 6335 5949
rect 6269 5944 7482 5946
rect 6269 5888 6274 5944
rect 6330 5888 7482 5944
rect 6269 5886 7482 5888
rect 6269 5883 6335 5886
rect 7422 5810 7482 5886
rect 8109 5810 8175 5813
rect 7422 5808 8175 5810
rect 7422 5752 8114 5808
rect 8170 5752 8175 5808
rect 7422 5750 8175 5752
rect 8109 5747 8175 5750
rect 21541 5810 21607 5813
rect 22200 5810 23000 5840
rect 21541 5808 23000 5810
rect 21541 5752 21546 5808
rect 21602 5752 23000 5808
rect 21541 5750 23000 5752
rect 21541 5747 21607 5750
rect 22200 5720 23000 5750
rect 1669 5538 1735 5541
rect 3417 5538 3483 5541
rect 1669 5536 3483 5538
rect 1669 5480 1674 5536
rect 1730 5480 3422 5536
rect 3478 5480 3483 5536
rect 1669 5478 3483 5480
rect 1669 5475 1735 5478
rect 0 5402 800 5432
rect 1485 5402 1551 5405
rect 0 5400 1551 5402
rect 0 5344 1490 5400
rect 1546 5344 1551 5400
rect 0 5342 1551 5344
rect 0 5312 800 5342
rect 1485 5339 1551 5342
rect 0 4994 800 5024
rect 2730 4994 2790 5478
rect 3417 5475 3483 5478
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 3417 5266 3483 5269
rect 9581 5266 9647 5269
rect 3417 5264 9647 5266
rect 3417 5208 3422 5264
rect 3478 5208 9586 5264
rect 9642 5208 9647 5264
rect 3417 5206 9647 5208
rect 3417 5203 3483 5206
rect 9581 5203 9647 5206
rect 3141 5130 3207 5133
rect 7189 5130 7255 5133
rect 9213 5130 9279 5133
rect 3141 5128 9279 5130
rect 3141 5072 3146 5128
rect 3202 5072 7194 5128
rect 7250 5072 9218 5128
rect 9274 5072 9279 5128
rect 3141 5070 9279 5072
rect 3141 5067 3207 5070
rect 7189 5067 7255 5070
rect 9213 5067 9279 5070
rect 11973 5130 12039 5133
rect 18597 5130 18663 5133
rect 11973 5128 18663 5130
rect 11973 5072 11978 5128
rect 12034 5072 18602 5128
rect 18658 5072 18663 5128
rect 11973 5070 18663 5072
rect 11973 5067 12039 5070
rect 18597 5067 18663 5070
rect 0 4934 2790 4994
rect 5625 4994 5691 4997
rect 5758 4994 5764 4996
rect 5625 4992 5764 4994
rect 5625 4936 5630 4992
rect 5686 4936 5764 4992
rect 5625 4934 5764 4936
rect 0 4904 800 4934
rect 5625 4931 5691 4934
rect 5758 4932 5764 4934
rect 5828 4932 5834 4996
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 1669 4858 1735 4861
rect 6085 4858 6151 4861
rect 1669 4856 6151 4858
rect 1669 4800 1674 4856
rect 1730 4800 6090 4856
rect 6146 4800 6151 4856
rect 1669 4798 6151 4800
rect 1669 4795 1735 4798
rect 6085 4795 6151 4798
rect 9765 4858 9831 4861
rect 13997 4858 14063 4861
rect 9765 4856 14063 4858
rect 9765 4800 9770 4856
rect 9826 4800 14002 4856
rect 14058 4800 14063 4856
rect 9765 4798 14063 4800
rect 9765 4795 9831 4798
rect 13997 4795 14063 4798
rect 1853 4722 1919 4725
rect 2957 4722 3023 4725
rect 4981 4722 5047 4725
rect 1853 4720 5047 4722
rect 1853 4664 1858 4720
rect 1914 4664 2962 4720
rect 3018 4664 4986 4720
rect 5042 4664 5047 4720
rect 1853 4662 5047 4664
rect 1853 4659 1919 4662
rect 2957 4659 3023 4662
rect 4981 4659 5047 4662
rect 5758 4660 5764 4724
rect 5828 4722 5834 4724
rect 10501 4722 10567 4725
rect 5828 4720 10567 4722
rect 5828 4664 10506 4720
rect 10562 4664 10567 4720
rect 5828 4662 10567 4664
rect 5828 4660 5834 4662
rect 10501 4659 10567 4662
rect 1577 4586 1643 4589
rect 6453 4586 6519 4589
rect 1577 4584 6519 4586
rect 1577 4528 1582 4584
rect 1638 4528 6458 4584
rect 6514 4528 6519 4584
rect 1577 4526 6519 4528
rect 1577 4523 1643 4526
rect 6453 4523 6519 4526
rect 12065 4586 12131 4589
rect 14733 4586 14799 4589
rect 16849 4586 16915 4589
rect 12065 4584 16915 4586
rect 12065 4528 12070 4584
rect 12126 4528 14738 4584
rect 14794 4528 16854 4584
rect 16910 4528 16915 4584
rect 12065 4526 16915 4528
rect 12065 4523 12131 4526
rect 14733 4523 14799 4526
rect 16849 4523 16915 4526
rect 0 4450 800 4480
rect 3049 4450 3115 4453
rect 0 4448 3115 4450
rect 0 4392 3054 4448
rect 3110 4392 3115 4448
rect 0 4390 3115 4392
rect 0 4360 800 4390
rect 3049 4387 3115 4390
rect 4981 4450 5047 4453
rect 6545 4450 6611 4453
rect 4981 4448 6611 4450
rect 4981 4392 4986 4448
rect 5042 4392 6550 4448
rect 6606 4392 6611 4448
rect 4981 4390 6611 4392
rect 4981 4387 5047 4390
rect 6545 4387 6611 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 2497 4314 2563 4317
rect 4245 4314 4311 4317
rect 2497 4312 4311 4314
rect 2497 4256 2502 4312
rect 2558 4256 4250 4312
rect 4306 4256 4311 4312
rect 2497 4254 4311 4256
rect 2497 4251 2563 4254
rect 4245 4251 4311 4254
rect 7649 4314 7715 4317
rect 7649 4312 9690 4314
rect 7649 4256 7654 4312
rect 7710 4256 9690 4312
rect 7649 4254 9690 4256
rect 7649 4251 7715 4254
rect 2497 4178 2563 4181
rect 7373 4178 7439 4181
rect 2497 4176 7439 4178
rect 2497 4120 2502 4176
rect 2558 4120 7378 4176
rect 7434 4120 7439 4176
rect 2497 4118 7439 4120
rect 2497 4115 2563 4118
rect 7373 4115 7439 4118
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 3049 4042 3115 4045
rect 9397 4042 9463 4045
rect 3049 4040 9463 4042
rect 3049 3984 3054 4040
rect 3110 3984 9402 4040
rect 9458 3984 9463 4040
rect 3049 3982 9463 3984
rect 9630 4042 9690 4254
rect 11145 4178 11211 4181
rect 13261 4178 13327 4181
rect 18873 4178 18939 4181
rect 11145 4176 18939 4178
rect 11145 4120 11150 4176
rect 11206 4120 13266 4176
rect 13322 4120 18878 4176
rect 18934 4120 18939 4176
rect 11145 4118 18939 4120
rect 11145 4115 11211 4118
rect 13261 4115 13327 4118
rect 18873 4115 18939 4118
rect 12341 4042 12407 4045
rect 9630 4040 12407 4042
rect 9630 3984 12346 4040
rect 12402 3984 12407 4040
rect 9630 3982 12407 3984
rect 3049 3979 3115 3982
rect 9397 3979 9463 3982
rect 12341 3979 12407 3982
rect 4521 3906 4587 3909
rect 5809 3906 5875 3909
rect 4521 3904 5875 3906
rect 4521 3848 4526 3904
rect 4582 3848 5814 3904
rect 5870 3848 5875 3904
rect 4521 3846 5875 3848
rect 4521 3843 4587 3846
rect 5809 3843 5875 3846
rect 9765 3906 9831 3909
rect 11973 3906 12039 3909
rect 9765 3904 12039 3906
rect 9765 3848 9770 3904
rect 9826 3848 11978 3904
rect 12034 3848 12039 3904
rect 9765 3846 12039 3848
rect 9765 3843 9831 3846
rect 11973 3843 12039 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 5809 3770 5875 3773
rect 6821 3770 6887 3773
rect 5809 3768 6887 3770
rect 5809 3712 5814 3768
rect 5870 3712 6826 3768
rect 6882 3712 6887 3768
rect 5809 3710 6887 3712
rect 5809 3707 5875 3710
rect 6821 3707 6887 3710
rect 2589 3634 2655 3637
rect 3325 3634 3391 3637
rect 5441 3634 5507 3637
rect 2589 3632 2790 3634
rect 2589 3576 2594 3632
rect 2650 3576 2790 3632
rect 2589 3574 2790 3576
rect 2589 3571 2655 3574
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 2730 3498 2790 3574
rect 3325 3632 5507 3634
rect 3325 3576 3330 3632
rect 3386 3576 5446 3632
rect 5502 3576 5507 3632
rect 3325 3574 5507 3576
rect 3325 3571 3391 3574
rect 5441 3571 5507 3574
rect 6913 3498 6979 3501
rect 2730 3496 6979 3498
rect 2730 3440 6918 3496
rect 6974 3440 6979 3496
rect 2730 3438 6979 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 6913 3435 6979 3438
rect 8477 3498 8543 3501
rect 9397 3498 9463 3501
rect 8477 3496 9463 3498
rect 8477 3440 8482 3496
rect 8538 3440 9402 3496
rect 9458 3440 9463 3496
rect 8477 3438 9463 3440
rect 8477 3435 8543 3438
rect 9397 3435 9463 3438
rect 3509 3362 3575 3365
rect 3785 3362 3851 3365
rect 3509 3360 3851 3362
rect 3509 3304 3514 3360
rect 3570 3304 3790 3360
rect 3846 3304 3851 3360
rect 3509 3302 3851 3304
rect 3509 3299 3575 3302
rect 3785 3299 3851 3302
rect 4981 3362 5047 3365
rect 8753 3362 8819 3365
rect 4981 3360 8819 3362
rect 4981 3304 4986 3360
rect 5042 3304 8758 3360
rect 8814 3304 8819 3360
rect 4981 3302 8819 3304
rect 4981 3299 5047 3302
rect 8753 3299 8819 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 3325 3226 3391 3229
rect 3006 3224 3391 3226
rect 3006 3168 3330 3224
rect 3386 3168 3391 3224
rect 3006 3166 3391 3168
rect 0 3090 800 3120
rect 3006 3090 3066 3166
rect 3325 3163 3391 3166
rect 5574 3164 5580 3228
rect 5644 3226 5650 3228
rect 5809 3226 5875 3229
rect 5644 3224 5875 3226
rect 5644 3168 5814 3224
rect 5870 3168 5875 3224
rect 5644 3166 5875 3168
rect 5644 3164 5650 3166
rect 5809 3163 5875 3166
rect 0 3030 3066 3090
rect 10777 3090 10843 3093
rect 17861 3090 17927 3093
rect 10777 3088 17927 3090
rect 10777 3032 10782 3088
rect 10838 3032 17866 3088
rect 17922 3032 17927 3088
rect 10777 3030 17927 3032
rect 0 3000 800 3030
rect 10777 3027 10843 3030
rect 17861 3027 17927 3030
rect 2313 2954 2379 2957
rect 3601 2954 3667 2957
rect 2313 2952 3667 2954
rect 2313 2896 2318 2952
rect 2374 2896 3606 2952
rect 3662 2896 3667 2952
rect 2313 2894 3667 2896
rect 2313 2891 2379 2894
rect 3601 2891 3667 2894
rect 3785 2954 3851 2957
rect 4613 2954 4679 2957
rect 4889 2956 4955 2957
rect 3785 2952 4679 2954
rect 3785 2896 3790 2952
rect 3846 2896 4618 2952
rect 4674 2896 4679 2952
rect 3785 2894 4679 2896
rect 3785 2891 3851 2894
rect 4613 2891 4679 2894
rect 4838 2892 4844 2956
rect 4908 2954 4955 2956
rect 4908 2952 5000 2954
rect 4950 2896 5000 2952
rect 4908 2894 5000 2896
rect 4908 2892 4955 2894
rect 4889 2891 4955 2892
rect 3785 2818 3851 2821
rect 5758 2818 5764 2820
rect 3785 2816 5764 2818
rect 3785 2760 3790 2816
rect 3846 2760 5764 2816
rect 3785 2758 5764 2760
rect 3785 2755 3851 2758
rect 5758 2756 5764 2758
rect 5828 2756 5834 2820
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 1669 2682 1735 2685
rect 4981 2682 5047 2685
rect 6821 2684 6887 2685
rect 6821 2682 6868 2684
rect 1669 2680 5047 2682
rect 1669 2624 1674 2680
rect 1730 2624 4986 2680
rect 5042 2624 5047 2680
rect 1669 2622 5047 2624
rect 6776 2680 6868 2682
rect 6776 2624 6826 2680
rect 6776 2622 6868 2624
rect 1669 2619 1735 2622
rect 4981 2619 5047 2622
rect 6821 2620 6868 2622
rect 6932 2620 6938 2684
rect 6821 2619 6887 2620
rect 0 2546 800 2576
rect 1025 2546 1091 2549
rect 0 2544 1091 2546
rect 0 2488 1030 2544
rect 1086 2488 1091 2544
rect 0 2486 1091 2488
rect 0 2456 800 2486
rect 1025 2483 1091 2486
rect 2405 2546 2471 2549
rect 3693 2546 3759 2549
rect 2405 2544 3759 2546
rect 2405 2488 2410 2544
rect 2466 2488 3698 2544
rect 3754 2488 3759 2544
rect 2405 2486 3759 2488
rect 2405 2483 2471 2486
rect 3693 2483 3759 2486
rect 4409 2208 4729 2209
rect 0 2138 800 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 800 2078
rect 4061 2075 4127 2078
rect 0 1594 800 1624
rect 1209 1594 1275 1597
rect 0 1592 1275 1594
rect 0 1536 1214 1592
rect 1270 1536 1275 1592
rect 0 1534 1275 1536
rect 0 1504 800 1534
rect 1209 1531 1275 1534
rect 0 1186 800 1216
rect 3785 1186 3851 1189
rect 0 1184 3851 1186
rect 0 1128 3790 1184
rect 3846 1128 3851 1184
rect 0 1126 3851 1128
rect 0 1096 800 1126
rect 3785 1123 3851 1126
rect 0 642 800 672
rect 3141 642 3207 645
rect 0 640 3207 642
rect 0 584 3146 640
rect 3202 584 3207 640
rect 0 582 3207 584
rect 0 552 800 582
rect 3141 579 3207 582
rect 0 234 800 264
rect 1485 234 1551 237
rect 0 232 1551 234
rect 0 176 1490 232
rect 1546 176 1551 232
rect 0 174 1551 176
rect 0 144 800 174
rect 1485 171 1551 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 4844 11460 4908 11524
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4108 10236 4172 10300
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 4108 9692 4172 9756
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 6868 8196 6932 8260
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 6868 7380 6932 7444
rect 5580 7168 5644 7172
rect 5580 7112 5594 7168
rect 5594 7112 5644 7168
rect 5580 7108 5644 7112
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 5764 4932 5828 4996
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 5764 4660 5828 4724
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 5580 3164 5644 3228
rect 4844 2952 4908 2956
rect 4844 2896 4894 2952
rect 4894 2896 4908 2952
rect 4844 2892 4908 2896
rect 5764 2756 5828 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 6868 2680 6932 2684
rect 6868 2624 6882 2680
rect 6882 2624 6932 2680
rect 6868 2620 6932 2624
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 4843 11524 4909 11525
rect 4843 11460 4844 11524
rect 4908 11460 4909 11524
rect 4843 11459 4909 11460
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4107 10300 4173 10301
rect 4107 10236 4108 10300
rect 4172 10236 4173 10300
rect 4107 10235 4173 10236
rect 4110 9757 4170 10235
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4107 9756 4173 9757
rect 4107 9692 4108 9756
rect 4172 9692 4173 9756
rect 4107 9691 4173 9692
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4846 2957 4906 11459
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 6867 8260 6933 8261
rect 6867 8196 6868 8260
rect 6932 8196 6933 8260
rect 6867 8195 6933 8196
rect 6870 7445 6930 8195
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 6867 7444 6933 7445
rect 6867 7380 6868 7444
rect 6932 7380 6933 7444
rect 6867 7379 6933 7380
rect 5579 7172 5645 7173
rect 5579 7108 5580 7172
rect 5644 7108 5645 7172
rect 5579 7107 5645 7108
rect 5582 3229 5642 7107
rect 5763 4996 5829 4997
rect 5763 4932 5764 4996
rect 5828 4932 5829 4996
rect 5763 4931 5829 4932
rect 5766 4725 5826 4931
rect 5763 4724 5829 4725
rect 5763 4660 5764 4724
rect 5828 4660 5829 4724
rect 5763 4659 5829 4660
rect 5579 3228 5645 3229
rect 5579 3164 5580 3228
rect 5644 3164 5645 3228
rect 5579 3163 5645 3164
rect 4843 2956 4909 2957
rect 4843 2892 4844 2956
rect 4908 2892 4909 2956
rect 4843 2891 4909 2892
rect 5766 2821 5826 4659
rect 5763 2820 5829 2821
rect 5763 2756 5764 2820
rect 5828 2756 5829 2820
rect 5763 2755 5829 2756
rect 6870 2685 6930 7379
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 6867 2684 6933 2685
rect 6867 2620 6868 2684
rect 6932 2620 6933 2684
rect 6867 2619 6933 2620
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3588 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1624635492
transform 1 0 2208 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2208 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input71 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform -1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4416 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform -1 0 4876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1624635492
transform -1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1624635492
transform -1 0 3772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1624635492
transform -1 0 4232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform -1 0 5520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1624635492
transform -1 0 6348 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1624635492
transform -1 0 6256 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1624635492
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8924 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1624635492
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 8924 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1624635492
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12236 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1624635492
transform -1 0 12696 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624635492
transform -1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 12236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 13984 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 14536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 13064 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform -1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform -1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_146
timestamp 1624635492
transform 1 0 14536 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform -1 0 15272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform -1 0 14904 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 15180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_153
timestamp 1624635492
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform -1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform -1 0 15548 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 16100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_163
timestamp 1624635492
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1624635492
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform -1 0 16468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 16468 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1624635492
transform 1 0 16744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1624635492
transform 1 0 16468 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform -1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 16744 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624635492
transform -1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform -1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform -1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform -1 0 17388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1624635492
transform 1 0 17388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform -1 0 17848 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform 1 0 17572 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform -1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform 1 0 18124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform -1 0 18124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1624635492
transform -1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 18768 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1624635492
transform -1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform -1 0 19320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform -1 0 19320 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1624635492
transform 1 0 19320 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_198
timestamp 1624635492
transform 1 0 19320 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1624635492
transform -1 0 19872 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform -1 0 19780 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform -1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_206
timestamp 1624635492
transform 1 0 20056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1624635492
transform -1 0 20056 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform -1 0 20240 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 1624635492
transform 1 0 20240 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1624635492
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_212
timestamp 1624635492
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_213
timestamp 1624635492
transform 1 0 20700 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform -1 0 20700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform -1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1624635492
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform -1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform -1 0 21252 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform 1 0 21252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform -1 0 21620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3128 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1624635492
transform 1 0 3128 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1624635492
transform -1 0 6256 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7084 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1624635492
transform 1 0 5336 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7544 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform 1 0 8556 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform -1 0 7452 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_69
timestamp 1624635492
transform 1 0 7452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 10120 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1624635492
transform -1 0 9936 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 10120 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1624635492
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 11592 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_126
timestamp 1624635492
transform 1 0 12696 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 13616 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13340 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 13064 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_140
timestamp 1624635492
transform 1 0 13984 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1624635492
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1624635492
transform -1 0 15364 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1624635492
transform -1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1624635492
transform -1 0 16192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_164 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16192 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform -1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1624635492
transform -1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_176 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 17296 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_189
timestamp 1624635492
transform 1 0 18492 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1624635492
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_213
timestamp 1624635492
transform 1 0 20700 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 1748 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5888 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform 1 0 3496 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1624635492
transform 1 0 4048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1624635492
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 5888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1624635492
transform -1 0 8280 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1624635492
transform -1 0 9108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1624635492
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1624635492
transform -1 0 12604 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1624635492
transform -1 0 12880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 15088 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1624635492
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform -1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1624635492
transform 1 0 15272 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16376 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_170
timestamp 1624635492
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_177
timestamp 1624635492
transform 1 0 17388 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_189
timestamp 1624635492
transform 1 0 18492 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_201
timestamp 1624635492
transform 1 0 19596 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_213
timestamp 1624635492
transform 1 0 20700 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1624635492
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2024 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 2852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5980 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1624635492
transform 1 0 5980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624635492
transform -1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1624635492
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1624635492
transform -1 0 8464 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform -1 0 8832 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1624635492
transform -1 0 10488 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 9476 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1624635492
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1624635492
transform 1 0 10764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 1624635492
transform 1 0 11132 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15180 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1624635492
transform -1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1624635492
transform 1 0 13708 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1624635492
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1624635492
transform 1 0 15180 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1624635492
transform -1 0 17664 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1624635492
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform -1 0 20240 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1624635492
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1624635492
transform 1 0 20240 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_220
timestamp 1624635492
transform 1 0 21344 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1840 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1624635492
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1624635492
transform -1 0 4140 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 4508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1624635492
transform 1 0 4508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1624635492
transform -1 0 7452 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 5612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624635492
transform -1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624635492
transform -1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624635492
transform -1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624635492
transform -1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624635492
transform -1 0 6624 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8924 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1624635492
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1624635492
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_124 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 12512 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 13064 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15364 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15364 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 18124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_185
timestamp 1624635492
transform 1 0 18124 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp 1624635492
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_199
timestamp 1624635492
transform 1 0 19412 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_211
timestamp 1624635492
transform 1 0 20516 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3220 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 1840 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6
timestamp 1624635492
transform 1 0 1656 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1624635492
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1624635492
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4324 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4692 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624635492
transform -1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1624635492
transform 1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1624635492
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_56
timestamp 1624635492
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_53
timestamp 1624635492
transform 1 0 5980 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 6992 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 7912 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7912 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7820 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7820 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10764 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 10488 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1624635492
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_111
timestamp 1624635492
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10764 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 1624635492
transform 1 0 12512 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_118
timestamp 1624635492
transform 1 0 11960 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1624635492
transform -1 0 12604 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1624635492
transform 1 0 12604 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15272 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 15180 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1624635492
transform 1 0 13708 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1624635492
transform 1 0 15272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 16008 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1624635492
transform -1 0 16008 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp 1624635492
transform 1 0 15548 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1624635492
transform 1 0 16284 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1624635492
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1624635492
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_199
timestamp 1624635492
transform 1 0 19412 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_188
timestamp 1624635492
transform 1 0 18400 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_200
timestamp 1624635492
transform 1 0 19504 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1624635492
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_213
timestamp 1624635492
transform 1 0 20700 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_217
timestamp 1624635492
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_212
timestamp 1624635492
transform 1 0 20608 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 1624635492
transform 1 0 21344 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1624635492
transform -1 0 3772 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1624635492
transform 1 0 1656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1624635492
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1624635492
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_79
timestamp 1624635492
transform 1 0 8372 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform 1 0 10120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1624635492
transform -1 0 10120 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624635492
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1624635492
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 12328 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 12604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1624635492
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_125
timestamp 1624635492
transform 1 0 12604 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 15180 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_137
timestamp 1624635492
transform 1 0 13708 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1624635492
transform 1 0 15180 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1624635492
transform 1 0 16284 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1624635492
transform 1 0 17388 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_189
timestamp 1624635492
transform 1 0 18492 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1624635492
transform 1 0 19228 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1624635492
transform 1 0 20700 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1624635492
transform 1 0 21436 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1624635492
transform 1 0 2300 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1624635492
transform 1 0 1656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform -1 0 2208 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_12
timestamp 1624635492
transform 1 0 2208 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1624635492
transform 1 0 3404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1624635492
transform -1 0 6348 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 1624635492
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1624635492
transform 1 0 7268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1624635492
transform -1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_100
timestamp 1624635492
transform 1 0 10304 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12788 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14904 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1624635492
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_139
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1624635492
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1624635492
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1624635492
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1624635492
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1624635492
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 2852 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2852 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5888 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1624635492
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_52
timestamp 1624635492
transform 1 0 5888 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_56
timestamp 1624635492
transform 1 0 6256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_77
timestamp 1624635492
transform 1 0 8188 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10396 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9200 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1624635492
transform 1 0 8924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1624635492
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_117
timestamp 1624635492
transform 1 0 11868 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_123
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1624635492
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_176
timestamp 1624635492
transform 1 0 17296 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_188
timestamp 1624635492
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1624635492
transform 1 0 20700 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1624635492
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3312 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 1840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform -1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1624635492
transform -1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp 1624635492
transform 1 0 4324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1624635492
transform -1 0 9200 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7820 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1624635492
transform 1 0 7452 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp 1624635492
transform 1 0 8096 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform 1 0 10028 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1624635492
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1624635492
transform 1 0 10304 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_118
timestamp 1624635492
transform 1 0 11960 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_124
timestamp 1624635492
transform 1 0 12512 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1624635492
transform 1 0 13616 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1624635492
transform 1 0 14444 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_155
timestamp 1624635492
transform 1 0 15364 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_167
timestamp 1624635492
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1624635492
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1624635492
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1624635492
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1624635492
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1624635492
transform 1 0 2668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4324 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7636 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1624635492
transform 1 0 7268 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10580 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1624635492
transform 1 0 10580 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11776 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1624635492
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1624635492
transform -1 0 14076 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13248 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1624635492
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_151
timestamp 1624635492
transform 1 0 14996 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_163
timestamp 1624635492
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_175
timestamp 1624635492
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_187
timestamp 1624635492
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1624635492
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_213
timestamp 1624635492
transform 1 0 20700 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1624635492
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform -1 0 2208 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624635492
transform 1 0 1656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 1932 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_12
timestamp 1624635492
transform 1 0 2208 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 3772 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5336 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4876 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_22
timestamp 1624635492
transform 1 0 3128 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 1624635492
transform 1 0 3864 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_40
timestamp 1624635492
transform 1 0 4784 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1624635492
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8280 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_50
timestamp 1624635492
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1624635492
transform 1 0 6256 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_49
timestamp 1624635492
transform 1 0 5612 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1624635492
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1624635492
transform 1 0 8096 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9292 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9936 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9936 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9016 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1624635492
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform 1 0 12512 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1624635492
transform -1 0 12512 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11592 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_105
timestamp 1624635492
transform 1 0 10764 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1624635492
transform 1 0 11316 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15916 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13800 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1624635492
transform -1 0 14628 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1624635492
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp 1624635492
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1624635492
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1624635492
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_161
timestamp 1624635492
transform 1 0 15916 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1624635492
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_173
timestamp 1624635492
transform 1 0 17020 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_185
timestamp 1624635492
transform 1 0 18124 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1624635492
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1624635492
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1624635492
transform 1 0 19228 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1624635492
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1624635492
transform 1 0 20700 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1624635492
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1748 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_6
timestamp 1624635492
transform 1 0 1656 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4232 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp 1624635492
transform 1 0 3220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1624635492
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1624635492
transform -1 0 7360 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1624635492
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8372 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1624635492
transform -1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1624635492
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_95
timestamp 1624635492
transform 1 0 9844 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1624635492
transform 1 0 10212 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform -1 0 12512 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_111
timestamp 1624635492
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_124
timestamp 1624635492
transform 1 0 12512 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12696 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14996 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1624635492
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1624635492
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1624635492
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1624635492
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1624635492
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1624635492
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1624635492
transform 1 0 2300 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624635492
transform 1 0 1656 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1624635492
transform -1 0 5520 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_24
timestamp 1624635492
transform 1 0 3312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1624635492
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1624635492
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6532 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_48
timestamp 1624635492
transform 1 0 5520 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 1624635492
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1624635492
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11868 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_96
timestamp 1624635492
transform 1 0 9936 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12696 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12696 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14444 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_135
timestamp 1624635492
transform 1 0 13524 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_157
timestamp 1624635492
transform 1 0 15548 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_169
timestamp 1624635492
transform 1 0 16652 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_181
timestamp 1624635492
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_193
timestamp 1624635492
transform 1 0 18860 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_199
timestamp 1624635492
transform 1 0 19412 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_213
timestamp 1624635492
transform 1 0 20700 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1624635492
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_26
timestamp 1624635492
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1624635492
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5796 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1624635492
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_62
timestamp 1624635492
transform 1 0 6808 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform 1 0 6900 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 7176 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1624635492
transform 1 0 8648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9844 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_95
timestamp 1624635492
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1624635492
transform 1 0 10212 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_111
timestamp 1624635492
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1624635492
transform -1 0 14996 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_133
timestamp 1624635492
transform 1 0 13340 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1624635492
transform 1 0 14076 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16560 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_168
timestamp 1624635492
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1624635492
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1624635492
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1624635492
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1624635492
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3496 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 1932 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1624635492
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4140 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1624635492
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 5612 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1624635492
transform 1 0 7084 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_77
timestamp 1624635492
transform 1 0 8188 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9292 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624635492
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10764 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 15824 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1624635492
transform 1 0 13064 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1624635492
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 15824 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_169
timestamp 1624635492
transform 1 0 16652 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_181
timestamp 1624635492
transform 1 0 17756 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_193
timestamp 1624635492
transform 1 0 18860 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1624635492
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_213
timestamp 1624635492
transform 1 0 20700 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1624635492
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1624635492
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_18
timestamp 1624635492
transform 1 0 2760 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1624635492
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_24
timestamp 1624635492
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3496 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1624635492
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1624635492
transform 1 0 4508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5980 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_49
timestamp 1624635492
transform 1 0 5612 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7912 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1624635492
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10212 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11132 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 10212 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1624635492
transform 1 0 10212 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_101
timestamp 1624635492
transform 1 0 10396 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 11408 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12236 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_109
timestamp 1624635492
transform 1 0 11132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624635492
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_109
timestamp 1624635492
transform 1 0 11132 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 14352 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_138
timestamp 1624635492
transform 1 0 13800 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_139
timestamp 1624635492
transform 1 0 13892 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15364 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_155
timestamp 1624635492
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_160
timestamp 1624635492
transform 1 0 15824 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18400 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1624635492
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_172
timestamp 1624635492
transform 1 0 16928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1624635492
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_188
timestamp 1624635492
transform 1 0 18400 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_200
timestamp 1624635492
transform 1 0 19504 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_196
timestamp 1624635492
transform 1 0 19136 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_212
timestamp 1624635492
transform 1 0 20608 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1624635492
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_213
timestamp 1624635492
transform 1 0 20700 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1624635492
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1624635492
transform 1 0 2024 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform 1 0 2300 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1624635492
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_34
timestamp 1624635492
transform 1 0 4232 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_38
timestamp 1624635492
transform 1 0 4600 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 7636 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_48
timestamp 1624635492
transform 1 0 5520 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1624635492
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9292 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9292 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1624635492
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1624635492
transform -1 0 11868 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1624635492
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1624635492
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1624635492
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 13800 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_138
timestamp 1624635492
transform 1 0 13800 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1624635492
transform 1 0 14536 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1624635492
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1624635492
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1624635492
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1624635492
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1624635492
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1624635492
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform 1 0 2024 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1624635492
transform -1 0 3772 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1624635492
transform 1 0 2300 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_19
timestamp 1624635492
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5336 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp 1624635492
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1624635492
transform -1 0 7176 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7268 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1624635492
transform 1 0 7176 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_76
timestamp 1624635492
transform 1 0 8096 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10396 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9568 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_94
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_100
timestamp 1624635492
transform 1 0 10304 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1624635492
transform -1 0 13064 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 11500 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1624635492
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp 1624635492
transform 1 0 11500 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform 1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14444 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1624635492
transform 1 0 13064 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_142
timestamp 1624635492
transform 1 0 14168 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_161
timestamp 1624635492
transform 1 0 15916 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_173
timestamp 1624635492
transform 1 0 17020 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_185
timestamp 1624635492
transform 1 0 18124 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1624635492
transform 1 0 19228 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_213
timestamp 1624635492
transform 1 0 20700 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_7
timestamp 1624635492
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_16
timestamp 1624635492
transform 1 0 2576 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_35
timestamp 1624635492
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7912 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_47
timestamp 1624635492
transform 1 0 5428 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7912 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_23_83
timestamp 1624635492
transform 1 0 8740 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9844 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1624635492
transform -1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1624635492
transform -1 0 13340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_111
timestamp 1624635492
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 13340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15088 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1624635492
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1624635492
transform 1 0 15272 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_166
timestamp 1624635492
transform 1 0 16376 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1624635492
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1624635492
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1624635492
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1624635492
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1624635492
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 2024 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform -1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_16
timestamp 1624635492
transform 1 0 2576 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1624635492
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1624635492
transform -1 0 4784 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624635492
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6716 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_45
timestamp 1624635492
transform 1 0 5244 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1624635492
transform 1 0 6348 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_79
timestamp 1624635492
transform 1 0 8372 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1624635492
transform -1 0 10304 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624635492
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1624635492
transform 1 0 10304 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11224 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 12696 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_160
timestamp 1624635492
transform 1 0 15824 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1624635492
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1624635492
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1624635492
transform 1 0 19136 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1624635492
transform 1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_10
timestamp 1624635492
transform 1 0 2024 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_14
timestamp 1624635492
transform 1 0 2392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3864 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1624635492
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 6716 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_46
timestamp 1624635492
transform 1 0 5336 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_54
timestamp 1624635492
transform 1 0 6072 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1624635492
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_64
timestamp 1624635492
transform 1 0 6992 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1624635492
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1624635492
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12512 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_110
timestamp 1624635492
transform 1 0 11224 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_124
timestamp 1624635492
transform 1 0 12512 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1624635492
transform -1 0 13524 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1624635492
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1624635492
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1624635492
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1624635492
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1624635492
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1624635492
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1624635492
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform -1 0 2116 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform -1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform -1 0 2024 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_17
timestamp 1624635492
transform 1 0 2668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1624635492
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624635492
transform -1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624635492
transform -1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3404 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2300 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3404 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4876 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3956 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1624635492
transform -1 0 3496 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_23
timestamp 1624635492
transform 1 0 3220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1624635492
transform 1 0 4784 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5152 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1624635492
transform -1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7912 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1624635492
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10856 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9752 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11500 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9568 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1624635492
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1624635492
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_103
timestamp 1624635492
transform 1 0 10580 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12328 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_126
timestamp 1624635492
transform 1 0 12696 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_138
timestamp 1624635492
transform 1 0 13800 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1624635492
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_134
timestamp 1624635492
transform 1 0 13432 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1624635492
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_146
timestamp 1624635492
transform 1 0 14536 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_158
timestamp 1624635492
transform 1 0 15640 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1624635492
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1624635492
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_170
timestamp 1624635492
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1624635492
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1624635492
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1624635492
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1624635492
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_213
timestamp 1624635492
transform 1 0 20700 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1624635492
transform 1 0 20976 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform 1 0 1748 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform -1 0 2300 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2852 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3956 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624635492
transform -1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624635492
transform -1 0 3496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624635492
transform -1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624635492
transform -1 0 4968 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_28
timestamp 1624635492
transform 1 0 3680 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6716 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624635492
transform -1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_46
timestamp 1624635492
transform 1 0 5336 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1624635492
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1624635492
transform 1 0 7544 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_73
timestamp 1624635492
transform 1 0 7820 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform 1 0 9200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9752 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_91
timestamp 1624635492
transform 1 0 9476 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11776 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_28_110
timestamp 1624635492
transform 1 0 11224 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1624635492
transform -1 0 13800 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_132
timestamp 1624635492
transform 1 0 13248 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1624635492
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1624635492
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1624635492
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1624635492
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1624635492
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1624635492
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_213
timestamp 1624635492
transform 1 0 20700 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform 1 0 1748 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 2576 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1624635492
transform 1 0 2024 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1624635492
transform 1 0 2300 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform -1 0 4324 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4324 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624635492
transform -1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1624635492
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6624 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 6624 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1624635492
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1624635492
transform 1 0 7084 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1624635492
transform 1 0 7360 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1624635492
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1624635492
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1624635492
transform 1 0 9660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_105
timestamp 1624635492
transform 1 0 10764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1624635492
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_124
timestamp 1624635492
transform 1 0 12512 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_136
timestamp 1624635492
transform 1 0 13616 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_148
timestamp 1624635492
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1624635492
transform 1 0 15824 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_168
timestamp 1624635492
transform 1 0 16560 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1624635492
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1624635492
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1624635492
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform 1 0 1748 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform 1 0 2024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform -1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1624635492
transform 1 0 3128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1624635492
transform 1 0 3404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1624635492
transform 1 0 4692 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1624635492
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6532 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_42
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624635492
transform -1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_83
timestamp 1624635492
transform 1 0 8740 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 10120 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11592 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_114
timestamp 1624635492
transform 1 0 11592 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14260 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1624635492
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_128
timestamp 1624635492
transform 1 0 12880 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_134
timestamp 1624635492
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1624635492
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1624635492
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15088 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1624635492
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1624635492
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1624635492
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1624635492
transform 1 0 15088 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_158
timestamp 1624635492
transform 1 0 15640 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_162
timestamp 1624635492
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_165
timestamp 1624635492
transform 1 0 16284 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16928 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1624635492
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1624635492
transform 1 0 16560 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_172
timestamp 1624635492
transform 1 0 16928 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1624635492
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1624635492
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_190
timestamp 1624635492
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_194
timestamp 1624635492
transform 1 0 18952 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_213
timestamp 1624635492
transform 1 0 20700 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform 1 0 2024 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3128 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4600 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4600 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform -1 0 7084 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 6072 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6532 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8556 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8556 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform -1 0 9108 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10580 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 10764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1624635492
transform -1 0 13432 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1624635492
transform -1 0 13708 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1624635492
transform -1 0 13984 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1624635492
transform -1 0 14720 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1624635492
transform -1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1624635492
transform -1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform -1 0 15088 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1624635492
transform -1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1624635492
transform -1 0 15916 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1624635492
transform -1 0 16192 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1624635492
transform -1 0 16560 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1624635492
transform -1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_148
timestamp 1624635492
transform 1 0 14720 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1624635492
transform 1 0 15548 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_164
timestamp 1624635492
transform 1 0 16192 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1624635492
transform -1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1624635492
transform -1 0 18584 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1624635492
transform -1 0 16836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1624635492
transform -1 0 18860 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1624635492
transform -1 0 19320 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1624635492
transform -1 0 19872 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1624635492
transform -1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_200
timestamp 1624635492
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_204
timestamp 1624635492
transform 1 0 19872 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_216
timestamp 1624635492
transform 1 0 20976 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1624635492
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform -1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1624635492
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1624635492
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1624635492
transform 1 0 4784 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1624635492
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_39
timestamp 1624635492
transform 1 0 4692 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6532 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1624635492
transform -1 0 6900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_59
timestamp 1624635492
transform 1 0 6532 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8372 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1624635492
transform -1 0 8740 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1624635492
transform 1 0 8740 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10580 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10580 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12328 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12696 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_122
timestamp 1624635492
transform 1 0 12328 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1624635492
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1624635492
transform 1 0 13156 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 13984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1624635492
transform -1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_140
timestamp 1624635492
transform 1 0 13984 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_146
timestamp 1624635492
transform 1 0 14536 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_158
timestamp 1624635492
transform 1 0 15640 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1624635492
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1624635492
transform -1 0 17020 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624635492
transform -1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1624635492
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_179
timestamp 1624635492
transform 1 0 17572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_191
timestamp 1624635492
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1624635492
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624635492
transform -1 0 21620 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_213
timestamp 1624635492
transform 1 0 20700 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 2852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1624635492
transform 1 0 4324 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1624635492
transform 1 0 4692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_38
timestamp 1624635492
transform 1 0 4600 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5060 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1624635492
transform 1 0 5888 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624635492
transform -1 0 8832 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1624635492
transform -1 0 8096 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1624635492
transform -1 0 8464 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1624635492
transform 1 0 8832 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1624635492
transform -1 0 10396 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1624635492
transform -1 0 10764 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1624635492
transform 1 0 10764 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1624635492
transform 1 0 12604 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1624635492
transform -1 0 11592 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1624635492
transform -1 0 12236 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1624635492
transform -1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_109
timestamp 1624635492
transform 1 0 11132 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform -1 0 13432 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624635492
transform -1 0 13892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624635492
transform -1 0 14352 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 13064 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_134
timestamp 1624635492
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1624635492
transform 1 0 13892 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1624635492
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624635492
transform -1 0 14904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624635492
transform -1 0 15272 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624635492
transform -1 0 15732 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624635492
transform -1 0 16192 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624635492
transform -1 0 16652 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_154
timestamp 1624635492
transform 1 0 15272 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_159
timestamp 1624635492
transform 1 0 15732 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_164
timestamp 1624635492
transform 1 0 16192 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform -1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform -1 0 18492 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624635492
transform 1 0 17296 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624635492
transform -1 0 17112 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1624635492
transform 1 0 16652 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_184
timestamp 1624635492
transform 1 0 18032 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform -1 0 18952 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1624635492
transform -1 0 19412 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624635492
transform -1 0 20240 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624635492
transform -1 0 20608 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624635492
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1624635492
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_194
timestamp 1624635492
transform 1 0 18952 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1624635492
transform -1 0 21620 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624635492
transform -1 0 20976 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624635492
transform -1 0 21344 0 1 20128
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 0 nsew signal input
rlabel metal2 s 662 0 718 800 6 bottom_left_grid_pin_43_
port 1 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 bottom_left_grid_pin_44_
port 2 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 bottom_left_grid_pin_45_
port 3 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_46_
port 4 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 bottom_left_grid_pin_47_
port 5 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_48_
port 6 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 bottom_left_grid_pin_49_
port 7 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 bottom_right_grid_pin_1_
port 8 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 10 nsew signal tristate
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[0]
port 11 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[10]
port 12 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[11]
port 13 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[12]
port 14 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[13]
port 15 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 16 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 17 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[16]
port 18 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[17]
port 19 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[18]
port 20 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 21 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 22 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[2]
port 23 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[3]
port 24 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[4]
port 25 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[5]
port 26 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[6]
port 27 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[7]
port 28 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[8]
port 29 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[9]
port 30 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 31 nsew signal tristate
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 32 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 33 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 34 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 35 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 36 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 37 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 38 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 39 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 40 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 41 nsew signal tristate
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[1]
port 42 nsew signal tristate
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[2]
port 43 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 44 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 45 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[5]
port 46 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[6]
port 47 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[7]
port 48 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 49 nsew signal tristate
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[9]
port 50 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 51 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[10]
port 52 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[11]
port 53 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 54 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[13]
port 55 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[14]
port 56 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[15]
port 57 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[16]
port 58 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[17]
port 59 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[18]
port 60 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[19]
port 61 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[1]
port 62 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_in[2]
port 63 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[3]
port 64 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[4]
port 65 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[5]
port 66 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[6]
port 67 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[7]
port 68 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 69 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 70 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[0]
port 71 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 chany_bottom_out[10]
port 72 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[11]
port 73 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[12]
port 74 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[13]
port 75 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 76 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 chany_bottom_out[15]
port 77 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[16]
port 78 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 chany_bottom_out[17]
port 79 nsew signal tristate
rlabel metal2 s 21730 0 21786 800 6 chany_bottom_out[18]
port 80 nsew signal tristate
rlabel metal2 s 22190 0 22246 800 6 chany_bottom_out[19]
port 81 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[1]
port 82 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[2]
port 83 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[3]
port 84 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[4]
port 85 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[5]
port 86 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[6]
port 87 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[7]
port 88 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[8]
port 89 nsew signal tristate
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[9]
port 90 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 91 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 92 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 93 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 94 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 95 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 96 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 97 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 98 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 99 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 100 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 101 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 102 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 103 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 104 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 105 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 106 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 107 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 108 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 109 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 110 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 111 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 112 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 113 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 114 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 115 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 116 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 117 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 118 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 119 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 120 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 121 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 122 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 123 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 124 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 125 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 126 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 127 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 128 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 129 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 130 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 131 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 132 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 left_bottom_grid_pin_36_
port 133 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 134 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_38_
port 135 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 136 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_40_
port 137 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 138 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 139 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 140 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 141 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 142 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 143 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 144 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 145 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 146 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 147 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 148 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 149 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 150 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 151 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 152 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 153 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
