VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_left_tile
  CLASS BLOCK ;
  FOREIGN top_left_tile ;
  ORIGIN 0.000 0.000 ;
  SIZE 135.000 BY 285.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.720 10.640 91.320 272.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.720 10.640 16.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 10.640 66.320 272.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 10.640 116.320 272.240 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 281.000 129.630 285.000 ;
    END
  END ccff_head
  PIN ccff_head_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END ccff_head_0
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 3.440 135.000 4.040 ;
    END
  END ccff_tail
  PIN ccff_tail_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 281.000 5.430 285.000 ;
    END
  END ccff_tail_0
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 129.920 135.000 130.520 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 170.720 135.000 171.320 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 174.800 135.000 175.400 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 178.880 135.000 179.480 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 182.960 135.000 183.560 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 187.040 135.000 187.640 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 191.120 135.000 191.720 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 195.200 135.000 195.800 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 199.280 135.000 199.880 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 203.360 135.000 203.960 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 207.440 135.000 208.040 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 134.000 135.000 134.600 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 211.520 135.000 212.120 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 215.600 135.000 216.200 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 219.680 135.000 220.280 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 223.760 135.000 224.360 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 227.840 135.000 228.440 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 231.920 135.000 232.520 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 236.000 135.000 236.600 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 240.080 135.000 240.680 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 244.160 135.000 244.760 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 248.240 135.000 248.840 ;
    END
  END chanx_right_in[29]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 138.080 135.000 138.680 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 142.160 135.000 142.760 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 146.240 135.000 146.840 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 150.320 135.000 150.920 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 154.400 135.000 155.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 158.480 135.000 159.080 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 162.560 135.000 163.160 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 166.640 135.000 167.240 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 7.520 135.000 8.120 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 48.320 135.000 48.920 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 52.400 135.000 53.000 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 56.480 135.000 57.080 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 60.560 135.000 61.160 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 64.640 135.000 65.240 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 68.720 135.000 69.320 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 72.800 135.000 73.400 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 76.880 135.000 77.480 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 80.960 135.000 81.560 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 85.040 135.000 85.640 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 11.600 135.000 12.200 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 89.120 135.000 89.720 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 93.200 135.000 93.800 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 97.280 135.000 97.880 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 101.360 135.000 101.960 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 105.440 135.000 106.040 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 109.520 135.000 110.120 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 113.600 135.000 114.200 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 117.680 135.000 118.280 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 121.760 135.000 122.360 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 125.840 135.000 126.440 ;
    END
  END chanx_right_out[29]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 15.680 135.000 16.280 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 19.760 135.000 20.360 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 23.840 135.000 24.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 27.920 135.000 28.520 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 32.000 135.000 32.600 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 36.080 135.000 36.680 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 40.160 135.000 40.760 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 44.240 135.000 44.840 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END chany_bottom_in_0[0]
  PIN chany_bottom_in_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END chany_bottom_in_0[10]
  PIN chany_bottom_in_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END chany_bottom_in_0[11]
  PIN chany_bottom_in_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END chany_bottom_in_0[12]
  PIN chany_bottom_in_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END chany_bottom_in_0[13]
  PIN chany_bottom_in_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END chany_bottom_in_0[14]
  PIN chany_bottom_in_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END chany_bottom_in_0[15]
  PIN chany_bottom_in_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in_0[16]
  PIN chany_bottom_in_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END chany_bottom_in_0[17]
  PIN chany_bottom_in_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END chany_bottom_in_0[18]
  PIN chany_bottom_in_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END chany_bottom_in_0[19]
  PIN chany_bottom_in_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END chany_bottom_in_0[1]
  PIN chany_bottom_in_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END chany_bottom_in_0[20]
  PIN chany_bottom_in_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END chany_bottom_in_0[21]
  PIN chany_bottom_in_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END chany_bottom_in_0[22]
  PIN chany_bottom_in_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END chany_bottom_in_0[23]
  PIN chany_bottom_in_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END chany_bottom_in_0[24]
  PIN chany_bottom_in_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END chany_bottom_in_0[25]
  PIN chany_bottom_in_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END chany_bottom_in_0[26]
  PIN chany_bottom_in_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END chany_bottom_in_0[27]
  PIN chany_bottom_in_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END chany_bottom_in_0[28]
  PIN chany_bottom_in_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END chany_bottom_in_0[29]
  PIN chany_bottom_in_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END chany_bottom_in_0[2]
  PIN chany_bottom_in_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END chany_bottom_in_0[3]
  PIN chany_bottom_in_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END chany_bottom_in_0[4]
  PIN chany_bottom_in_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END chany_bottom_in_0[5]
  PIN chany_bottom_in_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END chany_bottom_in_0[6]
  PIN chany_bottom_in_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END chany_bottom_in_0[7]
  PIN chany_bottom_in_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END chany_bottom_in_0[8]
  PIN chany_bottom_in_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chany_bottom_in_0[9]
  PIN chany_bottom_out_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END chany_bottom_out_0[0]
  PIN chany_bottom_out_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END chany_bottom_out_0[10]
  PIN chany_bottom_out_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END chany_bottom_out_0[11]
  PIN chany_bottom_out_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END chany_bottom_out_0[12]
  PIN chany_bottom_out_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END chany_bottom_out_0[13]
  PIN chany_bottom_out_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chany_bottom_out_0[14]
  PIN chany_bottom_out_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END chany_bottom_out_0[15]
  PIN chany_bottom_out_0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END chany_bottom_out_0[16]
  PIN chany_bottom_out_0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END chany_bottom_out_0[17]
  PIN chany_bottom_out_0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END chany_bottom_out_0[18]
  PIN chany_bottom_out_0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END chany_bottom_out_0[19]
  PIN chany_bottom_out_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END chany_bottom_out_0[1]
  PIN chany_bottom_out_0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END chany_bottom_out_0[20]
  PIN chany_bottom_out_0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END chany_bottom_out_0[21]
  PIN chany_bottom_out_0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END chany_bottom_out_0[22]
  PIN chany_bottom_out_0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END chany_bottom_out_0[23]
  PIN chany_bottom_out_0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END chany_bottom_out_0[24]
  PIN chany_bottom_out_0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END chany_bottom_out_0[25]
  PIN chany_bottom_out_0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END chany_bottom_out_0[26]
  PIN chany_bottom_out_0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END chany_bottom_out_0[27]
  PIN chany_bottom_out_0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END chany_bottom_out_0[28]
  PIN chany_bottom_out_0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END chany_bottom_out_0[29]
  PIN chany_bottom_out_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END chany_bottom_out_0[2]
  PIN chany_bottom_out_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END chany_bottom_out_0[3]
  PIN chany_bottom_out_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END chany_bottom_out_0[4]
  PIN chany_bottom_out_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END chany_bottom_out_0[5]
  PIN chany_bottom_out_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END chany_bottom_out_0[6]
  PIN chany_bottom_out_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END chany_bottom_out_0[7]
  PIN chany_bottom_out_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END chany_bottom_out_0[8]
  PIN chany_bottom_out_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END chany_bottom_out_0[9]
  PIN gfpga_pad_io_soc_dir[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 281.000 12.330 285.000 ;
    END
  END gfpga_pad_io_soc_dir[0]
  PIN gfpga_pad_io_soc_dir[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 281.000 19.230 285.000 ;
    END
  END gfpga_pad_io_soc_dir[1]
  PIN gfpga_pad_io_soc_dir[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 281.000 26.130 285.000 ;
    END
  END gfpga_pad_io_soc_dir[2]
  PIN gfpga_pad_io_soc_dir[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 281.000 33.030 285.000 ;
    END
  END gfpga_pad_io_soc_dir[3]
  PIN gfpga_pad_io_soc_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 281.000 67.530 285.000 ;
    END
  END gfpga_pad_io_soc_in[0]
  PIN gfpga_pad_io_soc_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 281.000 74.430 285.000 ;
    END
  END gfpga_pad_io_soc_in[1]
  PIN gfpga_pad_io_soc_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 281.000 81.330 285.000 ;
    END
  END gfpga_pad_io_soc_in[2]
  PIN gfpga_pad_io_soc_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 281.000 88.230 285.000 ;
    END
  END gfpga_pad_io_soc_in[3]
  PIN gfpga_pad_io_soc_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 281.000 39.930 285.000 ;
    END
  END gfpga_pad_io_soc_out[0]
  PIN gfpga_pad_io_soc_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 281.000 46.830 285.000 ;
    END
  END gfpga_pad_io_soc_out[1]
  PIN gfpga_pad_io_soc_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 281.000 53.730 285.000 ;
    END
  END gfpga_pad_io_soc_out[2]
  PIN gfpga_pad_io_soc_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 281.000 60.630 285.000 ;
    END
  END gfpga_pad_io_soc_out[3]
  PIN isol_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 281.000 95.130 285.000 ;
    END
  END isol_n
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END prog_clk
  PIN prog_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END prog_reset
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END reset
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 252.320 135.000 252.920 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 256.400 135.000 257.000 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 260.480 135.000 261.080 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 264.560 135.000 265.160 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 268.640 135.000 269.240 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 272.720 135.000 273.320 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 276.800 135.000 277.400 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 131.000 280.880 135.000 281.480 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
  PIN right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 281.000 102.030 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 281.000 108.930 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 281.000 115.830 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
  PIN right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 281.000 122.730 285.000 ;
    END
  END right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
  PIN right_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END right_width_0_height_0_subtile_0__pin_inpad_0_
  PIN right_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END right_width_0_height_0_subtile_1__pin_inpad_0_
  PIN right_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END right_width_0_height_0_subtile_2__pin_inpad_0_
  PIN right_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END right_width_0_height_0_subtile_3__pin_inpad_0_
  PIN test_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END test_enable
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 129.260 272.085 ;
      LAYER met1 ;
        RECT 5.130 8.880 134.710 272.240 ;
      LAYER met2 ;
        RECT 5.710 280.720 11.770 281.250 ;
        RECT 12.610 280.720 18.670 281.250 ;
        RECT 19.510 280.720 25.570 281.250 ;
        RECT 26.410 280.720 32.470 281.250 ;
        RECT 33.310 280.720 39.370 281.250 ;
        RECT 40.210 280.720 46.270 281.250 ;
        RECT 47.110 280.720 53.170 281.250 ;
        RECT 54.010 280.720 60.070 281.250 ;
        RECT 60.910 280.720 66.970 281.250 ;
        RECT 67.810 280.720 73.870 281.250 ;
        RECT 74.710 280.720 80.770 281.250 ;
        RECT 81.610 280.720 87.670 281.250 ;
        RECT 88.510 280.720 94.570 281.250 ;
        RECT 95.410 280.720 101.470 281.250 ;
        RECT 102.310 280.720 108.370 281.250 ;
        RECT 109.210 280.720 115.270 281.250 ;
        RECT 116.110 280.720 122.170 281.250 ;
        RECT 123.010 280.720 129.070 281.250 ;
        RECT 129.910 280.720 134.680 281.250 ;
        RECT 5.160 4.280 134.680 280.720 ;
        RECT 5.160 3.555 7.170 4.280 ;
        RECT 8.010 3.555 9.010 4.280 ;
        RECT 9.850 3.555 10.850 4.280 ;
        RECT 11.690 3.555 12.690 4.280 ;
        RECT 13.530 3.555 14.530 4.280 ;
        RECT 15.370 3.555 16.370 4.280 ;
        RECT 17.210 3.555 18.210 4.280 ;
        RECT 19.050 3.555 20.050 4.280 ;
        RECT 20.890 3.555 21.890 4.280 ;
        RECT 22.730 3.555 23.730 4.280 ;
        RECT 24.570 3.555 25.570 4.280 ;
        RECT 26.410 3.555 27.410 4.280 ;
        RECT 28.250 3.555 29.250 4.280 ;
        RECT 30.090 3.555 31.090 4.280 ;
        RECT 31.930 3.555 32.930 4.280 ;
        RECT 33.770 3.555 34.770 4.280 ;
        RECT 35.610 3.555 36.610 4.280 ;
        RECT 37.450 3.555 38.450 4.280 ;
        RECT 39.290 3.555 40.290 4.280 ;
        RECT 41.130 3.555 42.130 4.280 ;
        RECT 42.970 3.555 43.970 4.280 ;
        RECT 44.810 3.555 45.810 4.280 ;
        RECT 46.650 3.555 47.650 4.280 ;
        RECT 48.490 3.555 49.490 4.280 ;
        RECT 50.330 3.555 51.330 4.280 ;
        RECT 52.170 3.555 53.170 4.280 ;
        RECT 54.010 3.555 55.010 4.280 ;
        RECT 55.850 3.555 56.850 4.280 ;
        RECT 57.690 3.555 58.690 4.280 ;
        RECT 59.530 3.555 60.530 4.280 ;
        RECT 61.370 3.555 62.370 4.280 ;
        RECT 63.210 3.555 64.210 4.280 ;
        RECT 65.050 3.555 66.050 4.280 ;
        RECT 66.890 3.555 67.890 4.280 ;
        RECT 68.730 3.555 69.730 4.280 ;
        RECT 70.570 3.555 71.570 4.280 ;
        RECT 72.410 3.555 73.410 4.280 ;
        RECT 74.250 3.555 75.250 4.280 ;
        RECT 76.090 3.555 77.090 4.280 ;
        RECT 77.930 3.555 78.930 4.280 ;
        RECT 79.770 3.555 80.770 4.280 ;
        RECT 81.610 3.555 82.610 4.280 ;
        RECT 83.450 3.555 84.450 4.280 ;
        RECT 85.290 3.555 86.290 4.280 ;
        RECT 87.130 3.555 88.130 4.280 ;
        RECT 88.970 3.555 89.970 4.280 ;
        RECT 90.810 3.555 91.810 4.280 ;
        RECT 92.650 3.555 93.650 4.280 ;
        RECT 94.490 3.555 95.490 4.280 ;
        RECT 96.330 3.555 97.330 4.280 ;
        RECT 98.170 3.555 99.170 4.280 ;
        RECT 100.010 3.555 101.010 4.280 ;
        RECT 101.850 3.555 102.850 4.280 ;
        RECT 103.690 3.555 104.690 4.280 ;
        RECT 105.530 3.555 106.530 4.280 ;
        RECT 107.370 3.555 108.370 4.280 ;
        RECT 109.210 3.555 110.210 4.280 ;
        RECT 111.050 3.555 112.050 4.280 ;
        RECT 112.890 3.555 113.890 4.280 ;
        RECT 114.730 3.555 115.730 4.280 ;
        RECT 116.570 3.555 117.570 4.280 ;
        RECT 118.410 3.555 119.410 4.280 ;
        RECT 120.250 3.555 121.250 4.280 ;
        RECT 122.090 3.555 123.090 4.280 ;
        RECT 123.930 3.555 124.930 4.280 ;
        RECT 125.770 3.555 134.680 4.280 ;
      LAYER met3 ;
        RECT 4.000 280.480 130.600 281.330 ;
        RECT 4.000 277.800 131.955 280.480 ;
        RECT 4.000 276.400 130.600 277.800 ;
        RECT 4.000 273.720 131.955 276.400 ;
        RECT 4.000 272.320 130.600 273.720 ;
        RECT 4.000 269.640 131.955 272.320 ;
        RECT 4.000 268.240 130.600 269.640 ;
        RECT 4.000 265.560 131.955 268.240 ;
        RECT 4.000 264.160 130.600 265.560 ;
        RECT 4.000 261.480 131.955 264.160 ;
        RECT 4.000 260.080 130.600 261.480 ;
        RECT 4.000 257.400 131.955 260.080 ;
        RECT 4.000 256.000 130.600 257.400 ;
        RECT 4.000 253.320 131.955 256.000 ;
        RECT 4.000 251.920 130.600 253.320 ;
        RECT 4.000 249.240 131.955 251.920 ;
        RECT 4.000 247.840 130.600 249.240 ;
        RECT 4.000 245.160 131.955 247.840 ;
        RECT 4.000 243.760 130.600 245.160 ;
        RECT 4.000 241.080 131.955 243.760 ;
        RECT 4.000 239.680 130.600 241.080 ;
        RECT 4.000 237.000 131.955 239.680 ;
        RECT 4.000 235.600 130.600 237.000 ;
        RECT 4.000 232.920 131.955 235.600 ;
        RECT 4.000 231.520 130.600 232.920 ;
        RECT 4.000 228.840 131.955 231.520 ;
        RECT 4.000 227.440 130.600 228.840 ;
        RECT 4.000 224.760 131.955 227.440 ;
        RECT 4.000 223.360 130.600 224.760 ;
        RECT 4.000 220.680 131.955 223.360 ;
        RECT 4.000 219.280 130.600 220.680 ;
        RECT 4.000 216.600 131.955 219.280 ;
        RECT 4.000 215.200 130.600 216.600 ;
        RECT 4.000 212.520 131.955 215.200 ;
        RECT 4.000 211.120 130.600 212.520 ;
        RECT 4.000 208.440 131.955 211.120 ;
        RECT 4.000 207.040 130.600 208.440 ;
        RECT 4.000 204.360 131.955 207.040 ;
        RECT 4.000 202.960 130.600 204.360 ;
        RECT 4.000 200.280 131.955 202.960 ;
        RECT 4.000 198.880 130.600 200.280 ;
        RECT 4.000 196.200 131.955 198.880 ;
        RECT 4.000 194.800 130.600 196.200 ;
        RECT 4.000 192.120 131.955 194.800 ;
        RECT 4.000 190.720 130.600 192.120 ;
        RECT 4.000 188.040 131.955 190.720 ;
        RECT 4.000 186.640 130.600 188.040 ;
        RECT 4.000 183.960 131.955 186.640 ;
        RECT 4.000 182.560 130.600 183.960 ;
        RECT 4.000 179.880 131.955 182.560 ;
        RECT 4.000 178.480 130.600 179.880 ;
        RECT 4.000 175.800 131.955 178.480 ;
        RECT 4.000 174.400 130.600 175.800 ;
        RECT 4.000 171.720 131.955 174.400 ;
        RECT 4.000 170.320 130.600 171.720 ;
        RECT 4.000 167.640 131.955 170.320 ;
        RECT 4.000 166.240 130.600 167.640 ;
        RECT 4.000 163.560 131.955 166.240 ;
        RECT 4.000 162.160 130.600 163.560 ;
        RECT 4.000 159.480 131.955 162.160 ;
        RECT 4.000 158.080 130.600 159.480 ;
        RECT 4.000 155.400 131.955 158.080 ;
        RECT 4.000 154.000 130.600 155.400 ;
        RECT 4.000 151.320 131.955 154.000 ;
        RECT 4.000 149.920 130.600 151.320 ;
        RECT 4.000 147.240 131.955 149.920 ;
        RECT 4.000 145.840 130.600 147.240 ;
        RECT 4.000 143.160 131.955 145.840 ;
        RECT 4.000 141.760 130.600 143.160 ;
        RECT 4.000 139.080 131.955 141.760 ;
        RECT 4.000 137.680 130.600 139.080 ;
        RECT 4.000 135.000 131.955 137.680 ;
        RECT 4.000 133.600 130.600 135.000 ;
        RECT 4.000 130.920 131.955 133.600 ;
        RECT 4.000 129.520 130.600 130.920 ;
        RECT 4.000 126.840 131.955 129.520 ;
        RECT 4.000 125.440 130.600 126.840 ;
        RECT 4.000 122.760 131.955 125.440 ;
        RECT 4.000 121.360 130.600 122.760 ;
        RECT 4.000 118.680 131.955 121.360 ;
        RECT 4.000 117.280 130.600 118.680 ;
        RECT 4.000 114.600 131.955 117.280 ;
        RECT 4.000 113.200 130.600 114.600 ;
        RECT 4.000 110.520 131.955 113.200 ;
        RECT 4.000 109.120 130.600 110.520 ;
        RECT 4.000 106.440 131.955 109.120 ;
        RECT 4.000 105.040 130.600 106.440 ;
        RECT 4.000 102.360 131.955 105.040 ;
        RECT 4.000 100.960 130.600 102.360 ;
        RECT 4.000 98.280 131.955 100.960 ;
        RECT 4.000 96.880 130.600 98.280 ;
        RECT 4.000 94.200 131.955 96.880 ;
        RECT 4.000 92.800 130.600 94.200 ;
        RECT 4.000 90.120 131.955 92.800 ;
        RECT 4.000 88.720 130.600 90.120 ;
        RECT 4.000 86.040 131.955 88.720 ;
        RECT 4.000 84.640 130.600 86.040 ;
        RECT 4.000 81.960 131.955 84.640 ;
        RECT 4.000 80.560 130.600 81.960 ;
        RECT 4.000 77.880 131.955 80.560 ;
        RECT 4.000 76.480 130.600 77.880 ;
        RECT 4.000 73.800 131.955 76.480 ;
        RECT 4.000 72.400 130.600 73.800 ;
        RECT 4.000 69.720 131.955 72.400 ;
        RECT 4.000 68.320 130.600 69.720 ;
        RECT 4.000 65.640 131.955 68.320 ;
        RECT 4.000 64.240 130.600 65.640 ;
        RECT 4.000 61.560 131.955 64.240 ;
        RECT 4.000 60.160 130.600 61.560 ;
        RECT 4.000 57.480 131.955 60.160 ;
        RECT 4.000 56.080 130.600 57.480 ;
        RECT 4.000 53.400 131.955 56.080 ;
        RECT 4.000 52.000 130.600 53.400 ;
        RECT 4.000 49.320 131.955 52.000 ;
        RECT 4.000 47.920 130.600 49.320 ;
        RECT 4.000 45.240 131.955 47.920 ;
        RECT 4.000 44.560 130.600 45.240 ;
        RECT 4.400 43.840 130.600 44.560 ;
        RECT 4.400 43.160 131.955 43.840 ;
        RECT 4.000 41.160 131.955 43.160 ;
        RECT 4.000 39.760 130.600 41.160 ;
        RECT 4.000 37.080 131.955 39.760 ;
        RECT 4.000 35.680 130.600 37.080 ;
        RECT 4.000 33.000 131.955 35.680 ;
        RECT 4.400 31.600 130.600 33.000 ;
        RECT 4.000 28.920 131.955 31.600 ;
        RECT 4.000 27.520 130.600 28.920 ;
        RECT 4.000 24.840 131.955 27.520 ;
        RECT 4.000 23.440 130.600 24.840 ;
        RECT 4.000 21.440 131.955 23.440 ;
        RECT 4.400 20.760 131.955 21.440 ;
        RECT 4.400 20.040 130.600 20.760 ;
        RECT 4.000 19.360 130.600 20.040 ;
        RECT 4.000 16.680 131.955 19.360 ;
        RECT 4.000 15.280 130.600 16.680 ;
        RECT 4.000 12.600 131.955 15.280 ;
        RECT 4.000 11.200 130.600 12.600 ;
        RECT 4.000 9.880 131.955 11.200 ;
        RECT 4.400 8.520 131.955 9.880 ;
        RECT 4.400 8.480 130.600 8.520 ;
        RECT 4.000 7.120 130.600 8.480 ;
        RECT 4.000 4.440 131.955 7.120 ;
        RECT 4.000 3.575 130.600 4.440 ;
      LAYER met4 ;
        RECT 61.935 10.240 64.320 207.225 ;
        RECT 66.720 10.240 89.320 207.225 ;
        RECT 91.720 10.240 114.320 207.225 ;
        RECT 116.720 10.240 123.905 207.225 ;
        RECT 61.935 9.015 123.905 10.240 ;
  END
END top_left_tile
END LIBRARY

